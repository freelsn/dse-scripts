// verilog_out version 6.79.2
// options:  veriloggen jpeg_E.IFF
// bdlpars options:  -DDSE ../rle.cpp
// bdltran options:  -c1000 -s -Zresource_fcnt=GENERATE -Zresource_mcnt=GENERATE -lb /home/shuangnan/share/packages/zynq-1.BLIB -lfl /home/shuangnan/share/packages/zynq-1.FLIB jpeg.IFF -OX -a8196 -Zfu_cnt_incr_rate=0 -tcio 
// timestamp_0: 20180213183027_13048_66414
// timestamp_5: 20180213183033_14589_48057
// timestamp_9: 20180213183049_14589_66745
// timestamp_C: 20180213183049_14589_80597
// timestamp_E: 20180213183050_14589_50370
// timestamp_V: 20180213183053_18897_80448

module jpeg ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,jpeg_in_a04 ,
	jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,jpeg_in_a10 ,
	jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,jpeg_in_a16 ,
	jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,jpeg_in_a22 ,
	jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,jpeg_in_a28 ,
	jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,jpeg_in_a34 ,
	jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,jpeg_in_a40 ,
	jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,jpeg_in_a46 ,
	jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,jpeg_in_a52 ,
	jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,jpeg_in_a58 ,
	jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,jpeg_in_a64 ,
	jpeg_in_a65 ,jpeg_in_a66 ,jpeg_in_a67 ,jpeg_in_a68 ,jpeg_in_a69 ,jpeg_in_a70 ,
	jpeg_in_a71 ,jpeg_in_a72 ,jpeg_in_a73 ,jpeg_in_a74 ,jpeg_in_a75 ,jpeg_in_a76 ,
	jpeg_in_a77 ,jpeg_in_a78 ,jpeg_in_a79 ,jpeg_in_a80 ,jpeg_in_a81 ,jpeg_in_a82 ,
	jpeg_in_a83 ,jpeg_in_a84 ,jpeg_in_a85 ,jpeg_in_a86 ,jpeg_in_a87 ,jpeg_in_a88 ,
	jpeg_in_a89 ,jpeg_in_a90 ,jpeg_in_a91 ,jpeg_in_a92 ,jpeg_in_a93 ,jpeg_in_a94 ,
	jpeg_in_a95 ,jpeg_in_a96 ,jpeg_in_a97 ,jpeg_in_a98 ,jpeg_in_a99 ,jpeg_in_a100 ,
	jpeg_in_a101 ,jpeg_in_a102 ,jpeg_in_a103 ,jpeg_in_a104 ,jpeg_in_a105 ,jpeg_in_a106 ,
	jpeg_in_a107 ,jpeg_in_a108 ,jpeg_in_a109 ,jpeg_in_a110 ,jpeg_in_a111 ,jpeg_in_a112 ,
	jpeg_in_a113 ,jpeg_in_a114 ,jpeg_in_a115 ,jpeg_in_a116 ,jpeg_in_a117 ,jpeg_in_a118 ,
	jpeg_in_a119 ,jpeg_in_a120 ,jpeg_in_a121 ,jpeg_in_a122 ,jpeg_in_a123 ,jpeg_in_a124 ,
	jpeg_in_a125 ,jpeg_in_a126 ,jpeg_in_a127 ,jpeg_len_in ,jpeg_out_a00 ,jpeg_out_a01 ,
	jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,jpeg_out_a06 ,jpeg_out_a07 ,
	jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,jpeg_out_a12 ,jpeg_out_a13 ,
	jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,jpeg_out_a18 ,jpeg_out_a19 ,
	jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,jpeg_out_a24 ,jpeg_out_a25 ,
	jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,jpeg_out_a30 ,jpeg_out_a31 ,
	jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,jpeg_out_a36 ,jpeg_out_a37 ,
	jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,jpeg_out_a42 ,jpeg_out_a43 ,
	jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,jpeg_out_a48 ,jpeg_out_a49 ,
	jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,jpeg_out_a54 ,jpeg_out_a55 ,
	jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,jpeg_out_a60 ,jpeg_out_a61 ,
	jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,jpeg_out_a66 ,jpeg_out_a67 ,
	jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,jpeg_out_a72 ,jpeg_out_a73 ,
	jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,jpeg_out_a78 ,jpeg_out_a79 ,
	jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,jpeg_out_a84 ,jpeg_out_a85 ,
	jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,jpeg_out_a90 ,jpeg_out_a91 ,
	jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,jpeg_out_a96 ,jpeg_out_a97 ,
	jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,jpeg_out_a102 ,
	jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,jpeg_out_a107 ,
	jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,jpeg_out_a112 ,
	jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,jpeg_out_a117 ,
	jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,jpeg_out_a122 ,
	jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,jpeg_out_a127 ,
	jpeg_len_out ,valid );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a64 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a65 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a66 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a67 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a68 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a69 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a70 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a71 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a72 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a73 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a74 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a75 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a76 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a77 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a78 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a79 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a80 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a81 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a82 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a83 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a84 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a85 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a86 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a87 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a88 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a89 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a90 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a91 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a92 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a93 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a94 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a95 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a96 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a97 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a98 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a99 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a100 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a101 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a102 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a103 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a104 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a105 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a106 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a107 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a108 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a109 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a110 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a111 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a112 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a113 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a114 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a115 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a116 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a117 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a118 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a119 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a120 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a121 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a122 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a123 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a124 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a125 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a126 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a127 ;	// line#=../rle.h:56
input	[11:0]	jpeg_len_in ;	// line#=../rle.h:57
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
wire		ST1_01d ;
wire		ST1_02d ;
wire		ST1_03d ;
wire		ST1_04d ;
wire		ST1_05d ;
wire		ST1_06d ;
wire		ST1_07d ;
wire		ST1_08d ;
wire		ST1_09d ;
wire		ST1_10d ;
wire		ST1_11d ;
wire		ST1_12d ;
wire		ST1_13d ;
wire		ST1_14d ;
wire		ST1_15d ;
wire		ST1_16d ;
wire		ST1_17d ;
wire		ST1_18d ;
wire		ST1_19d ;
wire		ST1_20d ;
wire		ST1_21d ;
wire		ST1_22d ;
wire		ST1_23d ;
wire		ST1_24d ;
wire		ST1_25d ;
wire		ST1_26d ;
wire		ST1_27d ;
wire		ST1_28d ;
wire		ST1_29d ;
wire		ST1_30d ;
wire		ST1_31d ;
wire		ST1_32d ;
wire		ST1_33d ;
wire		ST1_34d ;
wire		ST1_35d ;
wire		ST1_36d ;
wire		ST1_37d ;
wire		ST1_38d ;
wire		ST1_39d ;
wire		ST1_40d ;
wire		ST1_41d ;
wire		ST1_42d ;
wire		ST1_43d ;
wire		ST1_44d ;
wire		ST1_45d ;
wire		ST1_46d ;
wire		ST1_47d ;
wire		ST1_48d ;
wire		ST1_49d ;
wire		ST1_50d ;
wire		ST1_51d ;
wire		ST1_52d ;
wire		ST1_53d ;
wire		ST1_54d ;
wire		JF_01 ;
wire		lop8u_11ot ;
wire		JF_03 ;
wire		CT_30 ;
wire		CT_35 ;
wire		JF_06 ;
wire		FL01_01_Leos_all ;

jpeg_fsm INST_fsm ( .clk(clk) ,.rst(rst) ,.ST1_54d(ST1_54d) ,.ST1_53d(ST1_53d) ,
	.ST1_52d(ST1_52d) ,.ST1_51d(ST1_51d) ,.ST1_50d(ST1_50d) ,.ST1_49d(ST1_49d) ,
	.ST1_48d(ST1_48d) ,.ST1_47d(ST1_47d) ,.ST1_46d(ST1_46d) ,.ST1_45d(ST1_45d) ,
	.ST1_44d(ST1_44d) ,.ST1_43d(ST1_43d) ,.ST1_42d(ST1_42d) ,.ST1_41d(ST1_41d) ,
	.ST1_40d(ST1_40d) ,.ST1_39d(ST1_39d) ,.ST1_38d(ST1_38d) ,.ST1_37d(ST1_37d) ,
	.ST1_36d(ST1_36d) ,.ST1_35d(ST1_35d) ,.ST1_34d(ST1_34d) ,.ST1_33d(ST1_33d) ,
	.ST1_32d(ST1_32d) ,.ST1_31d(ST1_31d) ,.ST1_30d(ST1_30d) ,.ST1_29d(ST1_29d) ,
	.ST1_28d(ST1_28d) ,.ST1_27d(ST1_27d) ,.ST1_26d(ST1_26d) ,.ST1_25d(ST1_25d) ,
	.ST1_24d(ST1_24d) ,.ST1_23d(ST1_23d) ,.ST1_22d(ST1_22d) ,.ST1_21d(ST1_21d) ,
	.ST1_20d(ST1_20d) ,.ST1_19d(ST1_19d) ,.ST1_18d(ST1_18d) ,.ST1_17d(ST1_17d) ,
	.ST1_16d(ST1_16d) ,.ST1_15d(ST1_15d) ,.ST1_14d(ST1_14d) ,.ST1_13d(ST1_13d) ,
	.ST1_12d(ST1_12d) ,.ST1_11d(ST1_11d) ,.ST1_10d(ST1_10d) ,.ST1_09d(ST1_09d) ,
	.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,
	.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,
	.JF_01(JF_01) ,.lop8u_11ot(lop8u_11ot) ,.JF_03(JF_03) ,.CT_30(CT_30) ,.CT_35(CT_35) ,
	.JF_06(JF_06) ,.FL01_01_Leos_all(FL01_01_Leos_all) );
jpeg_dat INST_dat ( .clk(clk) ,.rst(rst) ,.jpeg_in_a00(jpeg_in_a00) ,.jpeg_in_a01(jpeg_in_a01) ,
	.jpeg_in_a02(jpeg_in_a02) ,.jpeg_in_a03(jpeg_in_a03) ,.jpeg_in_a04(jpeg_in_a04) ,
	.jpeg_in_a05(jpeg_in_a05) ,.jpeg_in_a06(jpeg_in_a06) ,.jpeg_in_a07(jpeg_in_a07) ,
	.jpeg_in_a08(jpeg_in_a08) ,.jpeg_in_a09(jpeg_in_a09) ,.jpeg_in_a10(jpeg_in_a10) ,
	.jpeg_in_a11(jpeg_in_a11) ,.jpeg_in_a12(jpeg_in_a12) ,.jpeg_in_a13(jpeg_in_a13) ,
	.jpeg_in_a14(jpeg_in_a14) ,.jpeg_in_a15(jpeg_in_a15) ,.jpeg_in_a16(jpeg_in_a16) ,
	.jpeg_in_a17(jpeg_in_a17) ,.jpeg_in_a18(jpeg_in_a18) ,.jpeg_in_a19(jpeg_in_a19) ,
	.jpeg_in_a20(jpeg_in_a20) ,.jpeg_in_a21(jpeg_in_a21) ,.jpeg_in_a22(jpeg_in_a22) ,
	.jpeg_in_a23(jpeg_in_a23) ,.jpeg_in_a24(jpeg_in_a24) ,.jpeg_in_a25(jpeg_in_a25) ,
	.jpeg_in_a26(jpeg_in_a26) ,.jpeg_in_a27(jpeg_in_a27) ,.jpeg_in_a28(jpeg_in_a28) ,
	.jpeg_in_a29(jpeg_in_a29) ,.jpeg_in_a30(jpeg_in_a30) ,.jpeg_in_a31(jpeg_in_a31) ,
	.jpeg_in_a32(jpeg_in_a32) ,.jpeg_in_a33(jpeg_in_a33) ,.jpeg_in_a34(jpeg_in_a34) ,
	.jpeg_in_a35(jpeg_in_a35) ,.jpeg_in_a36(jpeg_in_a36) ,.jpeg_in_a37(jpeg_in_a37) ,
	.jpeg_in_a38(jpeg_in_a38) ,.jpeg_in_a39(jpeg_in_a39) ,.jpeg_in_a40(jpeg_in_a40) ,
	.jpeg_in_a41(jpeg_in_a41) ,.jpeg_in_a42(jpeg_in_a42) ,.jpeg_in_a43(jpeg_in_a43) ,
	.jpeg_in_a44(jpeg_in_a44) ,.jpeg_in_a45(jpeg_in_a45) ,.jpeg_in_a46(jpeg_in_a46) ,
	.jpeg_in_a47(jpeg_in_a47) ,.jpeg_in_a48(jpeg_in_a48) ,.jpeg_in_a49(jpeg_in_a49) ,
	.jpeg_in_a50(jpeg_in_a50) ,.jpeg_in_a51(jpeg_in_a51) ,.jpeg_in_a52(jpeg_in_a52) ,
	.jpeg_in_a53(jpeg_in_a53) ,.jpeg_in_a54(jpeg_in_a54) ,.jpeg_in_a55(jpeg_in_a55) ,
	.jpeg_in_a56(jpeg_in_a56) ,.jpeg_in_a57(jpeg_in_a57) ,.jpeg_in_a58(jpeg_in_a58) ,
	.jpeg_in_a59(jpeg_in_a59) ,.jpeg_in_a60(jpeg_in_a60) ,.jpeg_in_a61(jpeg_in_a61) ,
	.jpeg_in_a62(jpeg_in_a62) ,.jpeg_in_a63(jpeg_in_a63) ,.jpeg_out_a00(jpeg_out_a00) ,
	.jpeg_out_a01(jpeg_out_a01) ,.jpeg_out_a02(jpeg_out_a02) ,.jpeg_out_a03(jpeg_out_a03) ,
	.jpeg_out_a04(jpeg_out_a04) ,.jpeg_out_a05(jpeg_out_a05) ,.jpeg_out_a06(jpeg_out_a06) ,
	.jpeg_out_a07(jpeg_out_a07) ,.jpeg_out_a08(jpeg_out_a08) ,.jpeg_out_a09(jpeg_out_a09) ,
	.jpeg_out_a10(jpeg_out_a10) ,.jpeg_out_a11(jpeg_out_a11) ,.jpeg_out_a12(jpeg_out_a12) ,
	.jpeg_out_a13(jpeg_out_a13) ,.jpeg_out_a14(jpeg_out_a14) ,.jpeg_out_a15(jpeg_out_a15) ,
	.jpeg_out_a16(jpeg_out_a16) ,.jpeg_out_a17(jpeg_out_a17) ,.jpeg_out_a18(jpeg_out_a18) ,
	.jpeg_out_a19(jpeg_out_a19) ,.jpeg_out_a20(jpeg_out_a20) ,.jpeg_out_a21(jpeg_out_a21) ,
	.jpeg_out_a22(jpeg_out_a22) ,.jpeg_out_a23(jpeg_out_a23) ,.jpeg_out_a24(jpeg_out_a24) ,
	.jpeg_out_a25(jpeg_out_a25) ,.jpeg_out_a26(jpeg_out_a26) ,.jpeg_out_a27(jpeg_out_a27) ,
	.jpeg_out_a28(jpeg_out_a28) ,.jpeg_out_a29(jpeg_out_a29) ,.jpeg_out_a30(jpeg_out_a30) ,
	.jpeg_out_a31(jpeg_out_a31) ,.jpeg_out_a32(jpeg_out_a32) ,.jpeg_out_a33(jpeg_out_a33) ,
	.jpeg_out_a34(jpeg_out_a34) ,.jpeg_out_a35(jpeg_out_a35) ,.jpeg_out_a36(jpeg_out_a36) ,
	.jpeg_out_a37(jpeg_out_a37) ,.jpeg_out_a38(jpeg_out_a38) ,.jpeg_out_a39(jpeg_out_a39) ,
	.jpeg_out_a40(jpeg_out_a40) ,.jpeg_out_a41(jpeg_out_a41) ,.jpeg_out_a42(jpeg_out_a42) ,
	.jpeg_out_a43(jpeg_out_a43) ,.jpeg_out_a44(jpeg_out_a44) ,.jpeg_out_a45(jpeg_out_a45) ,
	.jpeg_out_a46(jpeg_out_a46) ,.jpeg_out_a47(jpeg_out_a47) ,.jpeg_out_a48(jpeg_out_a48) ,
	.jpeg_out_a49(jpeg_out_a49) ,.jpeg_out_a50(jpeg_out_a50) ,.jpeg_out_a51(jpeg_out_a51) ,
	.jpeg_out_a52(jpeg_out_a52) ,.jpeg_out_a53(jpeg_out_a53) ,.jpeg_out_a54(jpeg_out_a54) ,
	.jpeg_out_a55(jpeg_out_a55) ,.jpeg_out_a56(jpeg_out_a56) ,.jpeg_out_a57(jpeg_out_a57) ,
	.jpeg_out_a58(jpeg_out_a58) ,.jpeg_out_a59(jpeg_out_a59) ,.jpeg_out_a60(jpeg_out_a60) ,
	.jpeg_out_a61(jpeg_out_a61) ,.jpeg_out_a62(jpeg_out_a62) ,.jpeg_out_a63(jpeg_out_a63) ,
	.jpeg_out_a64(jpeg_out_a64) ,.jpeg_out_a65(jpeg_out_a65) ,.jpeg_out_a66(jpeg_out_a66) ,
	.jpeg_out_a67(jpeg_out_a67) ,.jpeg_out_a68(jpeg_out_a68) ,.jpeg_out_a69(jpeg_out_a69) ,
	.jpeg_out_a70(jpeg_out_a70) ,.jpeg_out_a71(jpeg_out_a71) ,.jpeg_out_a72(jpeg_out_a72) ,
	.jpeg_out_a73(jpeg_out_a73) ,.jpeg_out_a74(jpeg_out_a74) ,.jpeg_out_a75(jpeg_out_a75) ,
	.jpeg_out_a76(jpeg_out_a76) ,.jpeg_out_a77(jpeg_out_a77) ,.jpeg_out_a78(jpeg_out_a78) ,
	.jpeg_out_a79(jpeg_out_a79) ,.jpeg_out_a80(jpeg_out_a80) ,.jpeg_out_a81(jpeg_out_a81) ,
	.jpeg_out_a82(jpeg_out_a82) ,.jpeg_out_a83(jpeg_out_a83) ,.jpeg_out_a84(jpeg_out_a84) ,
	.jpeg_out_a85(jpeg_out_a85) ,.jpeg_out_a86(jpeg_out_a86) ,.jpeg_out_a87(jpeg_out_a87) ,
	.jpeg_out_a88(jpeg_out_a88) ,.jpeg_out_a89(jpeg_out_a89) ,.jpeg_out_a90(jpeg_out_a90) ,
	.jpeg_out_a91(jpeg_out_a91) ,.jpeg_out_a92(jpeg_out_a92) ,.jpeg_out_a93(jpeg_out_a93) ,
	.jpeg_out_a94(jpeg_out_a94) ,.jpeg_out_a95(jpeg_out_a95) ,.jpeg_out_a96(jpeg_out_a96) ,
	.jpeg_out_a97(jpeg_out_a97) ,.jpeg_out_a98(jpeg_out_a98) ,.jpeg_out_a99(jpeg_out_a99) ,
	.jpeg_out_a100(jpeg_out_a100) ,.jpeg_out_a101(jpeg_out_a101) ,.jpeg_out_a102(jpeg_out_a102) ,
	.jpeg_out_a103(jpeg_out_a103) ,.jpeg_out_a104(jpeg_out_a104) ,.jpeg_out_a105(jpeg_out_a105) ,
	.jpeg_out_a106(jpeg_out_a106) ,.jpeg_out_a107(jpeg_out_a107) ,.jpeg_out_a108(jpeg_out_a108) ,
	.jpeg_out_a109(jpeg_out_a109) ,.jpeg_out_a110(jpeg_out_a110) ,.jpeg_out_a111(jpeg_out_a111) ,
	.jpeg_out_a112(jpeg_out_a112) ,.jpeg_out_a113(jpeg_out_a113) ,.jpeg_out_a114(jpeg_out_a114) ,
	.jpeg_out_a115(jpeg_out_a115) ,.jpeg_out_a116(jpeg_out_a116) ,.jpeg_out_a117(jpeg_out_a117) ,
	.jpeg_out_a118(jpeg_out_a118) ,.jpeg_out_a119(jpeg_out_a119) ,.jpeg_out_a120(jpeg_out_a120) ,
	.jpeg_out_a121(jpeg_out_a121) ,.jpeg_out_a122(jpeg_out_a122) ,.jpeg_out_a123(jpeg_out_a123) ,
	.jpeg_out_a124(jpeg_out_a124) ,.jpeg_out_a125(jpeg_out_a125) ,.jpeg_out_a126(jpeg_out_a126) ,
	.jpeg_out_a127(jpeg_out_a127) ,.jpeg_len_out(jpeg_len_out) ,.valid(valid) ,
	.ST1_54d(ST1_54d) ,.ST1_53d(ST1_53d) ,.ST1_52d(ST1_52d) ,.ST1_51d(ST1_51d) ,
	.ST1_50d(ST1_50d) ,.ST1_49d(ST1_49d) ,.ST1_48d(ST1_48d) ,.ST1_47d(ST1_47d) ,
	.ST1_46d(ST1_46d) ,.ST1_45d(ST1_45d) ,.ST1_44d(ST1_44d) ,.ST1_43d(ST1_43d) ,
	.ST1_42d(ST1_42d) ,.ST1_41d(ST1_41d) ,.ST1_40d(ST1_40d) ,.ST1_39d(ST1_39d) ,
	.ST1_38d(ST1_38d) ,.ST1_37d(ST1_37d) ,.ST1_36d(ST1_36d) ,.ST1_35d(ST1_35d) ,
	.ST1_34d(ST1_34d) ,.ST1_33d(ST1_33d) ,.ST1_32d(ST1_32d) ,.ST1_31d(ST1_31d) ,
	.ST1_30d(ST1_30d) ,.ST1_29d(ST1_29d) ,.ST1_28d(ST1_28d) ,.ST1_27d(ST1_27d) ,
	.ST1_26d(ST1_26d) ,.ST1_25d(ST1_25d) ,.ST1_24d(ST1_24d) ,.ST1_23d(ST1_23d) ,
	.ST1_22d(ST1_22d) ,.ST1_21d(ST1_21d) ,.ST1_20d(ST1_20d) ,.ST1_19d(ST1_19d) ,
	.ST1_18d(ST1_18d) ,.ST1_17d(ST1_17d) ,.ST1_16d(ST1_16d) ,.ST1_15d(ST1_15d) ,
	.ST1_14d(ST1_14d) ,.ST1_13d(ST1_13d) ,.ST1_12d(ST1_12d) ,.ST1_11d(ST1_11d) ,
	.ST1_10d(ST1_10d) ,.ST1_09d(ST1_09d) ,.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,
	.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,
	.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,.JF_01(JF_01) ,.lop8u_11ot_port(lop8u_11ot) ,
	.JF_03(JF_03) ,.CT_30_port(CT_30) ,.CT_35_port(CT_35) ,.JF_06_port(JF_06) ,
	.FL01_01_Leos_all(FL01_01_Leos_all) );

endmodule

module jpeg_fsm ( clk ,rst ,ST1_54d ,ST1_53d ,ST1_52d ,ST1_51d ,ST1_50d ,ST1_49d ,
	ST1_48d ,ST1_47d ,ST1_46d ,ST1_45d ,ST1_44d ,ST1_43d ,ST1_42d ,ST1_41d ,
	ST1_40d ,ST1_39d ,ST1_38d ,ST1_37d ,ST1_36d ,ST1_35d ,ST1_34d ,ST1_33d ,
	ST1_32d ,ST1_31d ,ST1_30d ,ST1_29d ,ST1_28d ,ST1_27d ,ST1_26d ,ST1_25d ,
	ST1_24d ,ST1_23d ,ST1_22d ,ST1_21d ,ST1_20d ,ST1_19d ,ST1_18d ,ST1_17d ,
	ST1_16d ,ST1_15d ,ST1_14d ,ST1_13d ,ST1_12d ,ST1_11d ,ST1_10d ,ST1_09d ,
	ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,ST1_02d ,ST1_01d ,
	JF_01 ,lop8u_11ot ,JF_03 ,CT_30 ,CT_35 ,JF_06 ,FL01_01_Leos_all );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
output		ST1_54d ;
output		ST1_53d ;
output		ST1_52d ;
output		ST1_51d ;
output		ST1_50d ;
output		ST1_49d ;
output		ST1_48d ;
output		ST1_47d ;
output		ST1_46d ;
output		ST1_45d ;
output		ST1_44d ;
output		ST1_43d ;
output		ST1_42d ;
output		ST1_41d ;
output		ST1_40d ;
output		ST1_39d ;
output		ST1_38d ;
output		ST1_37d ;
output		ST1_36d ;
output		ST1_35d ;
output		ST1_34d ;
output		ST1_33d ;
output		ST1_32d ;
output		ST1_31d ;
output		ST1_30d ;
output		ST1_29d ;
output		ST1_28d ;
output		ST1_27d ;
output		ST1_26d ;
output		ST1_25d ;
output		ST1_24d ;
output		ST1_23d ;
output		ST1_22d ;
output		ST1_21d ;
output		ST1_20d ;
output		ST1_19d ;
output		ST1_18d ;
output		ST1_17d ;
output		ST1_16d ;
output		ST1_15d ;
output		ST1_14d ;
output		ST1_13d ;
output		ST1_12d ;
output		ST1_11d ;
output		ST1_10d ;
output		ST1_09d ;
output		ST1_08d ;
output		ST1_07d ;
output		ST1_06d ;
output		ST1_05d ;
output		ST1_04d ;
output		ST1_03d ;
output		ST1_02d ;
output		ST1_01d ;
input		JF_01 ;
input		lop8u_11ot ;
input		JF_03 ;
input		CT_30 ;
input		CT_35 ;
input		JF_06 ;
input		FL01_01_Leos_all ;
reg	[5:0]	B01_streg ;

parameter	ST1_01 = 6'h00 ;
parameter	ST1_02 = 6'h01 ;
parameter	ST1_03 = 6'h02 ;
parameter	ST1_04 = 6'h03 ;
parameter	ST1_05 = 6'h04 ;
parameter	ST1_06 = 6'h05 ;
parameter	ST1_07 = 6'h06 ;
parameter	ST1_08 = 6'h07 ;
parameter	ST1_09 = 6'h08 ;
parameter	ST1_10 = 6'h09 ;
parameter	ST1_11 = 6'h0a ;
parameter	ST1_12 = 6'h0b ;
parameter	ST1_13 = 6'h0c ;
parameter	ST1_14 = 6'h0d ;
parameter	ST1_15 = 6'h0e ;
parameter	ST1_16 = 6'h0f ;
parameter	ST1_17 = 6'h10 ;
parameter	ST1_18 = 6'h11 ;
parameter	ST1_19 = 6'h12 ;
parameter	ST1_20 = 6'h13 ;
parameter	ST1_21 = 6'h14 ;
parameter	ST1_22 = 6'h15 ;
parameter	ST1_23 = 6'h16 ;
parameter	ST1_24 = 6'h17 ;
parameter	ST1_25 = 6'h18 ;
parameter	ST1_26 = 6'h19 ;
parameter	ST1_27 = 6'h1a ;
parameter	ST1_28 = 6'h1b ;
parameter	ST1_29 = 6'h1c ;
parameter	ST1_30 = 6'h1d ;
parameter	ST1_31 = 6'h1e ;
parameter	ST1_32 = 6'h1f ;
parameter	ST1_33 = 6'h20 ;
parameter	ST1_34 = 6'h21 ;
parameter	ST1_35 = 6'h22 ;
parameter	ST1_36 = 6'h23 ;
parameter	ST1_37 = 6'h24 ;
parameter	ST1_38 = 6'h25 ;
parameter	ST1_39 = 6'h26 ;
parameter	ST1_40 = 6'h27 ;
parameter	ST1_41 = 6'h28 ;
parameter	ST1_42 = 6'h29 ;
parameter	ST1_43 = 6'h2a ;
parameter	ST1_44 = 6'h2b ;
parameter	ST1_45 = 6'h2c ;
parameter	ST1_46 = 6'h2d ;
parameter	ST1_47 = 6'h2e ;
parameter	ST1_48 = 6'h2f ;
parameter	ST1_49 = 6'h30 ;
parameter	ST1_50 = 6'h31 ;
parameter	ST1_51 = 6'h32 ;
parameter	ST1_52 = 6'h33 ;
parameter	ST1_53 = 6'h34 ;
parameter	ST1_54 = 6'h35 ;

assign	ST1_01d = ( ( B01_streg == ST1_01 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_02d = ( ( B01_streg == ST1_02 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_03d = ( ( B01_streg == ST1_03 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_04d = ( ( B01_streg == ST1_04 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_05d = ( ( B01_streg == ST1_05 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_06d = ( ( B01_streg == ST1_06 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_07d = ( ( B01_streg == ST1_07 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_08d = ( ( B01_streg == ST1_08 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_09d = ( ( B01_streg == ST1_09 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_10d = ( ( B01_streg == ST1_10 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_11d = ( ( B01_streg == ST1_11 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_12d = ( ( B01_streg == ST1_12 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_13d = ( ( B01_streg == ST1_13 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_14d = ( ( B01_streg == ST1_14 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_15d = ( ( B01_streg == ST1_15 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_16d = ( ( B01_streg == ST1_16 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_17d = ( ( B01_streg == ST1_17 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_18d = ( ( B01_streg == ST1_18 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_19d = ( ( B01_streg == ST1_19 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_20d = ( ( B01_streg == ST1_20 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_21d = ( ( B01_streg == ST1_21 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_22d = ( ( B01_streg == ST1_22 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_23d = ( ( B01_streg == ST1_23 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_24d = ( ( B01_streg == ST1_24 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_25d = ( ( B01_streg == ST1_25 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_26d = ( ( B01_streg == ST1_26 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_27d = ( ( B01_streg == ST1_27 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_28d = ( ( B01_streg == ST1_28 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_29d = ( ( B01_streg == ST1_29 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_30d = ( ( B01_streg == ST1_30 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_31d = ( ( B01_streg == ST1_31 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_32d = ( ( B01_streg == ST1_32 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_33d = ( ( B01_streg == ST1_33 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_34d = ( ( B01_streg == ST1_34 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_35d = ( ( B01_streg == ST1_35 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_36d = ( ( B01_streg == ST1_36 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_37d = ( ( B01_streg == ST1_37 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_38d = ( ( B01_streg == ST1_38 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_39d = ( ( B01_streg == ST1_39 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_40d = ( ( B01_streg == ST1_40 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_41d = ( ( B01_streg == ST1_41 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_42d = ( ( B01_streg == ST1_42 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_43d = ( ( B01_streg == ST1_43 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_44d = ( ( B01_streg == ST1_44 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_45d = ( ( B01_streg == ST1_45 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_46d = ( ( B01_streg == ST1_46 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_47d = ( ( B01_streg == ST1_47 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_48d = ( ( B01_streg == ST1_48 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_49d = ( ( B01_streg == ST1_49 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_50d = ( ( B01_streg == ST1_50 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_51d = ( ( B01_streg == ST1_51 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_52d = ( ( B01_streg == ST1_52 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_53d = ( ( B01_streg == ST1_53 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_54d = ( ( B01_streg == ST1_54 ) ? 1'h1 : 1'h0 ) ;
always @ ( posedge clk )
	if ( !rst )
		B01_streg <= ST1_01 ;
	else
		case ( B01_streg )
		ST1_01 :
			B01_streg <= ST1_02 ;
		ST1_02 :
			if ( ( JF_01 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_03 ;
		ST1_03 :
			if ( ( lop8u_11ot != 1'h0 ) )
				B01_streg <= ST1_03 ;
			else
				B01_streg <= ST1_04 ;
		ST1_04 :
			if ( ( JF_03 != 1'h0 ) )
				B01_streg <= ST1_04 ;
			else
				B01_streg <= ST1_05 ;
		ST1_05 :
			if ( ( CT_30 != 1'h0 ) )
				B01_streg <= ST1_05 ;
			else
				B01_streg <= ST1_06 ;
		ST1_06 :
			B01_streg <= ST1_07 ;
		ST1_07 :
			if ( ( CT_35 != 1'h0 ) )
				B01_streg <= ST1_05 ;
			else
				B01_streg <= ST1_08 ;
		ST1_08 :
			B01_streg <= ST1_09 ;
		ST1_09 :
			if ( ( JF_06 != 1'h0 ) )
				B01_streg <= ST1_10 ;
			else
				B01_streg <= ST1_11 ;
		ST1_10 :
			B01_streg <= ST1_11 ;
		ST1_11 :
			if ( ( FL01_01_Leos_all != 1'h0 ) )
				B01_streg <= ST1_12 ;
			else
				B01_streg <= ST1_11 ;
		ST1_12 :
			B01_streg <= ST1_13 ;
		ST1_13 :
			B01_streg <= ST1_14 ;
		ST1_14 :
			B01_streg <= ST1_15 ;
		ST1_15 :
			B01_streg <= ST1_16 ;
		ST1_16 :
			B01_streg <= ST1_17 ;
		ST1_17 :
			B01_streg <= ST1_18 ;
		ST1_18 :
			B01_streg <= ST1_19 ;
		ST1_19 :
			B01_streg <= ST1_20 ;
		ST1_20 :
			B01_streg <= ST1_21 ;
		ST1_21 :
			B01_streg <= ST1_22 ;
		ST1_22 :
			B01_streg <= ST1_23 ;
		ST1_23 :
			B01_streg <= ST1_24 ;
		ST1_24 :
			B01_streg <= ST1_25 ;
		ST1_25 :
			B01_streg <= ST1_26 ;
		ST1_26 :
			B01_streg <= ST1_27 ;
		ST1_27 :
			B01_streg <= ST1_28 ;
		ST1_28 :
			B01_streg <= ST1_29 ;
		ST1_29 :
			B01_streg <= ST1_30 ;
		ST1_30 :
			B01_streg <= ST1_31 ;
		ST1_31 :
			B01_streg <= ST1_32 ;
		ST1_32 :
			B01_streg <= ST1_33 ;
		ST1_33 :
			B01_streg <= ST1_34 ;
		ST1_34 :
			B01_streg <= ST1_35 ;
		ST1_35 :
			B01_streg <= ST1_36 ;
		ST1_36 :
			B01_streg <= ST1_37 ;
		ST1_37 :
			B01_streg <= ST1_38 ;
		ST1_38 :
			B01_streg <= ST1_39 ;
		ST1_39 :
			B01_streg <= ST1_40 ;
		ST1_40 :
			B01_streg <= ST1_41 ;
		ST1_41 :
			B01_streg <= ST1_42 ;
		ST1_42 :
			B01_streg <= ST1_43 ;
		ST1_43 :
			B01_streg <= ST1_44 ;
		ST1_44 :
			B01_streg <= ST1_45 ;
		ST1_45 :
			B01_streg <= ST1_46 ;
		ST1_46 :
			B01_streg <= ST1_47 ;
		ST1_47 :
			B01_streg <= ST1_48 ;
		ST1_48 :
			B01_streg <= ST1_49 ;
		ST1_49 :
			B01_streg <= ST1_50 ;
		ST1_50 :
			B01_streg <= ST1_51 ;
		ST1_51 :
			B01_streg <= ST1_52 ;
		ST1_52 :
			B01_streg <= ST1_53 ;
		ST1_53 :
			B01_streg <= ST1_54 ;
		ST1_54 :
			B01_streg <= ST1_02 ;
		default :
			B01_streg <= ST1_01 ;
		endcase

endmodule

module jpeg_dat ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,
	jpeg_in_a04 ,jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,
	jpeg_in_a10 ,jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,
	jpeg_in_a16 ,jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,
	jpeg_in_a22 ,jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,
	jpeg_in_a28 ,jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,
	jpeg_in_a34 ,jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,
	jpeg_in_a40 ,jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,
	jpeg_in_a46 ,jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,
	jpeg_in_a52 ,jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,
	jpeg_in_a58 ,jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,
	jpeg_out_a00 ,jpeg_out_a01 ,jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,
	jpeg_out_a06 ,jpeg_out_a07 ,jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,
	jpeg_out_a12 ,jpeg_out_a13 ,jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,
	jpeg_out_a18 ,jpeg_out_a19 ,jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,
	jpeg_out_a24 ,jpeg_out_a25 ,jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,
	jpeg_out_a30 ,jpeg_out_a31 ,jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,
	jpeg_out_a36 ,jpeg_out_a37 ,jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,
	jpeg_out_a42 ,jpeg_out_a43 ,jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,
	jpeg_out_a48 ,jpeg_out_a49 ,jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,
	jpeg_out_a54 ,jpeg_out_a55 ,jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,
	jpeg_out_a60 ,jpeg_out_a61 ,jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,
	jpeg_out_a66 ,jpeg_out_a67 ,jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,
	jpeg_out_a72 ,jpeg_out_a73 ,jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,
	jpeg_out_a78 ,jpeg_out_a79 ,jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,
	jpeg_out_a84 ,jpeg_out_a85 ,jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,
	jpeg_out_a90 ,jpeg_out_a91 ,jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,
	jpeg_out_a96 ,jpeg_out_a97 ,jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,
	jpeg_out_a102 ,jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,
	jpeg_out_a107 ,jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,
	jpeg_out_a112 ,jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,
	jpeg_out_a117 ,jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,
	jpeg_out_a122 ,jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,
	jpeg_out_a127 ,jpeg_len_out ,valid ,ST1_54d ,ST1_53d ,ST1_52d ,ST1_51d ,
	ST1_50d ,ST1_49d ,ST1_48d ,ST1_47d ,ST1_46d ,ST1_45d ,ST1_44d ,ST1_43d ,
	ST1_42d ,ST1_41d ,ST1_40d ,ST1_39d ,ST1_38d ,ST1_37d ,ST1_36d ,ST1_35d ,
	ST1_34d ,ST1_33d ,ST1_32d ,ST1_31d ,ST1_30d ,ST1_29d ,ST1_28d ,ST1_27d ,
	ST1_26d ,ST1_25d ,ST1_24d ,ST1_23d ,ST1_22d ,ST1_21d ,ST1_20d ,ST1_19d ,
	ST1_18d ,ST1_17d ,ST1_16d ,ST1_15d ,ST1_14d ,ST1_13d ,ST1_12d ,ST1_11d ,
	ST1_10d ,ST1_09d ,ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,
	ST1_02d ,ST1_01d ,JF_01 ,lop8u_11ot_port ,JF_03 ,CT_30_port ,CT_35_port ,
	JF_06_port ,FL01_01_Leos_all );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
input		ST1_54d ;
input		ST1_53d ;
input		ST1_52d ;
input		ST1_51d ;
input		ST1_50d ;
input		ST1_49d ;
input		ST1_48d ;
input		ST1_47d ;
input		ST1_46d ;
input		ST1_45d ;
input		ST1_44d ;
input		ST1_43d ;
input		ST1_42d ;
input		ST1_41d ;
input		ST1_40d ;
input		ST1_39d ;
input		ST1_38d ;
input		ST1_37d ;
input		ST1_36d ;
input		ST1_35d ;
input		ST1_34d ;
input		ST1_33d ;
input		ST1_32d ;
input		ST1_31d ;
input		ST1_30d ;
input		ST1_29d ;
input		ST1_28d ;
input		ST1_27d ;
input		ST1_26d ;
input		ST1_25d ;
input		ST1_24d ;
input		ST1_23d ;
input		ST1_22d ;
input		ST1_21d ;
input		ST1_20d ;
input		ST1_19d ;
input		ST1_18d ;
input		ST1_17d ;
input		ST1_16d ;
input		ST1_15d ;
input		ST1_14d ;
input		ST1_13d ;
input		ST1_12d ;
input		ST1_11d ;
input		ST1_10d ;
input		ST1_09d ;
input		ST1_08d ;
input		ST1_07d ;
input		ST1_06d ;
input		ST1_05d ;
input		ST1_04d ;
input		ST1_03d ;
input		ST1_02d ;
input		ST1_01d ;
output		JF_01 ;
output		lop8u_11ot_port ;
output		JF_03 ;
output		CT_30_port ;
output		CT_35_port ;
output		JF_06_port ;
output		FL01_01_Leos_all ;
wire		M_219 ;
wire		M_216 ;
wire		M_215 ;
wire		M_213 ;
wire		M_212 ;
wire		M_211 ;
wire		M_210 ;
wire		M_209 ;
wire		M_208 ;
wire		M_207 ;
wire		M_206 ;
wire		M_205 ;
wire		M_204 ;
wire		M_203 ;
wire		M_202 ;
wire		M_201 ;
wire		M_200 ;
wire		M_199 ;
wire		M_198 ;
wire		M_197 ;
wire		M_196 ;
wire		M_195 ;
wire		M_194 ;
wire		M_193 ;
wire		M_192 ;
wire		M_191 ;
wire		M_190 ;
wire		M_189 ;
wire		M_188 ;
wire		M_186 ;
wire		M_185 ;
wire		M_184 ;
wire		M_183 ;
wire		M_182 ;
wire		M_181 ;
wire		M_180 ;
wire		M_179 ;
wire		M_178 ;
wire		M_177 ;
wire		M_176 ;
wire		M_175 ;
wire		M_174 ;
wire		M_173 ;
wire		M_172 ;
wire		M_171 ;
wire		M_170 ;
wire		M_169 ;
wire		M_168 ;
wire		M_167 ;
wire		M_166 ;
wire		M_165 ;
wire		M_164 ;
wire		M_163 ;
wire		M_162 ;
wire		M_161 ;
wire		M_160 ;
wire		M_159 ;
wire		M_158 ;
wire		M_157 ;
wire		M_156 ;
wire		M_155 ;
wire		M_154 ;
wire		M_153 ;
wire		M_152 ;
wire		M_151 ;
wire		M_150 ;
wire		M_149 ;
wire		M_148 ;
wire		M_147 ;
wire		M_146 ;
wire		M_145 ;
wire		M_144 ;
wire		M_143 ;
wire		M_142 ;
wire		M_141 ;
wire		M_140 ;
wire		M_139 ;
wire		M_138 ;
wire		M_137 ;
wire		M_136 ;
wire		M_135 ;
wire		M_134 ;
wire		M_133 ;
wire		M_132 ;
wire		M_131 ;
wire		M_130 ;
wire		M_128 ;
wire		M_126 ;
wire		M_124 ;
wire		M_122 ;
wire		M_120 ;
wire		M_118 ;
wire		M_116 ;
wire		M_115 ;
wire		M_114 ;
wire		M_110 ;
wire		M_107 ;
wire		M_106 ;
wire		U_280 ;
wire		U_278 ;
wire		U_273 ;
wire		U_269 ;
wire		U_268 ;
wire		U_263 ;
wire		U_262 ;
wire		U_257 ;
wire		U_254 ;
wire		U_252 ;
wire		U_251 ;
wire		U_248 ;
wire		U_179 ;
wire		U_178 ;
wire		U_177 ;
wire		U_176 ;
wire		U_175 ;
wire		U_169 ;
wire		U_166 ;
wire		U_165 ;
wire		U_164 ;
wire		U_163 ;
wire		U_162 ;
wire		C_05 ;
wire		U_161 ;
wire		U_88 ;
wire		U_87 ;
wire		U_84 ;
wire		U_83 ;
wire		U_82 ;
wire		U_81 ;
wire		U_80 ;
wire		C_02 ;
wire		U_79 ;
wire		U_06 ;
wire		U_05 ;
wire	[1:0]	sub8u_7_11i2 ;
wire	[6:0]	sub8u_7_11ot ;
wire	[2:0]	sub8u_71i2 ;
wire	[6:0]	sub8u_71i1 ;
wire	[6:0]	sub8u_71ot ;
wire	[31:0]	decr32s2i1 ;
wire	[31:0]	decr32s2ot ;
wire	[31:0]	decr32s1i1 ;
wire	[31:0]	decr32s1ot ;
wire	[6:0]	decr8u_71i1 ;
wire	[6:0]	decr8u_71ot ;
wire	[31:0]	incr32s2i1 ;
wire	[31:0]	incr32s2ot ;
wire	[31:0]	incr32s1i1 ;
wire	[31:0]	incr32s1ot ;
wire	[7:0]	incr8u2ot ;
wire	[7:0]	incr8u1i1 ;
wire	[7:0]	incr8u1ot ;
wire	[3:0]	incr4s1i1 ;
wire	[3:0]	incr4s1ot ;
wire	[5:0]	lop8u_11i2 ;
wire	[5:0]	lop8u_11i1 ;
wire		lop8u_11ot ;
wire	[8:0]	sub12s_91i2 ;
wire	[8:0]	sub12s_91i1 ;
wire	[8:0]	sub12s_91ot ;
wire	[1:0]	sub8u1i2 ;
wire	[7:0]	sub8u1i1 ;
wire	[7:0]	sub8u1ot ;
wire		FL01_02_ndat ;
wire		FL01_01_ndat ;
wire		FL01_03_eos ;
wire		FL01_02_eos ;
wire		FL01_01_eos ;
wire		FL01_01_Leos_all ;
wire		FJ_13_14 ;
wire		FL01_03_01a ;
wire		FL01_02_01a ;
wire		FL01_01_01a ;
wire		FL01_03_break ;
wire		JF_06 ;
wire		CT_35 ;
wire		CT_33 ;
wire		CT_30 ;
wire		CT_18 ;
wire		JF_03 ;
wire		CT_03 ;
wire		JF_01 ;
wire		rl_WE1 ;
wire	[8:0]	rl_RD1 ;
wire	[8:0]	rl_RD3 ;
wire	[8:0]	rl_RD2 ;
wire		RG_previous_dc_en ;
wire		RG_quantized_block_en ;
wire		RG_quantized_block_1_en ;
wire		RG_quantized_block_2_en ;
wire		RG_quantized_block_3_en ;
wire		RG_quantized_block_4_en ;
wire		RG_quantized_block_5_en ;
wire		RG_quantized_block_6_en ;
wire		RG_quantized_block_7_en ;
wire		RG_quantized_block_8_en ;
wire		RG_quantized_block_9_en ;
wire		RG_quantized_block_10_en ;
wire		RG_quantized_block_11_en ;
wire		RG_quantized_block_12_en ;
wire		RG_quantized_block_13_en ;
wire		RG_quantized_block_14_en ;
wire		RG_quantized_block_15_en ;
wire		RG_quantized_block_16_en ;
wire		RG_quantized_block_17_en ;
wire		RG_quantized_block_18_en ;
wire		RG_quantized_block_19_en ;
wire		RG_quantized_block_20_en ;
wire		RG_quantized_block_21_en ;
wire		RG_quantized_block_22_en ;
wire		RG_quantized_block_23_en ;
wire		RG_quantized_block_24_en ;
wire		RG_quantized_block_25_en ;
wire		RG_quantized_block_26_en ;
wire		RG_quantized_block_27_en ;
wire		RG_quantized_block_28_en ;
wire		RG_quantized_block_29_en ;
wire		RG_quantized_block_30_en ;
wire		RG_quantized_block_31_en ;
wire		RG_quantized_block_32_en ;
wire		RG_quantized_block_33_en ;
wire		RG_quantized_block_34_en ;
wire		RG_quantized_block_35_en ;
wire		RG_quantized_block_36_en ;
wire		RG_quantized_block_37_en ;
wire		RG_quantized_block_38_en ;
wire		RG_quantized_block_39_en ;
wire		RG_quantized_block_40_en ;
wire		RG_quantized_block_41_en ;
wire		RG_quantized_block_42_en ;
wire		RG_quantized_block_43_en ;
wire		RG_quantized_block_44_en ;
wire		RG_quantized_block_45_en ;
wire		RG_quantized_block_46_en ;
wire		RG_quantized_block_47_en ;
wire		RG_quantized_block_48_en ;
wire		RG_quantized_block_49_en ;
wire		RG_quantized_block_50_en ;
wire		RG_quantized_block_51_en ;
wire		RG_quantized_block_52_en ;
wire		RG_quantized_block_53_en ;
wire		RG_quantized_block_54_en ;
wire		RG_quantized_block_55_en ;
wire		RG_quantized_block_56_en ;
wire		RG_quantized_block_57_en ;
wire		RG_quantized_block_58_en ;
wire		RG_quantized_block_59_en ;
wire		RG_quantized_block_60_en ;
wire		FF_j_en ;
wire		RG_len_03_en ;
wire		jpeg_out_a00_r_en ;
wire		jpeg_out_a01_r_en ;
wire		jpeg_out_a02_r_en ;
wire		jpeg_out_a03_r_en ;
wire		jpeg_out_a04_r_en ;
wire		jpeg_out_a05_r_en ;
wire		jpeg_out_a06_r_en ;
wire		jpeg_out_a07_r_en ;
wire		jpeg_out_a08_r_en ;
wire		jpeg_out_a09_r_en ;
wire		jpeg_out_a10_r_en ;
wire		jpeg_out_a11_r_en ;
wire		jpeg_out_a12_r_en ;
wire		jpeg_out_a13_r_en ;
wire		jpeg_out_a14_r_en ;
wire		jpeg_out_a15_r_en ;
wire		jpeg_out_a16_r_en ;
wire		jpeg_out_a17_r_en ;
wire		jpeg_out_a18_r_en ;
wire		jpeg_out_a19_r_en ;
wire		jpeg_out_a20_r_en ;
wire		jpeg_out_a21_r_en ;
wire		jpeg_out_a22_r_en ;
wire		jpeg_out_a23_r_en ;
wire		jpeg_out_a24_r_en ;
wire		jpeg_out_a25_r_en ;
wire		jpeg_out_a26_r_en ;
wire		jpeg_out_a27_r_en ;
wire		jpeg_out_a28_r_en ;
wire		jpeg_out_a29_r_en ;
wire		jpeg_out_a30_r_en ;
wire		jpeg_out_a31_r_en ;
wire		jpeg_out_a32_r_en ;
wire		jpeg_out_a33_r_en ;
wire		jpeg_out_a34_r_en ;
wire		jpeg_out_a35_r_en ;
wire		jpeg_out_a36_r_en ;
wire		jpeg_out_a37_r_en ;
wire		jpeg_out_a38_r_en ;
wire		jpeg_out_a39_r_en ;
wire		jpeg_out_a40_r_en ;
wire		jpeg_out_a41_r_en ;
wire		jpeg_out_a42_r_en ;
wire		jpeg_out_a43_r_en ;
wire		jpeg_out_a44_r_en ;
wire		jpeg_out_a45_r_en ;
wire		jpeg_out_a46_r_en ;
wire		jpeg_out_a47_r_en ;
wire		jpeg_out_a48_r_en ;
wire		jpeg_out_a49_r_en ;
wire		jpeg_out_a50_r_en ;
wire		jpeg_out_a51_r_en ;
wire		jpeg_out_a52_r_en ;
wire		jpeg_out_a53_r_en ;
wire		jpeg_out_a54_r_en ;
wire		jpeg_out_a55_r_en ;
wire		jpeg_out_a56_r_en ;
wire		jpeg_out_a57_r_en ;
wire		jpeg_out_a58_r_en ;
wire		jpeg_out_a59_r_en ;
wire		jpeg_out_a60_r_en ;
wire		jpeg_out_a61_r_en ;
wire		jpeg_out_a62_r_en ;
wire		jpeg_out_a63_r_en ;
wire		jpeg_out_a64_r_en ;
wire		jpeg_out_a65_r_en ;
wire		jpeg_out_a66_r_en ;
wire		jpeg_out_a67_r_en ;
wire		jpeg_out_a68_r_en ;
wire		jpeg_out_a69_r_en ;
wire		jpeg_out_a70_r_en ;
wire		jpeg_out_a71_r_en ;
wire		jpeg_out_a72_r_en ;
wire		jpeg_out_a73_r_en ;
wire		jpeg_out_a74_r_en ;
wire		jpeg_out_a75_r_en ;
wire		jpeg_out_a76_r_en ;
wire		jpeg_out_a77_r_en ;
wire		jpeg_out_a78_r_en ;
wire		jpeg_out_a79_r_en ;
wire		jpeg_out_a80_r_en ;
wire		jpeg_out_a81_r_en ;
wire		jpeg_out_a82_r_en ;
wire		jpeg_out_a83_r_en ;
wire		jpeg_out_a84_r_en ;
wire		jpeg_out_a85_r_en ;
wire		jpeg_out_a86_r_en ;
wire		jpeg_out_a87_r_en ;
wire		jpeg_out_a88_r_en ;
wire		jpeg_out_a89_r_en ;
wire		jpeg_out_a90_r_en ;
wire		jpeg_out_a91_r_en ;
wire		jpeg_out_a92_r_en ;
wire		jpeg_out_a93_r_en ;
wire		jpeg_out_a94_r_en ;
wire		jpeg_out_a95_r_en ;
wire		jpeg_out_a96_r_en ;
wire		jpeg_out_a97_r_en ;
wire		jpeg_out_a98_r_en ;
wire		jpeg_out_a99_r_en ;
wire		jpeg_out_a100_r_en ;
wire		jpeg_out_a101_r_en ;
wire		jpeg_out_a102_r_en ;
wire		jpeg_out_a103_r_en ;
wire		jpeg_out_a104_r_en ;
wire		jpeg_out_a105_r_en ;
wire		jpeg_out_a106_r_en ;
wire		jpeg_out_a107_r_en ;
wire		jpeg_out_a108_r_en ;
wire		jpeg_out_a109_r_en ;
wire		jpeg_out_a110_r_en ;
wire		jpeg_out_a111_r_en ;
wire		jpeg_out_a112_r_en ;
wire		jpeg_out_a113_r_en ;
wire		jpeg_out_a114_r_en ;
wire		jpeg_out_a115_r_en ;
wire		jpeg_out_a116_r_en ;
wire		jpeg_out_a117_r_en ;
wire		jpeg_out_a118_r_en ;
wire		jpeg_out_a119_r_en ;
wire		jpeg_out_a120_r_en ;
wire		jpeg_out_a121_r_en ;
wire		jpeg_out_a122_r_en ;
wire		jpeg_out_a123_r_en ;
wire		jpeg_out_a124_r_en ;
wire		jpeg_out_a125_r_en ;
wire		jpeg_out_a126_r_en ;
wire		jpeg_out_a127_r_en ;
wire		jpeg_len_out_r_en ;
wire		RG_previous_dc_zz_en ;
wire		RG_zz_en ;
wire		RG_zz_1_en ;
wire		RG_zz_2_en ;
wire		RG_zz_3_en ;
wire		RG_zz_4_en ;
wire		RG_zz_5_en ;
wire		RG_zz_6_en ;
wire		RG_zz_7_en ;
wire		RG_zz_8_en ;
wire		RG_zz_9_en ;
wire		RG_zz_10_en ;
wire		RG_zz_11_en ;
wire		RG_zz_12_en ;
wire		RG_zz_13_en ;
wire		RG_zz_14_en ;
wire		RG_zz_15_en ;
wire		RG_zz_16_en ;
wire		RG_zz_17_en ;
wire		RG_zz_18_en ;
wire		RG_zz_19_en ;
wire		RG_zz_20_en ;
wire		RG_zz_21_en ;
wire		RG_zz_22_en ;
wire		RG_zz_23_en ;
wire		RG_zz_24_en ;
wire		RG_zz_25_en ;
wire		RG_zz_26_en ;
wire		RG_zz_27_en ;
wire		RG_zz_28_en ;
wire		RG_zz_29_en ;
wire		RG_zz_30_en ;
wire		RG_zz_31_en ;
wire		RG_zz_32_en ;
wire		RG_zz_33_en ;
wire		RG_zz_34_en ;
wire		RG_zz_35_en ;
wire		RG_zz_36_en ;
wire		RG_zz_37_en ;
wire		RG_zz_38_en ;
wire		RG_zz_39_en ;
wire		RG_zz_40_en ;
wire		RG_zz_41_en ;
wire		RG_zz_42_en ;
wire		RG_zz_43_en ;
wire		RG_zz_44_en ;
wire		RG_zz_45_en ;
wire		RG_zz_46_en ;
wire		RG_zz_47_en ;
wire		RG_zz_48_en ;
wire		RG_zz_49_en ;
wire		RG_zz_50_en ;
wire		RG_zz_51_en ;
wire		RG_zz_52_en ;
wire		RG_zz_53_en ;
wire		RG_zz_54_en ;
wire		RG_zz_55_en ;
wire		RG_zz_56_en ;
wire		RG_zz_57_en ;
wire		RG_zz_58_en ;
wire		RG_zz_59_en ;
wire		RG_zz_60_en ;
wire		RG_zz_61_en ;
wire		RG_zz_62_en ;
wire		RG_j_03_en ;
wire		RG_i_en ;
wire		RG_j_k_en ;
wire		RG_quantized_block_rl_02_en ;
wire		RG_quantized_block_rl_02_1_en ;
wire		RG_quantized_block_zz_en ;
wire		FF_d_en ;
wire		FF_i_en ;
wire		FF_len_en ;
wire		RG_len_01_1_en ;
wire		FL01_01_streg_en ;
wire		FL01_02_streg_en ;
wire		FL01_03_streg_en ;
wire		valid_r_en ;
reg	FL01_03_streg ;
reg	FL01_02_streg ;
reg	FL01_01_streg ;
reg	[8:0]	RG_previous_dc ;	// line#=../rle.h:66
reg	[8:0]	RG_previous_dc_zz ;	// line#=../rle.h:65,66
reg	[8:0]	RG_zz ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_1 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_2 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_3 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_4 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_5 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_6 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_7 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_8 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_9 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_10 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_11 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_12 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_13 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_14 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_15 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_16 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_17 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_18 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_19 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_20 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_21 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_22 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_23 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_24 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_25 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_26 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_27 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_28 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_29 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_30 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_31 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_32 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_33 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_34 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_35 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_36 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_37 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_38 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_39 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_40 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_41 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_42 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_43 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_44 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_45 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_46 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_47 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_48 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_49 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_50 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_51 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_52 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_53 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_54 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_55 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_56 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_57 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_58 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_59 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_60 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_61 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_62 ;	// line#=../rle.h:65
reg	[3:0]	RG_j_03 ;	// line#=../rle.cpp:27
reg	[31:0]	RG_i ;	// line#=../rle.cpp:25,105
reg	[31:0]	RG_j_k ;	// line#=../rle.cpp:25,105
reg	[8:0]	RG_quantized_block ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_1 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_2 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_3 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_4 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_5 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_6 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_7 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_8 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_9 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_10 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_11 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_12 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_13 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_14 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_15 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_16 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_17 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_18 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_19 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_20 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_21 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_22 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_23 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_24 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_25 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_26 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_27 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_28 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_29 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_30 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_31 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_32 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_33 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_34 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_35 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_36 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_37 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_38 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_39 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_40 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_41 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_42 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_43 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_44 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_45 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_46 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_47 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_48 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_49 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_50 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_51 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_52 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_53 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_54 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_55 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_56 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_57 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_58 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_59 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_60 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_rl_02 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_02_1 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_zz ;	// line#=../rle.cpp:22 ../rle.h:65
reg	[5:0]	RG_k ;	// line#=../rle.cpp:105
reg	FF_d ;	// line#=../rle.cpp:105
reg	FF_j ;	// line#=../rle.cpp:27
reg	FF_i ;	// line#=../rle.cpp:25
reg	RG_136 ;
reg	FF_len ;	// line#=../rle.cpp:24
reg	[7:0]	RG_len_03 ;	// line#=../rle.cpp:24
reg	[7:0]	RG_len_02 ;	// line#=../rle.cpp:24
reg	[6:0]	RG_140_02 ;
reg	[7:0]	RG_len_01 ;	// line#=../rle.cpp:24
reg	[6:0]	RG_142_01 ;
reg	[7:0]	RG_len_01_1 ;	// line#=../rle.cpp:24
reg	[6:0]	RG_k_01 ;	// line#=../rle.cpp:105
reg	[8:0]	jpeg_out_a00_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a01_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a02_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a03_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a04_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a05_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a06_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a07_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a08_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a09_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a10_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a11_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a12_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a13_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a14_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a15_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a16_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a17_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a18_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a19_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a20_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a21_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a22_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a23_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a24_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a25_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a26_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a27_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a28_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a29_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a30_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a31_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a32_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a33_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a34_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a35_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a36_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a37_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a38_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a39_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a40_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a41_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a42_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a43_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a44_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a45_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a46_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a47_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a48_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a49_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a50_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a51_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a52_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a53_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a54_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a55_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a56_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a57_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a58_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a59_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a60_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a61_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a62_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a63_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a64_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a65_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a66_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a67_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a68_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a69_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a70_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a71_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a72_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a73_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a74_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a75_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a76_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a77_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a78_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a79_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a80_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a81_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a82_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a83_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a84_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a85_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a86_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a87_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a88_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a89_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a90_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a91_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a92_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a93_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a94_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a95_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a96_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a97_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a98_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a99_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a100_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a101_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a102_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a103_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a104_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a105_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a106_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a107_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a108_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a109_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a110_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a111_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a112_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a113_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a114_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a115_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a116_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a117_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a118_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a119_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a120_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a121_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a122_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a123_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a124_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a125_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a126_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a127_r ;	// line#=../rle.h:60
reg	[11:0]	jpeg_len_out_r ;	// line#=../rle.h:61
reg	valid_r ;	// line#=../rle.h:62
reg	M_02_t1 ;
reg	M_03_t1 ;
reg	FL01_01_next ;
reg	[8:0]	RG_previous_dc_zz_t ;
reg	RG_previous_dc_zz_t_c1 ;
reg	RG_previous_dc_zz_t_c2 ;
reg	[8:0]	RG_zz_t ;
reg	RG_zz_t_c1 ;
reg	RG_zz_t_c2 ;
reg	[8:0]	RG_zz_1_t ;
reg	RG_zz_1_t_c1 ;
reg	RG_zz_1_t_c2 ;
reg	[8:0]	RG_zz_2_t ;
reg	RG_zz_2_t_c1 ;
reg	RG_zz_2_t_c2 ;
reg	[8:0]	RG_zz_3_t ;
reg	RG_zz_3_t_c1 ;
reg	RG_zz_3_t_c2 ;
reg	[8:0]	RG_zz_4_t ;
reg	RG_zz_4_t_c1 ;
reg	RG_zz_4_t_c2 ;
reg	[8:0]	RG_zz_5_t ;
reg	RG_zz_5_t_c1 ;
reg	RG_zz_5_t_c2 ;
reg	[8:0]	RG_zz_6_t ;
reg	RG_zz_6_t_c1 ;
reg	RG_zz_6_t_c2 ;
reg	[8:0]	RG_zz_7_t ;
reg	RG_zz_7_t_c1 ;
reg	RG_zz_7_t_c2 ;
reg	[8:0]	RG_zz_8_t ;
reg	RG_zz_8_t_c1 ;
reg	RG_zz_8_t_c2 ;
reg	[8:0]	RG_zz_9_t ;
reg	RG_zz_9_t_c1 ;
reg	RG_zz_9_t_c2 ;
reg	[8:0]	RG_zz_10_t ;
reg	RG_zz_10_t_c1 ;
reg	RG_zz_10_t_c2 ;
reg	[8:0]	RG_zz_11_t ;
reg	RG_zz_11_t_c1 ;
reg	RG_zz_11_t_c2 ;
reg	[8:0]	RG_zz_12_t ;
reg	RG_zz_12_t_c1 ;
reg	RG_zz_12_t_c2 ;
reg	[8:0]	RG_zz_13_t ;
reg	RG_zz_13_t_c1 ;
reg	RG_zz_13_t_c2 ;
reg	[8:0]	RG_zz_14_t ;
reg	RG_zz_14_t_c1 ;
reg	RG_zz_14_t_c2 ;
reg	[8:0]	RG_zz_15_t ;
reg	RG_zz_15_t_c1 ;
reg	RG_zz_15_t_c2 ;
reg	[8:0]	RG_zz_16_t ;
reg	RG_zz_16_t_c1 ;
reg	RG_zz_16_t_c2 ;
reg	[8:0]	RG_zz_17_t ;
reg	RG_zz_17_t_c1 ;
reg	RG_zz_17_t_c2 ;
reg	[8:0]	RG_zz_18_t ;
reg	RG_zz_18_t_c1 ;
reg	RG_zz_18_t_c2 ;
reg	[8:0]	RG_zz_19_t ;
reg	RG_zz_19_t_c1 ;
reg	RG_zz_19_t_c2 ;
reg	[8:0]	RG_zz_20_t ;
reg	RG_zz_20_t_c1 ;
reg	RG_zz_20_t_c2 ;
reg	[8:0]	RG_zz_21_t ;
reg	RG_zz_21_t_c1 ;
reg	RG_zz_21_t_c2 ;
reg	[8:0]	RG_zz_22_t ;
reg	RG_zz_22_t_c1 ;
reg	RG_zz_22_t_c2 ;
reg	[8:0]	RG_zz_23_t ;
reg	RG_zz_23_t_c1 ;
reg	RG_zz_23_t_c2 ;
reg	[8:0]	RG_zz_24_t ;
reg	RG_zz_24_t_c1 ;
reg	RG_zz_24_t_c2 ;
reg	[8:0]	RG_zz_25_t ;
reg	RG_zz_25_t_c1 ;
reg	RG_zz_25_t_c2 ;
reg	[8:0]	RG_zz_26_t ;
reg	RG_zz_26_t_c1 ;
reg	RG_zz_26_t_c2 ;
reg	[8:0]	RG_zz_27_t ;
reg	RG_zz_27_t_c1 ;
reg	RG_zz_27_t_c2 ;
reg	[8:0]	RG_zz_28_t ;
reg	RG_zz_28_t_c1 ;
reg	RG_zz_28_t_c2 ;
reg	[8:0]	RG_zz_29_t ;
reg	RG_zz_29_t_c1 ;
reg	RG_zz_29_t_c2 ;
reg	[8:0]	RG_zz_30_t ;
reg	RG_zz_30_t_c1 ;
reg	RG_zz_30_t_c2 ;
reg	[8:0]	RG_zz_31_t ;
reg	RG_zz_31_t_c1 ;
reg	RG_zz_31_t_c2 ;
reg	[8:0]	RG_zz_32_t ;
reg	RG_zz_32_t_c1 ;
reg	RG_zz_32_t_c2 ;
reg	[8:0]	RG_zz_33_t ;
reg	RG_zz_33_t_c1 ;
reg	RG_zz_33_t_c2 ;
reg	[8:0]	RG_zz_34_t ;
reg	RG_zz_34_t_c1 ;
reg	RG_zz_34_t_c2 ;
reg	[8:0]	RG_zz_35_t ;
reg	RG_zz_35_t_c1 ;
reg	RG_zz_35_t_c2 ;
reg	[8:0]	RG_zz_36_t ;
reg	RG_zz_36_t_c1 ;
reg	RG_zz_36_t_c2 ;
reg	[8:0]	RG_zz_37_t ;
reg	RG_zz_37_t_c1 ;
reg	RG_zz_37_t_c2 ;
reg	[8:0]	RG_zz_38_t ;
reg	RG_zz_38_t_c1 ;
reg	RG_zz_38_t_c2 ;
reg	[8:0]	RG_zz_39_t ;
reg	RG_zz_39_t_c1 ;
reg	RG_zz_39_t_c2 ;
reg	[8:0]	RG_zz_40_t ;
reg	RG_zz_40_t_c1 ;
reg	RG_zz_40_t_c2 ;
reg	[8:0]	RG_zz_41_t ;
reg	RG_zz_41_t_c1 ;
reg	RG_zz_41_t_c2 ;
reg	[8:0]	RG_zz_42_t ;
reg	RG_zz_42_t_c1 ;
reg	RG_zz_42_t_c2 ;
reg	[8:0]	RG_zz_43_t ;
reg	RG_zz_43_t_c1 ;
reg	RG_zz_43_t_c2 ;
reg	[8:0]	RG_zz_44_t ;
reg	RG_zz_44_t_c1 ;
reg	RG_zz_44_t_c2 ;
reg	[8:0]	RG_zz_45_t ;
reg	RG_zz_45_t_c1 ;
reg	RG_zz_45_t_c2 ;
reg	[8:0]	RG_zz_46_t ;
reg	RG_zz_46_t_c1 ;
reg	RG_zz_46_t_c2 ;
reg	[8:0]	RG_zz_47_t ;
reg	RG_zz_47_t_c1 ;
reg	RG_zz_47_t_c2 ;
reg	[8:0]	RG_zz_48_t ;
reg	RG_zz_48_t_c1 ;
reg	RG_zz_48_t_c2 ;
reg	[8:0]	RG_zz_49_t ;
reg	RG_zz_49_t_c1 ;
reg	RG_zz_49_t_c2 ;
reg	[8:0]	RG_zz_50_t ;
reg	RG_zz_50_t_c1 ;
reg	RG_zz_50_t_c2 ;
reg	[8:0]	RG_zz_51_t ;
reg	RG_zz_51_t_c1 ;
reg	RG_zz_51_t_c2 ;
reg	[8:0]	RG_zz_52_t ;
reg	RG_zz_52_t_c1 ;
reg	RG_zz_52_t_c2 ;
reg	[8:0]	RG_zz_53_t ;
reg	RG_zz_53_t_c1 ;
reg	RG_zz_53_t_c2 ;
reg	[8:0]	RG_zz_54_t ;
reg	RG_zz_54_t_c1 ;
reg	RG_zz_54_t_c2 ;
reg	[8:0]	RG_zz_55_t ;
reg	RG_zz_55_t_c1 ;
reg	RG_zz_55_t_c2 ;
reg	[8:0]	RG_zz_56_t ;
reg	RG_zz_56_t_c1 ;
reg	RG_zz_56_t_c2 ;
reg	[8:0]	RG_zz_57_t ;
reg	RG_zz_57_t_c1 ;
reg	RG_zz_57_t_c2 ;
reg	[8:0]	RG_zz_58_t ;
reg	RG_zz_58_t_c1 ;
reg	RG_zz_58_t_c2 ;
reg	[8:0]	RG_zz_59_t ;
reg	RG_zz_59_t_c1 ;
reg	RG_zz_59_t_c2 ;
reg	[8:0]	RG_zz_60_t ;
reg	RG_zz_60_t_c1 ;
reg	RG_zz_60_t_c2 ;
reg	[8:0]	RG_zz_61_t ;
reg	RG_zz_61_t_c1 ;
reg	RG_zz_61_t_c2 ;
reg	[8:0]	RG_zz_62_t ;
reg	RG_zz_62_t_c1 ;
reg	RG_zz_62_t_c2 ;
reg	[3:0]	RG_j_03_t ;
reg	[2:0]	TR_01 ;
reg	[31:0]	RG_i_t ;
reg	RG_i_t_c1 ;
reg	RG_i_t_c2 ;
reg	RG_i_t_c3 ;
reg	[31:0]	RG_j_k_t ;
reg	RG_j_k_t_c1 ;
reg	RG_j_k_t_c2 ;
reg	RG_j_k_t_c3 ;
reg	[8:0]	RG_quantized_block_rl_02_t ;
reg	[8:0]	RG_quantized_block_rl_02_1_t ;
reg	[8:0]	RG_quantized_block_zz_t ;
reg	[5:0]	RG_k_t ;
reg	FF_d_t ;
reg	FF_d_t_c1 ;
reg	FF_d_t_c2 ;
reg	FF_i_t ;
reg	FF_len_t ;
reg	[6:0]	RG_142_01_t ;
reg	[7:0]	RG_len_01_1_t ;
reg	RG_len_01_1_t_c1 ;
reg	[6:0]	RG_k_01_t ;
reg	RG_k_01_t_c1 ;
reg	[8:0]	TR_44 ;
reg	[8:0]	TR_45 ;
reg	[8:0]	TR_46 ;
reg	[8:0]	TR_47 ;
reg	[8:0]	TR_48 ;
reg	[8:0]	TR_49 ;
reg	[8:0]	TR_50 ;
reg	[8:0]	TR_51 ;
reg	[8:0]	M_217 ;
reg	M_217_c1 ;
reg	M_217_c2 ;
reg	M_217_c3 ;
reg	M_217_c4 ;
reg	M_217_c5 ;
reg	M_217_c6 ;
reg	M_217_c7 ;
reg	M_217_c8 ;
reg	M_01_t64 ;
reg	M_01_t64_t1 ;
reg	FL01_01_streg_t ;
reg	FL01_01_streg_t_c1 ;
reg	FL01_02_streg_t ;
reg	FL01_02_streg_t_c1 ;
reg	FL01_02_streg_t_c2 ;
reg	FL01_03_streg_t ;
reg	FL01_03_streg_t_c1 ;
reg	FL01_03_streg_t_c2 ;
reg	valid_r_t ;
reg	[5:0]	TR_03 ;
reg	[7:0]	incr8u2i1 ;
reg	incr8u2i1_c1 ;
reg	[6:0]	sub8u_7_11i1 ;
reg	sub8u_7_11i1_c1 ;
reg	[1:0]	M_220 ;
reg	[1:0]	TR_17 ;
reg	[2:0]	TR_18 ;
reg	[3:0]	TR_05 ;
reg	TR_05_c1 ;
reg	[2:0]	TR_19 ;
reg	[2:0]	TR_32 ;
reg	[3:0]	TR_20 ;
reg	TR_20_c1 ;
reg	[4:0]	TR_06 ;
reg	TR_06_c1 ;
reg	[1:0]	TR_21 ;
reg	[2:0]	TR_22 ;
reg	[2:0]	TR_33 ;
reg	[3:0]	TR_23 ;
reg	TR_23_c1 ;
reg	[2:0]	TR_34 ;
reg	[1:0]	TR_41 ;
reg	[2:0]	TR_42 ;
reg	[3:0]	TR_35 ;
reg	TR_35_c1 ;
reg	[4:0]	TR_24 ;
reg	TR_24_c1 ;
reg	[5:0]	TR_07 ;
reg	TR_07_c1 ;
reg	[2:0]	TR_08 ;
reg	[2:0]	TR_25 ;
reg	[3:0]	TR_09 ;
reg	TR_09_c1 ;
reg	[1:0]	TR_26 ;
reg	[2:0]	TR_27 ;
reg	[2:0]	TR_36 ;
reg	[3:0]	TR_28 ;
reg	TR_28_c1 ;
reg	[4:0]	TR_10 ;
reg	TR_10_c1 ;
reg	[2:0]	TR_29 ;
reg	[1:0]	TR_37 ;
reg	[2:0]	TR_38 ;
reg	[3:0]	TR_30 ;
reg	TR_30_c1 ;
reg	[2:0]	TR_39 ;
reg	[2:0]	TR_43 ;
reg	[3:0]	TR_40 ;
reg	TR_40_c1 ;
reg	[4:0]	TR_31 ;
reg	TR_31_c1 ;
reg	[5:0]	TR_11 ;
reg	TR_11_c1 ;
reg	[6:0]	rl_AD1 ;
reg	rl_AD1_c1 ;
reg	rl_AD1_c2 ;
reg	rl_AD1_c3 ;
reg	[8:0]	rl_WD1 ;
reg	[8:0]	rl_WD1_t1 ;
reg	[5:0]	TR_12 ;
reg	[5:0]	TR_13 ;
reg	[6:0]	rl_RA2 ;
reg	rl_RA2_c1 ;
reg	[5:0]	TR_14 ;
reg	[5:0]	TR_15 ;
reg	[6:0]	rl_RA3 ;

jpeg_sub8u_7_1 INST_sub8u_7_1_1 ( .i1(sub8u_7_11i1) ,.i2(sub8u_7_11i2) ,.o1(sub8u_7_11ot) );	// line#=../rle.cpp:77,78,83,84
jpeg_sub8u_7 INST_sub8u_7_1 ( .i1(sub8u_71i1) ,.i2(sub8u_71i2) ,.o1(sub8u_71ot) );	// line#=../rle.cpp:83,84
jpeg_decr32s INST_decr32s_1 ( .i1(decr32s1i1) ,.o1(decr32s1ot) );	// line#=../rle.cpp:124,155
jpeg_decr32s INST_decr32s_2 ( .i1(decr32s2i1) ,.o1(decr32s2ot) );	// line#=../rle.cpp:130,161
jpeg_decr8u_7 INST_decr8u_7_1 ( .i1(decr8u_71i1) ,.o1(decr8u_71ot) );	// line#=../rle.cpp:77,78
jpeg_incr32s INST_incr32s_1 ( .i1(incr32s1i1) ,.o1(incr32s1ot) );	// line#=../rle.cpp:64,114,125,145,156
jpeg_incr32s INST_incr32s_2 ( .i1(incr32s2i1) ,.o1(incr32s2ot) );	// line#=../rle.cpp:63,74,119,129,150,160
jpeg_incr8u INST_incr8u_1 ( .i1(incr8u1i1) ,.o1(incr8u1ot) );	// line#=../rle.cpp:68,73,79
jpeg_incr8u INST_incr8u_2 ( .i1(incr8u2i1) ,.o1(incr8u2ot) );	// line#=../rle.cpp:69,74,80,111,142
jpeg_incr4s INST_incr4s_1 ( .i1(incr4s1i1) ,.o1(incr4s1ot) );	// line#=../rle.cpp:34
jpeg_lop8u_1 INST_lop8u_1_1 ( .i1(lop8u_11i1) ,.i2(lop8u_11i2) ,.o1(lop8u_11ot) );	// line#=../rle.cpp:109,110
assign	lop8u_11ot_port = lop8u_11ot ;
jpeg_sub12s_9 INST_sub12s_9_1 ( .i1(sub12s_91i1) ,.i2(sub12s_91i2) ,.o1(sub12s_91ot) );	// line#=../rle.cpp:52
jpeg_sub8u INST_sub8u_1 ( .i1(sub8u1i1) ,.i2(sub8u1i2) ,.o1(sub8u1ot) );	// line#=../rle.cpp:83,84,86
assign	jpeg_out_a00 = jpeg_out_a00_r ;	// line#=../rle.h:60
assign	jpeg_out_a01 = jpeg_out_a01_r ;	// line#=../rle.h:60
assign	jpeg_out_a02 = jpeg_out_a02_r ;	// line#=../rle.h:60
assign	jpeg_out_a03 = jpeg_out_a03_r ;	// line#=../rle.h:60
assign	jpeg_out_a04 = jpeg_out_a04_r ;	// line#=../rle.h:60
assign	jpeg_out_a05 = jpeg_out_a05_r ;	// line#=../rle.h:60
assign	jpeg_out_a06 = jpeg_out_a06_r ;	// line#=../rle.h:60
assign	jpeg_out_a07 = jpeg_out_a07_r ;	// line#=../rle.h:60
assign	jpeg_out_a08 = jpeg_out_a08_r ;	// line#=../rle.h:60
assign	jpeg_out_a09 = jpeg_out_a09_r ;	// line#=../rle.h:60
assign	jpeg_out_a10 = jpeg_out_a10_r ;	// line#=../rle.h:60
assign	jpeg_out_a11 = jpeg_out_a11_r ;	// line#=../rle.h:60
assign	jpeg_out_a12 = jpeg_out_a12_r ;	// line#=../rle.h:60
assign	jpeg_out_a13 = jpeg_out_a13_r ;	// line#=../rle.h:60
assign	jpeg_out_a14 = jpeg_out_a14_r ;	// line#=../rle.h:60
assign	jpeg_out_a15 = jpeg_out_a15_r ;	// line#=../rle.h:60
assign	jpeg_out_a16 = jpeg_out_a16_r ;	// line#=../rle.h:60
assign	jpeg_out_a17 = jpeg_out_a17_r ;	// line#=../rle.h:60
assign	jpeg_out_a18 = jpeg_out_a18_r ;	// line#=../rle.h:60
assign	jpeg_out_a19 = jpeg_out_a19_r ;	// line#=../rle.h:60
assign	jpeg_out_a20 = jpeg_out_a20_r ;	// line#=../rle.h:60
assign	jpeg_out_a21 = jpeg_out_a21_r ;	// line#=../rle.h:60
assign	jpeg_out_a22 = jpeg_out_a22_r ;	// line#=../rle.h:60
assign	jpeg_out_a23 = jpeg_out_a23_r ;	// line#=../rle.h:60
assign	jpeg_out_a24 = jpeg_out_a24_r ;	// line#=../rle.h:60
assign	jpeg_out_a25 = jpeg_out_a25_r ;	// line#=../rle.h:60
assign	jpeg_out_a26 = jpeg_out_a26_r ;	// line#=../rle.h:60
assign	jpeg_out_a27 = jpeg_out_a27_r ;	// line#=../rle.h:60
assign	jpeg_out_a28 = jpeg_out_a28_r ;	// line#=../rle.h:60
assign	jpeg_out_a29 = jpeg_out_a29_r ;	// line#=../rle.h:60
assign	jpeg_out_a30 = jpeg_out_a30_r ;	// line#=../rle.h:60
assign	jpeg_out_a31 = jpeg_out_a31_r ;	// line#=../rle.h:60
assign	jpeg_out_a32 = jpeg_out_a32_r ;	// line#=../rle.h:60
assign	jpeg_out_a33 = jpeg_out_a33_r ;	// line#=../rle.h:60
assign	jpeg_out_a34 = jpeg_out_a34_r ;	// line#=../rle.h:60
assign	jpeg_out_a35 = jpeg_out_a35_r ;	// line#=../rle.h:60
assign	jpeg_out_a36 = jpeg_out_a36_r ;	// line#=../rle.h:60
assign	jpeg_out_a37 = jpeg_out_a37_r ;	// line#=../rle.h:60
assign	jpeg_out_a38 = jpeg_out_a38_r ;	// line#=../rle.h:60
assign	jpeg_out_a39 = jpeg_out_a39_r ;	// line#=../rle.h:60
assign	jpeg_out_a40 = jpeg_out_a40_r ;	// line#=../rle.h:60
assign	jpeg_out_a41 = jpeg_out_a41_r ;	// line#=../rle.h:60
assign	jpeg_out_a42 = jpeg_out_a42_r ;	// line#=../rle.h:60
assign	jpeg_out_a43 = jpeg_out_a43_r ;	// line#=../rle.h:60
assign	jpeg_out_a44 = jpeg_out_a44_r ;	// line#=../rle.h:60
assign	jpeg_out_a45 = jpeg_out_a45_r ;	// line#=../rle.h:60
assign	jpeg_out_a46 = jpeg_out_a46_r ;	// line#=../rle.h:60
assign	jpeg_out_a47 = jpeg_out_a47_r ;	// line#=../rle.h:60
assign	jpeg_out_a48 = jpeg_out_a48_r ;	// line#=../rle.h:60
assign	jpeg_out_a49 = jpeg_out_a49_r ;	// line#=../rle.h:60
assign	jpeg_out_a50 = jpeg_out_a50_r ;	// line#=../rle.h:60
assign	jpeg_out_a51 = jpeg_out_a51_r ;	// line#=../rle.h:60
assign	jpeg_out_a52 = jpeg_out_a52_r ;	// line#=../rle.h:60
assign	jpeg_out_a53 = jpeg_out_a53_r ;	// line#=../rle.h:60
assign	jpeg_out_a54 = jpeg_out_a54_r ;	// line#=../rle.h:60
assign	jpeg_out_a55 = jpeg_out_a55_r ;	// line#=../rle.h:60
assign	jpeg_out_a56 = jpeg_out_a56_r ;	// line#=../rle.h:60
assign	jpeg_out_a57 = jpeg_out_a57_r ;	// line#=../rle.h:60
assign	jpeg_out_a58 = jpeg_out_a58_r ;	// line#=../rle.h:60
assign	jpeg_out_a59 = jpeg_out_a59_r ;	// line#=../rle.h:60
assign	jpeg_out_a60 = jpeg_out_a60_r ;	// line#=../rle.h:60
assign	jpeg_out_a61 = jpeg_out_a61_r ;	// line#=../rle.h:60
assign	jpeg_out_a62 = jpeg_out_a62_r ;	// line#=../rle.h:60
assign	jpeg_out_a63 = jpeg_out_a63_r ;	// line#=../rle.h:60
assign	jpeg_out_a64 = jpeg_out_a64_r ;	// line#=../rle.h:60
assign	jpeg_out_a65 = jpeg_out_a65_r ;	// line#=../rle.h:60
assign	jpeg_out_a66 = jpeg_out_a66_r ;	// line#=../rle.h:60
assign	jpeg_out_a67 = jpeg_out_a67_r ;	// line#=../rle.h:60
assign	jpeg_out_a68 = jpeg_out_a68_r ;	// line#=../rle.h:60
assign	jpeg_out_a69 = jpeg_out_a69_r ;	// line#=../rle.h:60
assign	jpeg_out_a70 = jpeg_out_a70_r ;	// line#=../rle.h:60
assign	jpeg_out_a71 = jpeg_out_a71_r ;	// line#=../rle.h:60
assign	jpeg_out_a72 = jpeg_out_a72_r ;	// line#=../rle.h:60
assign	jpeg_out_a73 = jpeg_out_a73_r ;	// line#=../rle.h:60
assign	jpeg_out_a74 = jpeg_out_a74_r ;	// line#=../rle.h:60
assign	jpeg_out_a75 = jpeg_out_a75_r ;	// line#=../rle.h:60
assign	jpeg_out_a76 = jpeg_out_a76_r ;	// line#=../rle.h:60
assign	jpeg_out_a77 = jpeg_out_a77_r ;	// line#=../rle.h:60
assign	jpeg_out_a78 = jpeg_out_a78_r ;	// line#=../rle.h:60
assign	jpeg_out_a79 = jpeg_out_a79_r ;	// line#=../rle.h:60
assign	jpeg_out_a80 = jpeg_out_a80_r ;	// line#=../rle.h:60
assign	jpeg_out_a81 = jpeg_out_a81_r ;	// line#=../rle.h:60
assign	jpeg_out_a82 = jpeg_out_a82_r ;	// line#=../rle.h:60
assign	jpeg_out_a83 = jpeg_out_a83_r ;	// line#=../rle.h:60
assign	jpeg_out_a84 = jpeg_out_a84_r ;	// line#=../rle.h:60
assign	jpeg_out_a85 = jpeg_out_a85_r ;	// line#=../rle.h:60
assign	jpeg_out_a86 = jpeg_out_a86_r ;	// line#=../rle.h:60
assign	jpeg_out_a87 = jpeg_out_a87_r ;	// line#=../rle.h:60
assign	jpeg_out_a88 = jpeg_out_a88_r ;	// line#=../rle.h:60
assign	jpeg_out_a89 = jpeg_out_a89_r ;	// line#=../rle.h:60
assign	jpeg_out_a90 = jpeg_out_a90_r ;	// line#=../rle.h:60
assign	jpeg_out_a91 = jpeg_out_a91_r ;	// line#=../rle.h:60
assign	jpeg_out_a92 = jpeg_out_a92_r ;	// line#=../rle.h:60
assign	jpeg_out_a93 = jpeg_out_a93_r ;	// line#=../rle.h:60
assign	jpeg_out_a94 = jpeg_out_a94_r ;	// line#=../rle.h:60
assign	jpeg_out_a95 = jpeg_out_a95_r ;	// line#=../rle.h:60
assign	jpeg_out_a96 = jpeg_out_a96_r ;	// line#=../rle.h:60
assign	jpeg_out_a97 = jpeg_out_a97_r ;	// line#=../rle.h:60
assign	jpeg_out_a98 = jpeg_out_a98_r ;	// line#=../rle.h:60
assign	jpeg_out_a99 = jpeg_out_a99_r ;	// line#=../rle.h:60
assign	jpeg_out_a100 = jpeg_out_a100_r ;	// line#=../rle.h:60
assign	jpeg_out_a101 = jpeg_out_a101_r ;	// line#=../rle.h:60
assign	jpeg_out_a102 = jpeg_out_a102_r ;	// line#=../rle.h:60
assign	jpeg_out_a103 = jpeg_out_a103_r ;	// line#=../rle.h:60
assign	jpeg_out_a104 = jpeg_out_a104_r ;	// line#=../rle.h:60
assign	jpeg_out_a105 = jpeg_out_a105_r ;	// line#=../rle.h:60
assign	jpeg_out_a106 = jpeg_out_a106_r ;	// line#=../rle.h:60
assign	jpeg_out_a107 = jpeg_out_a107_r ;	// line#=../rle.h:60
assign	jpeg_out_a108 = jpeg_out_a108_r ;	// line#=../rle.h:60
assign	jpeg_out_a109 = jpeg_out_a109_r ;	// line#=../rle.h:60
assign	jpeg_out_a110 = jpeg_out_a110_r ;	// line#=../rle.h:60
assign	jpeg_out_a111 = jpeg_out_a111_r ;	// line#=../rle.h:60
assign	jpeg_out_a112 = jpeg_out_a112_r ;	// line#=../rle.h:60
assign	jpeg_out_a113 = jpeg_out_a113_r ;	// line#=../rle.h:60
assign	jpeg_out_a114 = jpeg_out_a114_r ;	// line#=../rle.h:60
assign	jpeg_out_a115 = jpeg_out_a115_r ;	// line#=../rle.h:60
assign	jpeg_out_a116 = jpeg_out_a116_r ;	// line#=../rle.h:60
assign	jpeg_out_a117 = jpeg_out_a117_r ;	// line#=../rle.h:60
assign	jpeg_out_a118 = jpeg_out_a118_r ;	// line#=../rle.h:60
assign	jpeg_out_a119 = jpeg_out_a119_r ;	// line#=../rle.h:60
assign	jpeg_out_a120 = jpeg_out_a120_r ;	// line#=../rle.h:60
assign	jpeg_out_a121 = jpeg_out_a121_r ;	// line#=../rle.h:60
assign	jpeg_out_a122 = jpeg_out_a122_r ;	// line#=../rle.h:60
assign	jpeg_out_a123 = jpeg_out_a123_r ;	// line#=../rle.h:60
assign	jpeg_out_a124 = jpeg_out_a124_r ;	// line#=../rle.h:60
assign	jpeg_out_a125 = jpeg_out_a125_r ;	// line#=../rle.h:60
assign	jpeg_out_a126 = jpeg_out_a126_r ;	// line#=../rle.h:60
assign	jpeg_out_a127 = jpeg_out_a127_r ;	// line#=../rle.h:60
assign	jpeg_len_out = jpeg_len_out_r ;	// line#=../rle.h:61
assign	valid = valid_r ;	// line#=../rle.h:62
always @ ( posedge clk )	// line#=../rle.cpp:61,62
	RG_136 <= CT_30 ;
always @ ( posedge clk )
	RG_len_02 <= RG_len_01 ;
always @ ( posedge clk )	// line#=../rle.cpp:83,84
	RG_140_02 <= RG_142_01 ;
always @ ( posedge clk )
	RG_len_01 <= RG_len_01_1 ;
assign	CT_03 = ( ( ~|RG_j_k ) & M_106 ) ;	// line#=../rle.cpp:117,118
assign	M_106 = ~|{ ( RG_i [31] & RG_i [0] ) , ~RG_i [0] } ;	// line#=../rle.cpp:117,118,148,149
assign	CT_18 = ( ( ~|{ RG_j_k [31:3] , ~RG_j_k [2:0] } ) & M_106 ) ;	// line#=../rle.cpp:148,149
assign	CT_30 = ( M_01_t64 & ( RG_j_k [31] | ( ( ~|RG_j_k [30:4] ) & ( ~&RG_j_k [3:0] ) ) ) ) ;	// line#=../rle.cpp:61,62
assign	CT_30_port = CT_30 ;
assign	CT_33 = ~|{ RG_i [31:7] , ~RG_i [6] , RG_i [5:0] } ;	// line#=../rle.cpp:66,67
assign	CT_35 = ( RG_i [31] | ( ~|RG_i [30:6] ) ) ;	// line#=../rle.cpp:57,58,61,62
assign	CT_35_port = CT_35 ;
always @ ( M_184 or RG_quantized_block_rl_02 )	// line#=../rle.cpp:77,78
	case ( ~|RG_quantized_block_rl_02 )
	1'h1 :
		M_02_t1 = M_184 ;	// line#=../rle.cpp:77,78
	1'h0 :
		M_02_t1 = 1'h0 ;	// line#=../rle.cpp:77,78
	default :
		M_02_t1 = 1'hx ;
	endcase
assign	M_184 = ~|RG_quantized_block_rl_02_1 ;	// line#=../rle.cpp:77,78,83,84
always @ ( M_184 or RG_quantized_block_rl_02 )	// line#=../rle.cpp:83,84
	case ( ~|{ RG_quantized_block_rl_02 [8:4] , ~RG_quantized_block_rl_02 [3:0] } )
	1'h1 :
		M_03_t1 = M_184 ;	// line#=../rle.cpp:83,84
	1'h0 :
		M_03_t1 = 1'h0 ;	// line#=../rle.cpp:83,84
	default :
		M_03_t1 = 1'hx ;
	endcase
assign	FL01_01_Leos_all = ( ( FL01_01_eos & FL01_02_eos ) & FL01_03_eos ) ;
always @ ( FL01_01_streg )
	case ( FL01_01_streg )
	1'h0 :
		FL01_01_next = 1'h0 ;
	1'h1 :
		FL01_01_next = 1'h1 ;
	default :
		FL01_01_next = 1'hx ;
	endcase
assign	sub8u1i1 = RG_len_01_1 ;	// line#=../rle.cpp:83,84,86
assign	sub8u1i2 = 2'h2 ;	// line#=../rle.cpp:83,84,86
assign	sub12s_91i1 = RG_previous_dc_zz ;	// line#=../rle.cpp:52
assign	sub12s_91i2 = RG_previous_dc ;	// line#=../rle.cpp:52
assign	lop8u_11i1 = RG_k ;	// line#=../rle.cpp:109,110
assign	lop8u_11i2 = 6'h24 ;	// line#=../rle.cpp:109,110
assign	incr4s1i1 = RG_j_03 ;	// line#=../rle.cpp:34
assign	decr8u_71i1 = incr8u2ot [6:0] ;	// line#=../rle.cpp:69,74,77,78
assign	sub8u_71i1 = RG_len_01_1 [6:0] ;	// line#=../rle.cpp:83,84
assign	sub8u_71i2 = 3'h4 ;	// line#=../rle.cpp:83,84
assign	U_05 = ( ST1_03d & lop8u_11ot ) ;	// line#=../rle.cpp:109,110
assign	U_06 = ( ST1_03d & ( ~lop8u_11ot ) ) ;	// line#=../rle.cpp:109,110
assign	C_02 = ( ( ~|RG_i ) & M_183 ) ;	// line#=../rle.cpp:112,113
assign	U_79 = ( U_05 & C_02 ) ;	// line#=../rle.cpp:112,113
assign	U_80 = ( U_05 & ( ~C_02 ) ) ;	// line#=../rle.cpp:112,113
assign	U_81 = ( U_80 & CT_03 ) ;	// line#=../rle.cpp:117,118
assign	U_82 = ( U_80 & ( ~CT_03 ) ) ;	// line#=../rle.cpp:117,118
assign	U_83 = ( U_82 & ( ~FF_d ) ) ;	// line#=../rle.cpp:122,123
assign	U_84 = ( U_82 & FF_d ) ;	// line#=../rle.cpp:122,123
assign	U_87 = ( ST1_04d & ( ~RG_k_01 [6] ) ) ;	// line#=../rle.cpp:140,141
assign	U_88 = ( ST1_04d & RG_k_01 [6] ) ;	// line#=../rle.cpp:140,141
assign	M_183 = ~|{ ( RG_j_k [31] & RG_j_k [0] ) , RG_j_k [0] } ;	// line#=../rle.cpp:112,113,143,144
assign	C_05 = ( ( ~|{ RG_i [31:3] , ~RG_i [2:0] } ) & M_183 ) ;	// line#=../rle.cpp:143,144
assign	U_161 = ( U_87 & C_05 ) ;	// line#=../rle.cpp:143,144
assign	U_162 = ( U_87 & ( ~C_05 ) ) ;	// line#=../rle.cpp:143,144
assign	U_163 = ( U_162 & CT_18 ) ;	// line#=../rle.cpp:148,149
assign	U_164 = ( U_162 & ( ~CT_18 ) ) ;	// line#=../rle.cpp:148,149
assign	U_165 = ( U_164 & ( ~FF_d ) ) ;	// line#=../rle.cpp:153,154
assign	U_166 = ( U_164 & FF_d ) ;	// line#=../rle.cpp:153,154
assign	U_169 = ( ST1_05d & CT_30 ) ;	// line#=../rle.cpp:61,62
assign	U_175 = ( ST1_06d & ( ~RG_136 ) ) ;	// line#=../rle.cpp:61,62
assign	U_176 = ( U_175 & CT_33 ) ;	// line#=../rle.cpp:66,67
assign	U_177 = ( U_175 & ( ~CT_33 ) ) ;	// line#=../rle.cpp:66,67
assign	U_178 = ( ST1_07d & FF_i ) ;	// line#=../rle.cpp:66,67
assign	U_179 = ( ST1_07d & ( ~FF_i ) ) ;	// line#=../rle.cpp:66,67
assign	U_248 = ( ST1_09d & ( ~M_02_t1 ) ) ;	// line#=../rle.cpp:77,78
assign	U_251 = ( ST1_09d & ( ~JF_06 ) ) ;
assign	U_252 = ( ST1_11d & FL01_01_01a ) ;
assign	U_254 = ( ST1_11d & FL01_03_01a ) ;
assign	U_257 = ( U_254 & M_03_t1 ) ;	// line#=../rle.cpp:83,84
assign	U_262 = ( ST1_11d & ( ~FL01_02_streg ) ) ;
assign	U_263 = ( ST1_11d & FL01_02_streg ) ;
assign	U_268 = ( ST1_11d & ( ~FL01_03_streg ) ) ;
assign	U_269 = ( ST1_11d & FL01_03_streg ) ;
assign	U_273 = ( U_269 & ( ~FJ_13_14 ) ) ;
assign	U_278 = ( ST1_11d & FJ_13_14 ) ;
assign	U_280 = ( ST1_11d & FL01_03_break ) ;
assign	RG_previous_dc_en = ST1_54d ;
always @ ( posedge clk )
	if ( !rst )
		RG_previous_dc <= 9'h000 ;
	else if ( RG_previous_dc_en )
		RG_previous_dc <= RG_previous_dc_zz ;
always @ ( RG_quantized_block_zz or ST1_54d or RG_k_01 or U_87 or M_217 or M_110 or 
	U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_previous_dc_zz_t_c1 = ( U_05 & M_110 ) ;	// line#=../rle.cpp:111
	RG_previous_dc_zz_t_c2 = ( U_87 & ( ~|RG_k_01 [5:0] ) ) ;	// line#=../rle.cpp:142
	RG_previous_dc_zz_t = ( ( { 9{ RG_previous_dc_zz_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_previous_dc_zz_t_c2 } } & M_217 )			// line#=../rle.cpp:142
		| ( { 9{ ST1_54d } } & RG_quantized_block_zz ) ) ;
	end
assign	RG_previous_dc_zz_en = ( RG_previous_dc_zz_t_c1 | RG_previous_dc_zz_t_c2 | 
	ST1_54d ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_previous_dc_zz_en )
		RG_previous_dc_zz <= RG_previous_dc_zz_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_107 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_t_c1 = ( U_05 & M_107 ) ;	// line#=../rle.cpp:111
	RG_zz_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h01 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_t = ( ( { 9{ RG_zz_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_en = ( RG_zz_t_c1 | RG_zz_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_en )
		RG_zz <= RG_zz_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_116 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_1_t_c1 = ( U_05 & M_116 ) ;	// line#=../rle.cpp:111
	RG_zz_1_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h02 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_1_t = ( ( { 9{ RG_zz_1_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_1_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_1_en = ( RG_zz_1_t_c1 | RG_zz_1_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_1_en )
		RG_zz_1 <= RG_zz_1_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_124 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_2_t_c1 = ( U_05 & M_124 ) ;	// line#=../rle.cpp:111
	RG_zz_2_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h03 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_2_t = ( ( { 9{ RG_zz_2_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_2_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_2_en = ( RG_zz_2_t_c1 | RG_zz_2_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_2_en )
		RG_zz_2 <= RG_zz_2_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_122 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_3_t_c1 = ( U_05 & M_122 ) ;	// line#=../rle.cpp:111
	RG_zz_3_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h04 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_3_t = ( ( { 9{ RG_zz_3_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_3_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_3_en = ( RG_zz_3_t_c1 | RG_zz_3_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_3_en )
		RG_zz_3 <= RG_zz_3_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_126 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_4_t_c1 = ( U_05 & M_126 ) ;	// line#=../rle.cpp:111
	RG_zz_4_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h05 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_4_t = ( ( { 9{ RG_zz_4_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_4_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_4_en = ( RG_zz_4_t_c1 | RG_zz_4_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_4_en )
		RG_zz_4 <= RG_zz_4_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_128 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_5_t_c1 = ( U_05 & M_128 ) ;	// line#=../rle.cpp:111
	RG_zz_5_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h06 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_5_t = ( ( { 9{ RG_zz_5_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_5_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_5_en = ( RG_zz_5_t_c1 | RG_zz_5_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_5_en )
		RG_zz_5 <= RG_zz_5_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_118 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_6_t_c1 = ( U_05 & M_118 ) ;	// line#=../rle.cpp:111
	RG_zz_6_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h07 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_6_t = ( ( { 9{ RG_zz_6_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_6_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_6_en = ( RG_zz_6_t_c1 | RG_zz_6_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_6_en )
		RG_zz_6 <= RG_zz_6_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_114 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_7_t_c1 = ( U_05 & M_114 ) ;	// line#=../rle.cpp:111
	RG_zz_7_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h08 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_7_t = ( ( { 9{ RG_zz_7_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_7_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_7_en = ( RG_zz_7_t_c1 | RG_zz_7_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_7_en )
		RG_zz_7 <= RG_zz_7_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_182 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_8_t_c1 = ( U_05 & M_182 ) ;	// line#=../rle.cpp:111
	RG_zz_8_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h09 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_8_t = ( ( { 9{ RG_zz_8_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_8_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_8_en = ( RG_zz_8_t_c1 | RG_zz_8_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_8_en )
		RG_zz_8 <= RG_zz_8_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_181 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_9_t_c1 = ( U_05 & M_181 ) ;	// line#=../rle.cpp:111
	RG_zz_9_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h0a ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_9_t = ( ( { 9{ RG_zz_9_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_9_t_c2 } } & M_217 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_9_en = ( RG_zz_9_t_c1 | RG_zz_9_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_9_en )
		RG_zz_9 <= RG_zz_9_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_180 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_10_t_c1 = ( U_05 & M_180 ) ;	// line#=../rle.cpp:111
	RG_zz_10_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h0b ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_10_t = ( ( { 9{ RG_zz_10_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_10_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_10_en = ( RG_zz_10_t_c1 | RG_zz_10_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_10_en )
		RG_zz_10 <= RG_zz_10_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_179 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_11_t_c1 = ( U_05 & M_179 ) ;	// line#=../rle.cpp:111
	RG_zz_11_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h0c ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_11_t = ( ( { 9{ RG_zz_11_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_11_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_11_en = ( RG_zz_11_t_c1 | RG_zz_11_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_11_en )
		RG_zz_11 <= RG_zz_11_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_178 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_12_t_c1 = ( U_05 & M_178 ) ;	// line#=../rle.cpp:111
	RG_zz_12_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h0d ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_12_t = ( ( { 9{ RG_zz_12_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_12_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_12_en = ( RG_zz_12_t_c1 | RG_zz_12_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_12_en )
		RG_zz_12 <= RG_zz_12_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_177 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_13_t_c1 = ( U_05 & M_177 ) ;	// line#=../rle.cpp:111
	RG_zz_13_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h0e ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_13_t = ( ( { 9{ RG_zz_13_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_13_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_13_en = ( RG_zz_13_t_c1 | RG_zz_13_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_13_en )
		RG_zz_13 <= RG_zz_13_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_120 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_14_t_c1 = ( U_05 & M_120 ) ;	// line#=../rle.cpp:111
	RG_zz_14_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h0f ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_14_t = ( ( { 9{ RG_zz_14_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_14_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_14_en = ( RG_zz_14_t_c1 | RG_zz_14_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_14_en )
		RG_zz_14 <= RG_zz_14_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_176 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_15_t_c1 = ( U_05 & M_176 ) ;	// line#=../rle.cpp:111
	RG_zz_15_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h10 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_15_t = ( ( { 9{ RG_zz_15_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_15_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_15_en = ( RG_zz_15_t_c1 | RG_zz_15_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_15_en )
		RG_zz_15 <= RG_zz_15_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_175 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_16_t_c1 = ( U_05 & M_175 ) ;	// line#=../rle.cpp:111
	RG_zz_16_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h11 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_16_t = ( ( { 9{ RG_zz_16_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_16_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_16_en = ( RG_zz_16_t_c1 | RG_zz_16_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_16_en )
		RG_zz_16 <= RG_zz_16_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_174 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_17_t_c1 = ( U_05 & M_174 ) ;	// line#=../rle.cpp:111
	RG_zz_17_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h12 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_17_t = ( ( { 9{ RG_zz_17_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_17_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_17_en = ( RG_zz_17_t_c1 | RG_zz_17_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_17_en )
		RG_zz_17 <= RG_zz_17_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_173 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_18_t_c1 = ( U_05 & M_173 ) ;	// line#=../rle.cpp:111
	RG_zz_18_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h13 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_18_t = ( ( { 9{ RG_zz_18_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_18_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_18_en = ( RG_zz_18_t_c1 | RG_zz_18_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_18_en )
		RG_zz_18 <= RG_zz_18_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_172 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_19_t_c1 = ( U_05 & M_172 ) ;	// line#=../rle.cpp:111
	RG_zz_19_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h14 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_19_t = ( ( { 9{ RG_zz_19_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_19_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_19_en = ( RG_zz_19_t_c1 | RG_zz_19_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_19_en )
		RG_zz_19 <= RG_zz_19_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_171 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_20_t_c1 = ( U_05 & M_171 ) ;	// line#=../rle.cpp:111
	RG_zz_20_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h15 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_20_t = ( ( { 9{ RG_zz_20_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_20_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_20_en = ( RG_zz_20_t_c1 | RG_zz_20_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_20_en )
		RG_zz_20 <= RG_zz_20_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_170 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_21_t_c1 = ( U_05 & M_170 ) ;	// line#=../rle.cpp:111
	RG_zz_21_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h16 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_21_t = ( ( { 9{ RG_zz_21_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_21_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_21_en = ( RG_zz_21_t_c1 | RG_zz_21_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_21_en )
		RG_zz_21 <= RG_zz_21_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_169 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_22_t_c1 = ( U_05 & M_169 ) ;	// line#=../rle.cpp:111
	RG_zz_22_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h17 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_22_t = ( ( { 9{ RG_zz_22_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_22_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_22_en = ( RG_zz_22_t_c1 | RG_zz_22_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_22_en )
		RG_zz_22 <= RG_zz_22_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_168 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_23_t_c1 = ( U_05 & M_168 ) ;	// line#=../rle.cpp:111
	RG_zz_23_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h18 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_23_t = ( ( { 9{ RG_zz_23_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_23_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_23_en = ( RG_zz_23_t_c1 | RG_zz_23_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_23_en )
		RG_zz_23 <= RG_zz_23_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_167 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_24_t_c1 = ( U_05 & M_167 ) ;	// line#=../rle.cpp:111
	RG_zz_24_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h19 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_24_t = ( ( { 9{ RG_zz_24_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_24_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_24_en = ( RG_zz_24_t_c1 | RG_zz_24_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_24_en )
		RG_zz_24 <= RG_zz_24_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_166 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_25_t_c1 = ( U_05 & M_166 ) ;	// line#=../rle.cpp:111
	RG_zz_25_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h1a ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_25_t = ( ( { 9{ RG_zz_25_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_25_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_25_en = ( RG_zz_25_t_c1 | RG_zz_25_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_25_en )
		RG_zz_25 <= RG_zz_25_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_165 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_26_t_c1 = ( U_05 & M_165 ) ;	// line#=../rle.cpp:111
	RG_zz_26_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h1b ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_26_t = ( ( { 9{ RG_zz_26_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_26_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_26_en = ( RG_zz_26_t_c1 | RG_zz_26_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_26_en )
		RG_zz_26 <= RG_zz_26_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_164 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_27_t_c1 = ( U_05 & M_164 ) ;	// line#=../rle.cpp:111
	RG_zz_27_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h1c ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_27_t = ( ( { 9{ RG_zz_27_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_27_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_27_en = ( RG_zz_27_t_c1 | RG_zz_27_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_27_en )
		RG_zz_27 <= RG_zz_27_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_163 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_28_t_c1 = ( U_05 & M_163 ) ;	// line#=../rle.cpp:111
	RG_zz_28_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h1d ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_28_t = ( ( { 9{ RG_zz_28_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_28_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_28_en = ( RG_zz_28_t_c1 | RG_zz_28_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_28_en )
		RG_zz_28 <= RG_zz_28_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_162 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_29_t_c1 = ( U_05 & M_162 ) ;	// line#=../rle.cpp:111
	RG_zz_29_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h1e ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_29_t = ( ( { 9{ RG_zz_29_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_29_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_29_en = ( RG_zz_29_t_c1 | RG_zz_29_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_29_en )
		RG_zz_29 <= RG_zz_29_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_161 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_30_t_c1 = ( U_05 & M_161 ) ;	// line#=../rle.cpp:111
	RG_zz_30_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h1f ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_30_t = ( ( { 9{ RG_zz_30_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_30_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_30_en = ( RG_zz_30_t_c1 | RG_zz_30_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_30_en )
		RG_zz_30 <= RG_zz_30_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_160 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_31_t_c1 = ( U_05 & M_160 ) ;	// line#=../rle.cpp:111
	RG_zz_31_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h20 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_31_t = ( ( { 9{ RG_zz_31_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_31_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_31_en = ( RG_zz_31_t_c1 | RG_zz_31_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_31_en )
		RG_zz_31 <= RG_zz_31_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_159 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_32_t_c1 = ( U_05 & M_159 ) ;	// line#=../rle.cpp:111
	RG_zz_32_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h21 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_32_t = ( ( { 9{ RG_zz_32_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_32_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_32_en = ( RG_zz_32_t_c1 | RG_zz_32_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_32_en )
		RG_zz_32 <= RG_zz_32_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_158 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_33_t_c1 = ( U_05 & M_158 ) ;	// line#=../rle.cpp:111
	RG_zz_33_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h22 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_33_t = ( ( { 9{ RG_zz_33_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_33_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_33_en = ( RG_zz_33_t_c1 | RG_zz_33_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_33_en )
		RG_zz_33 <= RG_zz_33_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_157 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_34_t_c1 = ( U_05 & M_157 ) ;	// line#=../rle.cpp:111
	RG_zz_34_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h23 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_34_t = ( ( { 9{ RG_zz_34_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_34_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_34_en = ( RG_zz_34_t_c1 | RG_zz_34_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_34_en )
		RG_zz_34 <= RG_zz_34_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_115 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_35_t_c1 = ( U_05 & M_115 ) ;	// line#=../rle.cpp:111
	RG_zz_35_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h24 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_35_t = ( ( { 9{ RG_zz_35_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_35_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_35_en = ( RG_zz_35_t_c1 | RG_zz_35_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_35_en )
		RG_zz_35 <= RG_zz_35_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_156 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_36_t_c1 = ( U_05 & M_156 ) ;	// line#=../rle.cpp:111
	RG_zz_36_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h25 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_36_t = ( ( { 9{ RG_zz_36_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_36_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_36_en = ( RG_zz_36_t_c1 | RG_zz_36_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_36_en )
		RG_zz_36 <= RG_zz_36_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_155 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_37_t_c1 = ( U_05 & M_155 ) ;	// line#=../rle.cpp:111
	RG_zz_37_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h26 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_37_t = ( ( { 9{ RG_zz_37_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_37_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_37_en = ( RG_zz_37_t_c1 | RG_zz_37_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_37_en )
		RG_zz_37 <= RG_zz_37_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_154 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_38_t_c1 = ( U_05 & M_154 ) ;	// line#=../rle.cpp:111
	RG_zz_38_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h27 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_38_t = ( ( { 9{ RG_zz_38_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_38_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_38_en = ( RG_zz_38_t_c1 | RG_zz_38_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_38_en )
		RG_zz_38 <= RG_zz_38_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_153 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_39_t_c1 = ( U_05 & M_153 ) ;	// line#=../rle.cpp:111
	RG_zz_39_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h28 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_39_t = ( ( { 9{ RG_zz_39_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_39_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_39_en = ( RG_zz_39_t_c1 | RG_zz_39_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_39_en )
		RG_zz_39 <= RG_zz_39_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_152 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_40_t_c1 = ( U_05 & M_152 ) ;	// line#=../rle.cpp:111
	RG_zz_40_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h29 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_40_t = ( ( { 9{ RG_zz_40_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_40_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_40_en = ( RG_zz_40_t_c1 | RG_zz_40_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_40_en )
		RG_zz_40 <= RG_zz_40_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_151 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_41_t_c1 = ( U_05 & M_151 ) ;	// line#=../rle.cpp:111
	RG_zz_41_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h2a ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_41_t = ( ( { 9{ RG_zz_41_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_41_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_41_en = ( RG_zz_41_t_c1 | RG_zz_41_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_41_en )
		RG_zz_41 <= RG_zz_41_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_150 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_42_t_c1 = ( U_05 & M_150 ) ;	// line#=../rle.cpp:111
	RG_zz_42_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h2b ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_42_t = ( ( { 9{ RG_zz_42_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_42_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_42_en = ( RG_zz_42_t_c1 | RG_zz_42_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_42_en )
		RG_zz_42 <= RG_zz_42_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_149 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_43_t_c1 = ( U_05 & M_149 ) ;	// line#=../rle.cpp:111
	RG_zz_43_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h2c ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_43_t = ( ( { 9{ RG_zz_43_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_43_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_43_en = ( RG_zz_43_t_c1 | RG_zz_43_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_43_en )
		RG_zz_43 <= RG_zz_43_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_148 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_44_t_c1 = ( U_05 & M_148 ) ;	// line#=../rle.cpp:111
	RG_zz_44_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h2d ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_44_t = ( ( { 9{ RG_zz_44_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_44_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_44_en = ( RG_zz_44_t_c1 | RG_zz_44_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_44_en )
		RG_zz_44 <= RG_zz_44_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_147 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_45_t_c1 = ( U_05 & M_147 ) ;	// line#=../rle.cpp:111
	RG_zz_45_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h2e ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_45_t = ( ( { 9{ RG_zz_45_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_45_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_45_en = ( RG_zz_45_t_c1 | RG_zz_45_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_45_en )
		RG_zz_45 <= RG_zz_45_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_146 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_46_t_c1 = ( U_05 & M_146 ) ;	// line#=../rle.cpp:111
	RG_zz_46_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h2f ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_46_t = ( ( { 9{ RG_zz_46_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_46_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_46_en = ( RG_zz_46_t_c1 | RG_zz_46_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_46_en )
		RG_zz_46 <= RG_zz_46_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_145 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_47_t_c1 = ( U_05 & M_145 ) ;	// line#=../rle.cpp:111
	RG_zz_47_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h30 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_47_t = ( ( { 9{ RG_zz_47_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_47_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_47_en = ( RG_zz_47_t_c1 | RG_zz_47_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_47_en )
		RG_zz_47 <= RG_zz_47_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_144 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_48_t_c1 = ( U_05 & M_144 ) ;	// line#=../rle.cpp:111
	RG_zz_48_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h31 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_48_t = ( ( { 9{ RG_zz_48_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_48_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_48_en = ( RG_zz_48_t_c1 | RG_zz_48_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_48_en )
		RG_zz_48 <= RG_zz_48_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_143 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_49_t_c1 = ( U_05 & M_143 ) ;	// line#=../rle.cpp:111
	RG_zz_49_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h32 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_49_t = ( ( { 9{ RG_zz_49_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_49_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_49_en = ( RG_zz_49_t_c1 | RG_zz_49_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_49_en )
		RG_zz_49 <= RG_zz_49_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_142 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_50_t_c1 = ( U_05 & M_142 ) ;	// line#=../rle.cpp:111
	RG_zz_50_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h33 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_50_t = ( ( { 9{ RG_zz_50_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_50_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_50_en = ( RG_zz_50_t_c1 | RG_zz_50_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_50_en )
		RG_zz_50 <= RG_zz_50_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_141 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_51_t_c1 = ( U_05 & M_141 ) ;	// line#=../rle.cpp:111
	RG_zz_51_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h34 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_51_t = ( ( { 9{ RG_zz_51_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_51_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_51_en = ( RG_zz_51_t_c1 | RG_zz_51_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_51_en )
		RG_zz_51 <= RG_zz_51_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_140 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_52_t_c1 = ( U_05 & M_140 ) ;	// line#=../rle.cpp:111
	RG_zz_52_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h35 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_52_t = ( ( { 9{ RG_zz_52_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_52_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_52_en = ( RG_zz_52_t_c1 | RG_zz_52_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_52_en )
		RG_zz_52 <= RG_zz_52_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_139 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_53_t_c1 = ( U_05 & M_139 ) ;	// line#=../rle.cpp:111
	RG_zz_53_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h36 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_53_t = ( ( { 9{ RG_zz_53_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_53_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_53_en = ( RG_zz_53_t_c1 | RG_zz_53_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_53_en )
		RG_zz_53 <= RG_zz_53_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_138 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_54_t_c1 = ( U_05 & M_138 ) ;	// line#=../rle.cpp:111
	RG_zz_54_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h37 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_54_t = ( ( { 9{ RG_zz_54_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_54_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_54_en = ( RG_zz_54_t_c1 | RG_zz_54_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_54_en )
		RG_zz_54 <= RG_zz_54_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_137 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_55_t_c1 = ( U_05 & M_137 ) ;	// line#=../rle.cpp:111
	RG_zz_55_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h38 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_55_t = ( ( { 9{ RG_zz_55_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_55_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_55_en = ( RG_zz_55_t_c1 | RG_zz_55_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_55_en )
		RG_zz_55 <= RG_zz_55_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_136 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_56_t_c1 = ( U_05 & M_136 ) ;	// line#=../rle.cpp:111
	RG_zz_56_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h39 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_56_t = ( ( { 9{ RG_zz_56_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_56_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_56_en = ( RG_zz_56_t_c1 | RG_zz_56_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_56_en )
		RG_zz_56 <= RG_zz_56_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_135 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_57_t_c1 = ( U_05 & M_135 ) ;	// line#=../rle.cpp:111
	RG_zz_57_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h3a ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_57_t = ( ( { 9{ RG_zz_57_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_57_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_57_en = ( RG_zz_57_t_c1 | RG_zz_57_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_57_en )
		RG_zz_57 <= RG_zz_57_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_134 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_58_t_c1 = ( U_05 & M_134 ) ;	// line#=../rle.cpp:111
	RG_zz_58_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h3b ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_58_t = ( ( { 9{ RG_zz_58_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_58_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_58_en = ( RG_zz_58_t_c1 | RG_zz_58_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_58_en )
		RG_zz_58 <= RG_zz_58_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_133 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_59_t_c1 = ( U_05 & M_133 ) ;	// line#=../rle.cpp:111
	RG_zz_59_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h3c ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_59_t = ( ( { 9{ RG_zz_59_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_59_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_59_en = ( RG_zz_59_t_c1 | RG_zz_59_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_59_en )
		RG_zz_59 <= RG_zz_59_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_132 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_60_t_c1 = ( U_05 & M_132 ) ;	// line#=../rle.cpp:111
	RG_zz_60_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h3d ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_60_t = ( ( { 9{ RG_zz_60_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_60_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_60_en = ( RG_zz_60_t_c1 | RG_zz_60_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_60_en )
		RG_zz_60 <= RG_zz_60_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_131 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_61_t_c1 = ( U_05 & M_131 ) ;	// line#=../rle.cpp:111
	RG_zz_61_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h3e ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_61_t = ( ( { 9{ RG_zz_61_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_61_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_61_en = ( RG_zz_61_t_c1 | RG_zz_61_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_61_en )
		RG_zz_61 <= RG_zz_61_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_01 or U_87 or M_217 or M_130 or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_62_t_c1 = ( U_05 & M_130 ) ;	// line#=../rle.cpp:111
	RG_zz_62_t_c2 = ( U_87 & ( ~|( RG_k_01 [5:0] ^ 6'h3f ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_62_t = ( ( { 9{ RG_zz_62_t_c1 } } & M_217 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_62_t_c2 } } & M_217 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_62_en = ( RG_zz_62_t_c1 | RG_zz_62_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_62_en )
		RG_zz_62 <= RG_zz_62_t ;	// line#=../rle.cpp:111,142
always @ ( FF_j or U_254 or incr4s1ot or ST1_02d or ST1_01d )
	RG_j_03_t = ( ( { 4{ ST1_01d } } & 4'hf /*-4'h1*/ )	// line#=../rle.cpp:34
		| ( { 4{ ST1_02d } } & incr4s1ot )		// line#=../rle.cpp:34
		| ( { 4{ U_254 } } & { 3'h0 , FF_j } )		// line#=../rle.cpp:83,84
		) ;
assign	RG_j_03_en = ( ST1_01d | ST1_02d | U_254 ) ;
always @ ( posedge clk )
	if ( RG_j_03_en )
		RG_j_03 <= RG_j_03_t ;	// line#=../rle.cpp:34,83,84
assign	M_186 = ( ST1_02d | U_88 ) ;
always @ ( U_06 or FF_i or U_88 or M_186 )
	TR_01 = ( ( { 3{ M_186 } } & { 2'h0 , ( U_88 & FF_i ) } )	// line#=../rle.cpp:105
		| ( { 3{ U_06 } } & 3'h7 )				// line#=../rle.cpp:134
		) ;
always @ ( decr32s1ot or U_165 or U_83 or incr32s2ot or U_169 or U_177 or U_166 or 
	U_163 or U_84 or U_81 or TR_01 or U_88 or M_185 )
	begin
	RG_i_t_c1 = ( M_185 | U_88 ) ;	// line#=../rle.cpp:105,134
	RG_i_t_c2 = ( ( ( ( ( U_81 | U_84 ) | U_163 ) | U_166 ) | U_177 ) | U_169 ) ;	// line#=../rle.cpp:63,74,119,129,150,160
	RG_i_t_c3 = ( U_83 | U_165 ) ;	// line#=../rle.cpp:124,155
	RG_i_t = ( ( { 32{ RG_i_t_c1 } } & { 29'h00000000 , TR_01 } )	// line#=../rle.cpp:105,134
		| ( { 32{ RG_i_t_c2 } } & incr32s2ot )			// line#=../rle.cpp:63,74,119,129,150,160
		| ( { 32{ RG_i_t_c3 } } & decr32s1ot )			// line#=../rle.cpp:124,155
		) ;
	end
assign	RG_i_en = ( RG_i_t_c1 | RG_i_t_c2 | RG_i_t_c3 ) ;
always @ ( posedge clk )
	if ( RG_i_en )
		RG_i <= RG_i_t ;	// line#=../rle.cpp:63,74,105,119,124,129
					// ,134,150,155,160
always @ ( decr32s2ot or U_166 or U_84 or incr32s1ot or U_169 or U_165 or U_161 or 
	U_83 or U_79 or U_06 or ST1_07d or M_186 )
	begin
	RG_j_k_t_c1 = ( ( M_186 | ST1_07d ) | U_06 ) ;	// line#=../rle.cpp:59,105,135
	RG_j_k_t_c2 = ( ( ( ( U_79 | U_83 ) | U_161 ) | U_165 ) | U_169 ) ;	// line#=../rle.cpp:64,114,125,145,156
	RG_j_k_t_c3 = ( U_84 | U_166 ) ;	// line#=../rle.cpp:130,161
	RG_j_k_t = ( ( { 32{ RG_j_k_t_c1 } } & { 31'h00000000 , U_06 } )	// line#=../rle.cpp:59,105,135
		| ( { 32{ RG_j_k_t_c2 } } & incr32s1ot )			// line#=../rle.cpp:64,114,125,145,156
		| ( { 32{ RG_j_k_t_c3 } } & decr32s2ot )			// line#=../rle.cpp:130,161
		) ;
	end
assign	RG_j_k_en = ( RG_j_k_t_c1 | RG_j_k_t_c2 | RG_j_k_t_c3 ) ;
always @ ( posedge clk )
	if ( RG_j_k_en )
		RG_j_k <= RG_j_k_t ;	// line#=../rle.cpp:59,64,105,114,125,130
					// ,135,145,156,161
assign	RG_quantized_block_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_en )
		RG_quantized_block <= jpeg_in_a00 ;
assign	RG_quantized_block_1_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_1_en )
		RG_quantized_block_1 <= jpeg_in_a01 ;
assign	RG_quantized_block_2_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_2_en )
		RG_quantized_block_2 <= jpeg_in_a02 ;
assign	RG_quantized_block_3_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_3_en )
		RG_quantized_block_3 <= jpeg_in_a03 ;
assign	RG_quantized_block_4_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_4_en )
		RG_quantized_block_4 <= jpeg_in_a04 ;
assign	RG_quantized_block_5_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_5_en )
		RG_quantized_block_5 <= jpeg_in_a05 ;
assign	RG_quantized_block_6_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_6_en )
		RG_quantized_block_6 <= jpeg_in_a06 ;
assign	RG_quantized_block_7_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_7_en )
		RG_quantized_block_7 <= jpeg_in_a07 ;
assign	RG_quantized_block_8_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_8_en )
		RG_quantized_block_8 <= jpeg_in_a08 ;
assign	RG_quantized_block_9_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_9_en )
		RG_quantized_block_9 <= jpeg_in_a09 ;
assign	RG_quantized_block_10_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_10_en )
		RG_quantized_block_10 <= jpeg_in_a10 ;
assign	RG_quantized_block_11_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_11_en )
		RG_quantized_block_11 <= jpeg_in_a11 ;
assign	RG_quantized_block_12_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_12_en )
		RG_quantized_block_12 <= jpeg_in_a12 ;
assign	RG_quantized_block_13_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_13_en )
		RG_quantized_block_13 <= jpeg_in_a13 ;
assign	RG_quantized_block_14_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_14_en )
		RG_quantized_block_14 <= jpeg_in_a14 ;
assign	RG_quantized_block_15_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_15_en )
		RG_quantized_block_15 <= jpeg_in_a15 ;
assign	RG_quantized_block_16_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_16_en )
		RG_quantized_block_16 <= jpeg_in_a16 ;
assign	RG_quantized_block_17_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_17_en )
		RG_quantized_block_17 <= jpeg_in_a17 ;
assign	RG_quantized_block_18_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_18_en )
		RG_quantized_block_18 <= jpeg_in_a18 ;
assign	RG_quantized_block_19_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_19_en )
		RG_quantized_block_19 <= jpeg_in_a19 ;
assign	RG_quantized_block_20_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_20_en )
		RG_quantized_block_20 <= jpeg_in_a20 ;
assign	RG_quantized_block_21_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_21_en )
		RG_quantized_block_21 <= jpeg_in_a21 ;
assign	RG_quantized_block_22_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_22_en )
		RG_quantized_block_22 <= jpeg_in_a22 ;
assign	RG_quantized_block_23_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_23_en )
		RG_quantized_block_23 <= jpeg_in_a23 ;
assign	RG_quantized_block_24_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_24_en )
		RG_quantized_block_24 <= jpeg_in_a24 ;
assign	RG_quantized_block_25_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_25_en )
		RG_quantized_block_25 <= jpeg_in_a25 ;
assign	RG_quantized_block_26_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_26_en )
		RG_quantized_block_26 <= jpeg_in_a26 ;
assign	RG_quantized_block_27_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_27_en )
		RG_quantized_block_27 <= jpeg_in_a27 ;
assign	RG_quantized_block_28_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_28_en )
		RG_quantized_block_28 <= jpeg_in_a28 ;
assign	RG_quantized_block_29_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_29_en )
		RG_quantized_block_29 <= jpeg_in_a29 ;
assign	RG_quantized_block_30_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_30_en )
		RG_quantized_block_30 <= jpeg_in_a30 ;
assign	RG_quantized_block_31_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_31_en )
		RG_quantized_block_31 <= jpeg_in_a31 ;
assign	RG_quantized_block_32_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_32_en )
		RG_quantized_block_32 <= jpeg_in_a32 ;
assign	RG_quantized_block_33_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_33_en )
		RG_quantized_block_33 <= jpeg_in_a33 ;
assign	RG_quantized_block_34_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_34_en )
		RG_quantized_block_34 <= jpeg_in_a34 ;
assign	RG_quantized_block_35_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_35_en )
		RG_quantized_block_35 <= jpeg_in_a35 ;
assign	RG_quantized_block_36_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_36_en )
		RG_quantized_block_36 <= jpeg_in_a36 ;
assign	RG_quantized_block_37_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_37_en )
		RG_quantized_block_37 <= jpeg_in_a37 ;
assign	RG_quantized_block_38_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_38_en )
		RG_quantized_block_38 <= jpeg_in_a38 ;
assign	RG_quantized_block_39_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_39_en )
		RG_quantized_block_39 <= jpeg_in_a39 ;
assign	RG_quantized_block_40_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_40_en )
		RG_quantized_block_40 <= jpeg_in_a40 ;
assign	RG_quantized_block_41_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_41_en )
		RG_quantized_block_41 <= jpeg_in_a41 ;
assign	RG_quantized_block_42_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_42_en )
		RG_quantized_block_42 <= jpeg_in_a42 ;
assign	RG_quantized_block_43_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_43_en )
		RG_quantized_block_43 <= jpeg_in_a43 ;
assign	RG_quantized_block_44_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_44_en )
		RG_quantized_block_44 <= jpeg_in_a44 ;
assign	RG_quantized_block_45_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_45_en )
		RG_quantized_block_45 <= jpeg_in_a45 ;
assign	RG_quantized_block_46_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_46_en )
		RG_quantized_block_46 <= jpeg_in_a46 ;
assign	RG_quantized_block_47_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_47_en )
		RG_quantized_block_47 <= jpeg_in_a47 ;
assign	RG_quantized_block_48_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_48_en )
		RG_quantized_block_48 <= jpeg_in_a48 ;
assign	RG_quantized_block_49_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_49_en )
		RG_quantized_block_49 <= jpeg_in_a49 ;
assign	RG_quantized_block_50_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_50_en )
		RG_quantized_block_50 <= jpeg_in_a50 ;
assign	RG_quantized_block_51_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_51_en )
		RG_quantized_block_51 <= jpeg_in_a51 ;
assign	RG_quantized_block_52_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_52_en )
		RG_quantized_block_52 <= jpeg_in_a52 ;
assign	RG_quantized_block_53_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_53_en )
		RG_quantized_block_53 <= jpeg_in_a53 ;
assign	RG_quantized_block_54_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_54_en )
		RG_quantized_block_54 <= jpeg_in_a54 ;
assign	RG_quantized_block_55_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_55_en )
		RG_quantized_block_55 <= jpeg_in_a55 ;
assign	RG_quantized_block_56_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_56_en )
		RG_quantized_block_56 <= jpeg_in_a56 ;
assign	RG_quantized_block_57_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_57_en )
		RG_quantized_block_57 <= jpeg_in_a57 ;
assign	RG_quantized_block_58_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_58_en )
		RG_quantized_block_58 <= jpeg_in_a58 ;
assign	RG_quantized_block_59_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_59_en )
		RG_quantized_block_59 <= jpeg_in_a59 ;
assign	RG_quantized_block_60_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_60_en )
		RG_quantized_block_60 <= jpeg_in_a60 ;
jpeg_MEM_rl rl ( .AD1(rl_AD1) ,.RD1(rl_RD1) ,.WD1(rl_WD1) ,.WE1(rl_WE1) ,.CLK1(clk) ,
	.RA2(rl_RA2) ,.RD2(rl_RD2) ,.RA3(rl_RA3) ,.RD3(rl_RD3) );	// line#=../rle.cpp:23
always @ ( rl_RD2 or M_188 or jpeg_in_a61 or ST1_02d )
	RG_quantized_block_rl_02_t = ( ( { 9{ ST1_02d } } & jpeg_in_a61 )	// line#=../rle.cpp:45
		| ( { 9{ M_188 } } & rl_RD2 ) ) ;
assign	RG_quantized_block_rl_02_en = ( ST1_02d | M_188 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_02_en )
		RG_quantized_block_rl_02 <= RG_quantized_block_rl_02_t ;	// line#=../rle.cpp:45
assign	M_188 = ( ST1_08d | ( ST1_11d & FL01_02_01a ) ) ;
always @ ( rl_RD3 or M_188 or jpeg_in_a62 or ST1_02d )
	RG_quantized_block_rl_02_1_t = ( ( { 9{ ST1_02d } } & jpeg_in_a62 )	// line#=../rle.cpp:45
		| ( { 9{ M_188 } } & rl_RD3 )					// line#=../rle.cpp:77,78,83,84
		) ;
assign	RG_quantized_block_rl_02_1_en = ( ST1_02d | M_188 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_02_1_en )
		RG_quantized_block_rl_02_1 <= RG_quantized_block_rl_02_1_t ;	// line#=../rle.cpp:45,77,78,83,84
always @ ( RG_previous_dc_zz or U_88 or jpeg_in_a63 or ST1_02d )
	RG_quantized_block_zz_t = ( ( { 9{ ST1_02d } } & jpeg_in_a63 )	// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_previous_dc_zz ) ) ;
assign	RG_quantized_block_zz_en = ( ST1_02d | U_88 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_zz_en )
		RG_quantized_block_zz <= RG_quantized_block_zz_t ;	// line#=../rle.cpp:45
always @ ( RG_i or ST1_06d or incr8u2ot or ST1_03d )
	RG_k_t = ( ( { 6{ ST1_03d } } & incr8u2ot [5:0] )	// line#=../rle.cpp:111
		| ( { 6{ ST1_06d } } & RG_i [5:0] )		// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:105
always @ ( posedge clk )
	RG_k <= RG_k_t ;	// line#=../rle.cpp:74,105,111
assign	M_185 = ( ST1_02d | U_06 ) ;
always @ ( M_02_t1 or ST1_09d or U_163 or U_79 or U_161 or U_81 or M_185 )
	begin
	FF_d_t_c1 = ( ( M_185 | U_81 ) | U_161 ) ;	// line#=../rle.cpp:105,120,136,146
	FF_d_t_c2 = ( U_79 | U_163 ) ;	// line#=../rle.cpp:115,151
	FF_d_t = ( ( { 1{ FF_d_t_c2 } } & 1'h1 )	// line#=../rle.cpp:115,151
		| ( { 1{ ST1_09d } } & ( ~M_02_t1 ) )	// line#=../rle.cpp:77,78
		) ;	// line#=../rle.cpp:105,120,136,146
	end
assign	FF_d_en = ( FF_d_t_c1 | FF_d_t_c2 | ST1_09d ) ;
always @ ( posedge clk )
	if ( FF_d_en )
		FF_d <= FF_d_t ;	// line#=../rle.cpp:77,78,105,115,120,136
					// ,146,151
assign	FF_j_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:36
	if ( FF_j_en )
		FF_j <= 1'h0 ;
always @ ( CT_35 or ST1_07d or CT_33 or ST1_06d or ST1_02d )
	FF_i_t = ( ( { 1{ ST1_02d } } & 1'h1 )	// line#=../rle.cpp:37
		| ( { 1{ ST1_06d } } & CT_33 )	// line#=../rle.cpp:66,67
		| ( { 1{ ST1_07d } } & CT_35 )	// line#=../rle.cpp:57,58
		) ;
assign	FF_i_en = ( ST1_02d | ST1_06d | ST1_07d ) ;
always @ ( posedge clk )
	if ( FF_i_en )
		FF_i <= FF_i_t ;	// line#=../rle.cpp:37,57,58,66,67
always @ ( RG_136 or ST1_06d or ST1_02d )
	FF_len_t = ( ( { 1{ ST1_02d } } & 1'h1 )	// line#=../rle.cpp:39
		| ( { 1{ ST1_06d } } & RG_136 ) ) ;
assign	FF_len_en = ( ST1_02d | ST1_06d ) ;
always @ ( posedge clk )
	if ( FF_len_en )
		FF_len <= FF_len_t ;	// line#=../rle.cpp:39
assign	RG_len_03_en = U_254 ;
always @ ( posedge clk )
	if ( RG_len_03_en )
		RG_len_03 <= RG_len_02 ;
always @ ( sub8u_71ot or U_252 or decr8u_71ot or ST1_07d )
	RG_142_01_t = ( ( { 7{ ST1_07d } } & decr8u_71ot )	// line#=../rle.cpp:77,78
		| ( { 7{ U_252 } } & sub8u_71ot )		// line#=../rle.cpp:83,84
		) ;
always @ ( posedge clk )
	RG_142_01 <= RG_142_01_t ;	// line#=../rle.cpp:77,78,83,84
always @ ( sub8u1ot or U_252 or incr8u2ot or ST1_10d or ST1_07d or FF_len or ST1_04d )
	begin
	RG_len_01_1_t_c1 = ( ST1_07d | ST1_10d ) ;	// line#=../rle.cpp:69,74,80
	RG_len_01_1_t = ( ( { 8{ ST1_04d } } & { 7'h00 , FF_len } )
		| ( { 8{ RG_len_01_1_t_c1 } } & incr8u2ot )	// line#=../rle.cpp:69,74,80
		| ( { 8{ U_252 } } & sub8u1ot )			// line#=../rle.cpp:83,84,86
		) ;
	end
assign	RG_len_01_1_en = ( ST1_04d | RG_len_01_1_t_c1 | U_252 ) ;
always @ ( posedge clk )
	if ( RG_len_01_1_en )
		RG_len_01_1 <= RG_len_01_1_t ;	// line#=../rle.cpp:69,74,80,83,84,86
always @ ( sub8u_7_11ot or U_252 or ST1_07d or incr8u2ot or ST1_04d or RG_k or ST1_03d )
	begin
	RG_k_01_t_c1 = ( ST1_07d | U_252 ) ;	// line#=../rle.cpp:77,78,83,84
	RG_k_01_t = ( ( { 7{ ST1_03d } } & { 1'h0 , RG_k } )
		| ( { 7{ ST1_04d } } & incr8u2ot [6:0] )	// line#=../rle.cpp:142
		| ( { 7{ RG_k_01_t_c1 } } & sub8u_7_11ot )	// line#=../rle.cpp:77,78,83,84
		) ;
	end
always @ ( posedge clk )
	RG_k_01 <= RG_k_01_t ;	// line#=../rle.cpp:77,78,83,84,142
assign	JF_01 = ~( ~|{ ~incr4s1ot [3] , incr4s1ot [2:0] } ) ;	// line#=../rle.cpp:34,35
always @ ( RG_quantized_block_7 or RG_quantized_block_6 or RG_quantized_block_5 or 
	RG_quantized_block_4 or RG_quantized_block_3 or RG_quantized_block_2 or 
	RG_quantized_block_1 or RG_quantized_block or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_44 = RG_quantized_block ;	// line#=../rle.cpp:111
	3'h1 :
		TR_44 = RG_quantized_block_1 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_44 = RG_quantized_block_2 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_44 = RG_quantized_block_3 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_44 = RG_quantized_block_4 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_44 = RG_quantized_block_5 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_44 = RG_quantized_block_6 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_44 = RG_quantized_block_7 ;	// line#=../rle.cpp:111
	default :
		TR_44 = 9'hx ;
	endcase
always @ ( RG_quantized_block_15 or RG_quantized_block_14 or RG_quantized_block_13 or 
	RG_quantized_block_12 or RG_quantized_block_11 or RG_quantized_block_10 or 
	RG_quantized_block_9 or RG_quantized_block_8 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_45 = RG_quantized_block_8 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_45 = RG_quantized_block_9 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_45 = RG_quantized_block_10 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_45 = RG_quantized_block_11 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_45 = RG_quantized_block_12 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_45 = RG_quantized_block_13 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_45 = RG_quantized_block_14 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_45 = RG_quantized_block_15 ;	// line#=../rle.cpp:111
	default :
		TR_45 = 9'hx ;
	endcase
always @ ( RG_quantized_block_23 or RG_quantized_block_22 or RG_quantized_block_21 or 
	RG_quantized_block_20 or RG_quantized_block_19 or RG_quantized_block_18 or 
	RG_quantized_block_17 or RG_quantized_block_16 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_46 = RG_quantized_block_16 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_46 = RG_quantized_block_17 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_46 = RG_quantized_block_18 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_46 = RG_quantized_block_19 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_46 = RG_quantized_block_20 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_46 = RG_quantized_block_21 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_46 = RG_quantized_block_22 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_46 = RG_quantized_block_23 ;	// line#=../rle.cpp:111
	default :
		TR_46 = 9'hx ;
	endcase
always @ ( RG_quantized_block_31 or RG_quantized_block_30 or RG_quantized_block_29 or 
	RG_quantized_block_28 or RG_quantized_block_27 or RG_quantized_block_26 or 
	RG_quantized_block_25 or RG_quantized_block_24 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_47 = RG_quantized_block_24 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_47 = RG_quantized_block_25 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_47 = RG_quantized_block_26 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_47 = RG_quantized_block_27 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_47 = RG_quantized_block_28 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_47 = RG_quantized_block_29 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_47 = RG_quantized_block_30 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_47 = RG_quantized_block_31 ;	// line#=../rle.cpp:111
	default :
		TR_47 = 9'hx ;
	endcase
always @ ( RG_quantized_block_39 or RG_quantized_block_38 or RG_quantized_block_37 or 
	RG_quantized_block_36 or RG_quantized_block_35 or RG_quantized_block_34 or 
	RG_quantized_block_33 or RG_quantized_block_32 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_48 = RG_quantized_block_32 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_48 = RG_quantized_block_33 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_48 = RG_quantized_block_34 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_48 = RG_quantized_block_35 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_48 = RG_quantized_block_36 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_48 = RG_quantized_block_37 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_48 = RG_quantized_block_38 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_48 = RG_quantized_block_39 ;	// line#=../rle.cpp:111
	default :
		TR_48 = 9'hx ;
	endcase
always @ ( RG_quantized_block_47 or RG_quantized_block_46 or RG_quantized_block_45 or 
	RG_quantized_block_44 or RG_quantized_block_43 or RG_quantized_block_42 or 
	RG_quantized_block_41 or RG_quantized_block_40 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_49 = RG_quantized_block_40 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_49 = RG_quantized_block_41 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_49 = RG_quantized_block_42 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_49 = RG_quantized_block_43 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_49 = RG_quantized_block_44 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_49 = RG_quantized_block_45 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_49 = RG_quantized_block_46 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_49 = RG_quantized_block_47 ;	// line#=../rle.cpp:111
	default :
		TR_49 = 9'hx ;
	endcase
always @ ( RG_quantized_block_55 or RG_quantized_block_54 or RG_quantized_block_53 or 
	RG_quantized_block_52 or RG_quantized_block_51 or RG_quantized_block_50 or 
	RG_quantized_block_49 or RG_quantized_block_48 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_50 = RG_quantized_block_48 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_50 = RG_quantized_block_49 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_50 = RG_quantized_block_50 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_50 = RG_quantized_block_51 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_50 = RG_quantized_block_52 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_50 = RG_quantized_block_53 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_50 = RG_quantized_block_54 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_50 = RG_quantized_block_55 ;	// line#=../rle.cpp:111
	default :
		TR_50 = 9'hx ;
	endcase
always @ ( RG_quantized_block_zz or RG_quantized_block_rl_02_1 or RG_quantized_block_rl_02 or 
	RG_quantized_block_60 or RG_quantized_block_59 or RG_quantized_block_58 or 
	RG_quantized_block_57 or RG_quantized_block_56 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_51 = RG_quantized_block_56 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_51 = RG_quantized_block_57 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_51 = RG_quantized_block_58 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_51 = RG_quantized_block_59 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_51 = RG_quantized_block_60 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_51 = RG_quantized_block_rl_02 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_51 = RG_quantized_block_rl_02_1 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_51 = RG_quantized_block_zz ;	// line#=../rle.cpp:111
	default :
		TR_51 = 9'hx ;
	endcase
always @ ( TR_51 or TR_50 or TR_49 or TR_48 or TR_47 or TR_46 or TR_45 or TR_44 or 
	RG_i )	// line#=../rle.cpp:111,142
	begin
	M_217_c1 = ~|RG_i [2:0] ;	// line#=../rle.cpp:111,142
	M_217_c2 = ~|( RG_i [2:0] ^ 3'h1 ) ;	// line#=../rle.cpp:111,142
	M_217_c3 = ~|( RG_i [2:0] ^ 3'h2 ) ;	// line#=../rle.cpp:111,142
	M_217_c4 = ~|( RG_i [2:0] ^ 3'h3 ) ;	// line#=../rle.cpp:111,142
	M_217_c5 = ~|( RG_i [2:0] ^ 3'h4 ) ;	// line#=../rle.cpp:111,142
	M_217_c6 = ~|( RG_i [2:0] ^ 3'h5 ) ;	// line#=../rle.cpp:111,142
	M_217_c7 = ~|( RG_i [2:0] ^ 3'h6 ) ;	// line#=../rle.cpp:111,142
	M_217_c8 = ~|( RG_i [2:0] ^ 3'h7 ) ;	// line#=../rle.cpp:111,142
	M_217 = ( ( { 9{ M_217_c1 } } & TR_44 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_217_c2 } } & TR_45 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_217_c3 } } & TR_46 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_217_c4 } } & TR_47 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_217_c5 } } & TR_48 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_217_c6 } } & TR_49 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_217_c7 } } & TR_50 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_217_c8 } } & TR_51 )	// line#=../rle.cpp:111,142
		) ;
	end
assign	JF_03 = ~RG_k_01 [6] ;
always @ ( RG_zz_62 or RG_zz_61 or RG_zz_60 or RG_zz_59 or RG_zz_58 or RG_zz_57 or 
	RG_zz_56 or RG_zz_55 or RG_zz_54 or RG_zz_53 or RG_zz_52 or RG_zz_51 or 
	RG_zz_50 or RG_zz_49 or RG_zz_48 or RG_zz_47 or RG_zz_46 or RG_zz_45 or 
	RG_zz_44 or RG_zz_43 or RG_zz_42 or RG_zz_41 or RG_zz_40 or RG_zz_39 or 
	RG_zz_38 or RG_zz_37 or RG_zz_36 or RG_zz_35 or RG_zz_34 or RG_zz_33 or 
	RG_zz_32 or RG_zz_31 or RG_zz_30 or RG_zz_29 or RG_zz_28 or RG_zz_27 or 
	RG_zz_26 or RG_zz_25 or RG_zz_24 or RG_zz_23 or RG_zz_22 or RG_zz_21 or 
	RG_zz_20 or RG_zz_19 or RG_zz_18 or RG_zz_17 or RG_zz_16 or RG_zz_15 or 
	RG_zz_14 or RG_zz_13 or RG_zz_12 or RG_zz_11 or RG_zz_10 or RG_zz_9 or RG_zz_8 or 
	RG_zz_7 or RG_zz_6 or RG_zz_5 or RG_zz_4 or RG_zz_3 or RG_zz_2 or RG_zz_1 or 
	RG_zz or RG_quantized_block_zz or RG_i )	// line#=../rle.cpp:61,62
	case ( RG_i [5:0] )
	6'h00 :
		M_01_t64_t1 = ~|RG_quantized_block_zz ;	// line#=../rle.cpp:61,62
	6'h01 :
		M_01_t64_t1 = ~|RG_zz ;	// line#=../rle.cpp:61,62
	6'h02 :
		M_01_t64_t1 = ~|RG_zz_1 ;	// line#=../rle.cpp:61,62
	6'h03 :
		M_01_t64_t1 = ~|RG_zz_2 ;	// line#=../rle.cpp:61,62
	6'h04 :
		M_01_t64_t1 = ~|RG_zz_3 ;	// line#=../rle.cpp:61,62
	6'h05 :
		M_01_t64_t1 = ~|RG_zz_4 ;	// line#=../rle.cpp:61,62
	6'h06 :
		M_01_t64_t1 = ~|RG_zz_5 ;	// line#=../rle.cpp:61,62
	6'h07 :
		M_01_t64_t1 = ~|RG_zz_6 ;	// line#=../rle.cpp:61,62
	6'h08 :
		M_01_t64_t1 = ~|RG_zz_7 ;	// line#=../rle.cpp:61,62
	6'h09 :
		M_01_t64_t1 = ~|RG_zz_8 ;	// line#=../rle.cpp:61,62
	6'h0a :
		M_01_t64_t1 = ~|RG_zz_9 ;	// line#=../rle.cpp:61,62
	6'h0b :
		M_01_t64_t1 = ~|RG_zz_10 ;	// line#=../rle.cpp:61,62
	6'h0c :
		M_01_t64_t1 = ~|RG_zz_11 ;	// line#=../rle.cpp:61,62
	6'h0d :
		M_01_t64_t1 = ~|RG_zz_12 ;	// line#=../rle.cpp:61,62
	6'h0e :
		M_01_t64_t1 = ~|RG_zz_13 ;	// line#=../rle.cpp:61,62
	6'h0f :
		M_01_t64_t1 = ~|RG_zz_14 ;	// line#=../rle.cpp:61,62
	6'h10 :
		M_01_t64_t1 = ~|RG_zz_15 ;	// line#=../rle.cpp:61,62
	6'h11 :
		M_01_t64_t1 = ~|RG_zz_16 ;	// line#=../rle.cpp:61,62
	6'h12 :
		M_01_t64_t1 = ~|RG_zz_17 ;	// line#=../rle.cpp:61,62
	6'h13 :
		M_01_t64_t1 = ~|RG_zz_18 ;	// line#=../rle.cpp:61,62
	6'h14 :
		M_01_t64_t1 = ~|RG_zz_19 ;	// line#=../rle.cpp:61,62
	6'h15 :
		M_01_t64_t1 = ~|RG_zz_20 ;	// line#=../rle.cpp:61,62
	6'h16 :
		M_01_t64_t1 = ~|RG_zz_21 ;	// line#=../rle.cpp:61,62
	6'h17 :
		M_01_t64_t1 = ~|RG_zz_22 ;	// line#=../rle.cpp:61,62
	6'h18 :
		M_01_t64_t1 = ~|RG_zz_23 ;	// line#=../rle.cpp:61,62
	6'h19 :
		M_01_t64_t1 = ~|RG_zz_24 ;	// line#=../rle.cpp:61,62
	6'h1a :
		M_01_t64_t1 = ~|RG_zz_25 ;	// line#=../rle.cpp:61,62
	6'h1b :
		M_01_t64_t1 = ~|RG_zz_26 ;	// line#=../rle.cpp:61,62
	6'h1c :
		M_01_t64_t1 = ~|RG_zz_27 ;	// line#=../rle.cpp:61,62
	6'h1d :
		M_01_t64_t1 = ~|RG_zz_28 ;	// line#=../rle.cpp:61,62
	6'h1e :
		M_01_t64_t1 = ~|RG_zz_29 ;	// line#=../rle.cpp:61,62
	6'h1f :
		M_01_t64_t1 = ~|RG_zz_30 ;	// line#=../rle.cpp:61,62
	6'h20 :
		M_01_t64_t1 = ~|RG_zz_31 ;	// line#=../rle.cpp:61,62
	6'h21 :
		M_01_t64_t1 = ~|RG_zz_32 ;	// line#=../rle.cpp:61,62
	6'h22 :
		M_01_t64_t1 = ~|RG_zz_33 ;	// line#=../rle.cpp:61,62
	6'h23 :
		M_01_t64_t1 = ~|RG_zz_34 ;	// line#=../rle.cpp:61,62
	6'h24 :
		M_01_t64_t1 = ~|RG_zz_35 ;	// line#=../rle.cpp:61,62
	6'h25 :
		M_01_t64_t1 = ~|RG_zz_36 ;	// line#=../rle.cpp:61,62
	6'h26 :
		M_01_t64_t1 = ~|RG_zz_37 ;	// line#=../rle.cpp:61,62
	6'h27 :
		M_01_t64_t1 = ~|RG_zz_38 ;	// line#=../rle.cpp:61,62
	6'h28 :
		M_01_t64_t1 = ~|RG_zz_39 ;	// line#=../rle.cpp:61,62
	6'h29 :
		M_01_t64_t1 = ~|RG_zz_40 ;	// line#=../rle.cpp:61,62
	6'h2a :
		M_01_t64_t1 = ~|RG_zz_41 ;	// line#=../rle.cpp:61,62
	6'h2b :
		M_01_t64_t1 = ~|RG_zz_42 ;	// line#=../rle.cpp:61,62
	6'h2c :
		M_01_t64_t1 = ~|RG_zz_43 ;	// line#=../rle.cpp:61,62
	6'h2d :
		M_01_t64_t1 = ~|RG_zz_44 ;	// line#=../rle.cpp:61,62
	6'h2e :
		M_01_t64_t1 = ~|RG_zz_45 ;	// line#=../rle.cpp:61,62
	6'h2f :
		M_01_t64_t1 = ~|RG_zz_46 ;	// line#=../rle.cpp:61,62
	6'h30 :
		M_01_t64_t1 = ~|RG_zz_47 ;	// line#=../rle.cpp:61,62
	6'h31 :
		M_01_t64_t1 = ~|RG_zz_48 ;	// line#=../rle.cpp:61,62
	6'h32 :
		M_01_t64_t1 = ~|RG_zz_49 ;	// line#=../rle.cpp:61,62
	6'h33 :
		M_01_t64_t1 = ~|RG_zz_50 ;	// line#=../rle.cpp:61,62
	6'h34 :
		M_01_t64_t1 = ~|RG_zz_51 ;	// line#=../rle.cpp:61,62
	6'h35 :
		M_01_t64_t1 = ~|RG_zz_52 ;	// line#=../rle.cpp:61,62
	6'h36 :
		M_01_t64_t1 = ~|RG_zz_53 ;	// line#=../rle.cpp:61,62
	6'h37 :
		M_01_t64_t1 = ~|RG_zz_54 ;	// line#=../rle.cpp:61,62
	6'h38 :
		M_01_t64_t1 = ~|RG_zz_55 ;	// line#=../rle.cpp:61,62
	6'h39 :
		M_01_t64_t1 = ~|RG_zz_56 ;	// line#=../rle.cpp:61,62
	6'h3a :
		M_01_t64_t1 = ~|RG_zz_57 ;	// line#=../rle.cpp:61,62
	6'h3b :
		M_01_t64_t1 = ~|RG_zz_58 ;	// line#=../rle.cpp:61,62
	6'h3c :
		M_01_t64_t1 = ~|RG_zz_59 ;	// line#=../rle.cpp:61,62
	6'h3d :
		M_01_t64_t1 = ~|RG_zz_60 ;	// line#=../rle.cpp:61,62
	6'h3e :
		M_01_t64_t1 = ~|RG_zz_61 ;	// line#=../rle.cpp:61,62
	6'h3f :
		M_01_t64_t1 = ~|RG_zz_62 ;	// line#=../rle.cpp:61,62
	default :
		M_01_t64_t1 = 1'hx ;
	endcase
always @ ( M_01_t64_t1 or CT_35 )	// line#=../rle.cpp:61,62
	M_01_t64 = ( { 1{ CT_35 } } & M_01_t64_t1 )	// line#=../rle.cpp:61,62
		 ;	// line#=../rle.cpp:61,62
assign	JF_06 = ~M_02_t1 ;	// line#=../rle.cpp:77,78
assign	JF_06_port = JF_06 ;
assign	FL01_03_break = ( FL01_03_streg & FJ_13_14 ) ;
assign	M_219 = ( ST1_11d & FL01_01_streg ) ;
assign	FL01_01_01a = M_219 ;
assign	FL01_02_01a = U_263 ;
assign	FL01_03_01a = U_269 ;
assign	FJ_13_14 = ( U_254 & ( ~M_03_t1 ) ) ;	// line#=../rle.cpp:83,84
assign	FL01_01_eos = ( ( ST1_11d & ( ~FL01_01_streg ) ) | U_278 ) ;
assign	FL01_02_eos = ( M_215 | U_278 ) ;
assign	FL01_03_eos = ( M_216 | U_280 ) ;
always @ ( ST1_10d or U_251 or FL01_01_next or M_190 )
	begin
	FL01_01_streg_t_c1 = ( U_251 | ST1_10d ) ;
	FL01_01_streg_t = ( ( { 1{ M_190 } } & FL01_01_next )
		| ( { 1{ FL01_01_streg_t_c1 } } & 1'h1 ) ) ;
	end
assign	FL01_01_streg_en = ( U_278 | M_190 | FL01_01_streg_t_c1 ) ;
always @ ( posedge clk )
	if ( FL01_01_streg_en )
		FL01_01_streg <= FL01_01_streg_t ;
assign	M_190 = ( ST1_11d & ( ~FJ_13_14 ) ) ;
assign	M_215 = ( ( U_263 & ( ~FL01_01_ndat ) ) | ( U_262 & ( ~FL01_01_ndat ) ) ) ;
always @ ( U_262 or FL01_01_ndat or U_263 or M_215 or M_190 or ST1_10d or U_251 or 
	U_278 )
	begin
	FL01_02_streg_t_c1 = ( ( ( U_278 | U_251 ) | ST1_10d ) | ( M_190 & M_215 ) ) ;
	FL01_02_streg_t_c2 = ( M_190 & ( ( U_263 & FL01_01_ndat ) | ( U_262 & FL01_01_ndat ) ) ) ;
	FL01_02_streg_t = ( { 1{ FL01_02_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_02_streg_en = ( FL01_02_streg_t_c1 | FL01_02_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_02_streg_en )
		FL01_02_streg <= FL01_02_streg_t ;
assign	M_191 = ( ST1_11d & ( ~FL01_03_break ) ) ;
assign	M_216 = ( ( ( U_269 & FJ_13_14 ) | ( U_273 & ( ~FL01_02_ndat ) ) ) | ( U_268 & ( 
	~FL01_02_ndat ) ) ) ;
always @ ( U_268 or FL01_02_ndat or U_273 or M_216 or M_191 or ST1_10d or U_251 or 
	U_280 )
	begin
	FL01_03_streg_t_c1 = ( ( ( U_280 | U_251 ) | ST1_10d ) | ( M_191 & M_216 ) ) ;
	FL01_03_streg_t_c2 = ( M_191 & ( ( U_273 & FL01_02_ndat ) | ( U_268 & FL01_02_ndat ) ) ) ;
	FL01_03_streg_t = ( { 1{ FL01_03_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_03_streg_en = ( FL01_03_streg_t_c1 | FL01_03_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_03_streg_en )
		FL01_03_streg <= FL01_03_streg_t ;
assign	FL01_01_ndat = M_219 ;
assign	FL01_02_ndat = U_263 ;
assign	jpeg_out_a00_r_en = ST1_12d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a00_r_en )
		jpeg_out_a00_r <= rl_RD1 ;
assign	jpeg_out_a01_r_en = ST1_12d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a01_r_en )
		jpeg_out_a01_r <= rl_RD3 ;
assign	jpeg_out_a02_r_en = ST1_12d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a02_r_en )
		jpeg_out_a02_r <= rl_RD2 ;
assign	jpeg_out_a03_r_en = ST1_13d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a03_r_en )
		jpeg_out_a03_r <= rl_RD3 ;
assign	jpeg_out_a04_r_en = ST1_13d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a04_r_en )
		jpeg_out_a04_r <= rl_RD2 ;
assign	jpeg_out_a05_r_en = ST1_13d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a05_r_en )
		jpeg_out_a05_r <= rl_RD1 ;
assign	jpeg_out_a06_r_en = ST1_14d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a06_r_en )
		jpeg_out_a06_r <= rl_RD3 ;
assign	jpeg_out_a07_r_en = ST1_14d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a07_r_en )
		jpeg_out_a07_r <= rl_RD2 ;
assign	jpeg_out_a08_r_en = ST1_14d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a08_r_en )
		jpeg_out_a08_r <= rl_RD1 ;
assign	jpeg_out_a09_r_en = ST1_15d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a09_r_en )
		jpeg_out_a09_r <= rl_RD3 ;
assign	jpeg_out_a10_r_en = ST1_15d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a10_r_en )
		jpeg_out_a10_r <= rl_RD2 ;
assign	jpeg_out_a11_r_en = ST1_15d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a11_r_en )
		jpeg_out_a11_r <= rl_RD1 ;
assign	jpeg_out_a12_r_en = ST1_16d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a12_r_en )
		jpeg_out_a12_r <= rl_RD3 ;
assign	jpeg_out_a13_r_en = ST1_16d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a13_r_en )
		jpeg_out_a13_r <= rl_RD2 ;
assign	jpeg_out_a14_r_en = ST1_16d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a14_r_en )
		jpeg_out_a14_r <= rl_RD1 ;
assign	jpeg_out_a15_r_en = ST1_17d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a15_r_en )
		jpeg_out_a15_r <= rl_RD3 ;
assign	jpeg_out_a16_r_en = ST1_17d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a16_r_en )
		jpeg_out_a16_r <= rl_RD2 ;
assign	jpeg_out_a17_r_en = ST1_17d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a17_r_en )
		jpeg_out_a17_r <= rl_RD1 ;
assign	jpeg_out_a18_r_en = ST1_18d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a18_r_en )
		jpeg_out_a18_r <= rl_RD3 ;
assign	jpeg_out_a19_r_en = ST1_18d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a19_r_en )
		jpeg_out_a19_r <= rl_RD2 ;
assign	jpeg_out_a20_r_en = ST1_18d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a20_r_en )
		jpeg_out_a20_r <= rl_RD1 ;
assign	jpeg_out_a21_r_en = ST1_19d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a21_r_en )
		jpeg_out_a21_r <= rl_RD3 ;
assign	jpeg_out_a22_r_en = ST1_19d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a22_r_en )
		jpeg_out_a22_r <= rl_RD2 ;
assign	jpeg_out_a23_r_en = ST1_19d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a23_r_en )
		jpeg_out_a23_r <= rl_RD1 ;
assign	jpeg_out_a24_r_en = ST1_20d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a24_r_en )
		jpeg_out_a24_r <= rl_RD3 ;
assign	jpeg_out_a25_r_en = ST1_20d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a25_r_en )
		jpeg_out_a25_r <= rl_RD2 ;
assign	jpeg_out_a26_r_en = ST1_20d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a26_r_en )
		jpeg_out_a26_r <= rl_RD1 ;
assign	jpeg_out_a27_r_en = ST1_21d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a27_r_en )
		jpeg_out_a27_r <= rl_RD3 ;
assign	jpeg_out_a28_r_en = ST1_21d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a28_r_en )
		jpeg_out_a28_r <= rl_RD2 ;
assign	jpeg_out_a29_r_en = ST1_21d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a29_r_en )
		jpeg_out_a29_r <= rl_RD1 ;
assign	jpeg_out_a30_r_en = ST1_22d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a30_r_en )
		jpeg_out_a30_r <= rl_RD3 ;
assign	jpeg_out_a31_r_en = ST1_22d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a31_r_en )
		jpeg_out_a31_r <= rl_RD2 ;
assign	jpeg_out_a32_r_en = ST1_22d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a32_r_en )
		jpeg_out_a32_r <= rl_RD1 ;
assign	jpeg_out_a33_r_en = ST1_23d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a33_r_en )
		jpeg_out_a33_r <= rl_RD3 ;
assign	jpeg_out_a34_r_en = ST1_23d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a34_r_en )
		jpeg_out_a34_r <= rl_RD2 ;
assign	jpeg_out_a35_r_en = ST1_23d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a35_r_en )
		jpeg_out_a35_r <= rl_RD1 ;
assign	jpeg_out_a36_r_en = ST1_24d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a36_r_en )
		jpeg_out_a36_r <= rl_RD3 ;
assign	jpeg_out_a37_r_en = ST1_24d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a37_r_en )
		jpeg_out_a37_r <= rl_RD2 ;
assign	jpeg_out_a38_r_en = ST1_24d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a38_r_en )
		jpeg_out_a38_r <= rl_RD1 ;
assign	jpeg_out_a39_r_en = ST1_25d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a39_r_en )
		jpeg_out_a39_r <= rl_RD3 ;
assign	jpeg_out_a40_r_en = ST1_25d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a40_r_en )
		jpeg_out_a40_r <= rl_RD2 ;
assign	jpeg_out_a41_r_en = ST1_25d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a41_r_en )
		jpeg_out_a41_r <= rl_RD1 ;
assign	jpeg_out_a42_r_en = ST1_26d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a42_r_en )
		jpeg_out_a42_r <= rl_RD3 ;
assign	jpeg_out_a43_r_en = ST1_26d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a43_r_en )
		jpeg_out_a43_r <= rl_RD2 ;
assign	jpeg_out_a44_r_en = ST1_26d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a44_r_en )
		jpeg_out_a44_r <= rl_RD1 ;
assign	jpeg_out_a45_r_en = ST1_27d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a45_r_en )
		jpeg_out_a45_r <= rl_RD3 ;
assign	jpeg_out_a46_r_en = ST1_27d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a46_r_en )
		jpeg_out_a46_r <= rl_RD2 ;
assign	jpeg_out_a47_r_en = ST1_27d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a47_r_en )
		jpeg_out_a47_r <= rl_RD1 ;
assign	jpeg_out_a48_r_en = ST1_28d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a48_r_en )
		jpeg_out_a48_r <= rl_RD3 ;
assign	jpeg_out_a49_r_en = ST1_28d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a49_r_en )
		jpeg_out_a49_r <= rl_RD2 ;
assign	jpeg_out_a50_r_en = ST1_28d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a50_r_en )
		jpeg_out_a50_r <= rl_RD1 ;
assign	jpeg_out_a51_r_en = ST1_29d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a51_r_en )
		jpeg_out_a51_r <= rl_RD3 ;
assign	jpeg_out_a52_r_en = ST1_29d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a52_r_en )
		jpeg_out_a52_r <= rl_RD2 ;
assign	jpeg_out_a53_r_en = ST1_29d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a53_r_en )
		jpeg_out_a53_r <= rl_RD1 ;
assign	jpeg_out_a54_r_en = ST1_30d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a54_r_en )
		jpeg_out_a54_r <= rl_RD3 ;
assign	jpeg_out_a55_r_en = ST1_30d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a55_r_en )
		jpeg_out_a55_r <= rl_RD2 ;
assign	jpeg_out_a56_r_en = ST1_30d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a56_r_en )
		jpeg_out_a56_r <= rl_RD1 ;
assign	jpeg_out_a57_r_en = ST1_31d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a57_r_en )
		jpeg_out_a57_r <= rl_RD3 ;
assign	jpeg_out_a58_r_en = ST1_31d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a58_r_en )
		jpeg_out_a58_r <= rl_RD2 ;
assign	jpeg_out_a59_r_en = ST1_31d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a59_r_en )
		jpeg_out_a59_r <= rl_RD1 ;
assign	jpeg_out_a60_r_en = ST1_32d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a60_r_en )
		jpeg_out_a60_r <= rl_RD3 ;
assign	jpeg_out_a61_r_en = ST1_32d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a61_r_en )
		jpeg_out_a61_r <= rl_RD2 ;
assign	jpeg_out_a62_r_en = ST1_32d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a62_r_en )
		jpeg_out_a62_r <= rl_RD1 ;
assign	jpeg_out_a63_r_en = ST1_33d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a63_r_en )
		jpeg_out_a63_r <= rl_RD2 ;
assign	jpeg_out_a64_r_en = ST1_33d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a64_r_en )
		jpeg_out_a64_r <= rl_RD3 ;
assign	jpeg_out_a65_r_en = ST1_33d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a65_r_en )
		jpeg_out_a65_r <= rl_RD1 ;
assign	jpeg_out_a66_r_en = ST1_34d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a66_r_en )
		jpeg_out_a66_r <= rl_RD2 ;
assign	jpeg_out_a67_r_en = ST1_34d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a67_r_en )
		jpeg_out_a67_r <= rl_RD3 ;
assign	jpeg_out_a68_r_en = ST1_34d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a68_r_en )
		jpeg_out_a68_r <= rl_RD1 ;
assign	jpeg_out_a69_r_en = ST1_35d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a69_r_en )
		jpeg_out_a69_r <= rl_RD2 ;
assign	jpeg_out_a70_r_en = ST1_35d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a70_r_en )
		jpeg_out_a70_r <= rl_RD3 ;
assign	jpeg_out_a71_r_en = ST1_35d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a71_r_en )
		jpeg_out_a71_r <= rl_RD1 ;
assign	jpeg_out_a72_r_en = ST1_36d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a72_r_en )
		jpeg_out_a72_r <= rl_RD2 ;
assign	jpeg_out_a73_r_en = ST1_36d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a73_r_en )
		jpeg_out_a73_r <= rl_RD3 ;
assign	jpeg_out_a74_r_en = ST1_36d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a74_r_en )
		jpeg_out_a74_r <= rl_RD1 ;
assign	jpeg_out_a75_r_en = ST1_37d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a75_r_en )
		jpeg_out_a75_r <= rl_RD2 ;
assign	jpeg_out_a76_r_en = ST1_37d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a76_r_en )
		jpeg_out_a76_r <= rl_RD3 ;
assign	jpeg_out_a77_r_en = ST1_37d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a77_r_en )
		jpeg_out_a77_r <= rl_RD1 ;
assign	jpeg_out_a78_r_en = ST1_38d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a78_r_en )
		jpeg_out_a78_r <= rl_RD2 ;
assign	jpeg_out_a79_r_en = ST1_38d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a79_r_en )
		jpeg_out_a79_r <= rl_RD3 ;
assign	jpeg_out_a80_r_en = ST1_38d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a80_r_en )
		jpeg_out_a80_r <= rl_RD1 ;
assign	jpeg_out_a81_r_en = ST1_39d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a81_r_en )
		jpeg_out_a81_r <= rl_RD2 ;
assign	jpeg_out_a82_r_en = ST1_39d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a82_r_en )
		jpeg_out_a82_r <= rl_RD3 ;
assign	jpeg_out_a83_r_en = ST1_39d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a83_r_en )
		jpeg_out_a83_r <= rl_RD1 ;
assign	jpeg_out_a84_r_en = ST1_40d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a84_r_en )
		jpeg_out_a84_r <= rl_RD2 ;
assign	jpeg_out_a85_r_en = ST1_40d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a85_r_en )
		jpeg_out_a85_r <= rl_RD3 ;
assign	jpeg_out_a86_r_en = ST1_40d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a86_r_en )
		jpeg_out_a86_r <= rl_RD1 ;
assign	jpeg_out_a87_r_en = ST1_41d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a87_r_en )
		jpeg_out_a87_r <= rl_RD2 ;
assign	jpeg_out_a88_r_en = ST1_41d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a88_r_en )
		jpeg_out_a88_r <= rl_RD3 ;
assign	jpeg_out_a89_r_en = ST1_41d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a89_r_en )
		jpeg_out_a89_r <= rl_RD1 ;
assign	jpeg_out_a90_r_en = ST1_42d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a90_r_en )
		jpeg_out_a90_r <= rl_RD2 ;
assign	jpeg_out_a91_r_en = ST1_42d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a91_r_en )
		jpeg_out_a91_r <= rl_RD3 ;
assign	jpeg_out_a92_r_en = ST1_42d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a92_r_en )
		jpeg_out_a92_r <= rl_RD1 ;
assign	jpeg_out_a93_r_en = ST1_43d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a93_r_en )
		jpeg_out_a93_r <= rl_RD2 ;
assign	jpeg_out_a94_r_en = ST1_43d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a94_r_en )
		jpeg_out_a94_r <= rl_RD3 ;
assign	jpeg_out_a95_r_en = ST1_43d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a95_r_en )
		jpeg_out_a95_r <= rl_RD1 ;
assign	jpeg_out_a96_r_en = ST1_44d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a96_r_en )
		jpeg_out_a96_r <= rl_RD2 ;
assign	jpeg_out_a97_r_en = ST1_44d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a97_r_en )
		jpeg_out_a97_r <= rl_RD3 ;
assign	jpeg_out_a98_r_en = ST1_44d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a98_r_en )
		jpeg_out_a98_r <= rl_RD1 ;
assign	jpeg_out_a99_r_en = ST1_45d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a99_r_en )
		jpeg_out_a99_r <= rl_RD2 ;
assign	jpeg_out_a100_r_en = ST1_45d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a100_r_en )
		jpeg_out_a100_r <= rl_RD3 ;
assign	jpeg_out_a101_r_en = ST1_45d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a101_r_en )
		jpeg_out_a101_r <= rl_RD1 ;
assign	jpeg_out_a102_r_en = ST1_46d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a102_r_en )
		jpeg_out_a102_r <= rl_RD2 ;
assign	jpeg_out_a103_r_en = ST1_46d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a103_r_en )
		jpeg_out_a103_r <= rl_RD3 ;
assign	jpeg_out_a104_r_en = ST1_46d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a104_r_en )
		jpeg_out_a104_r <= rl_RD1 ;
assign	jpeg_out_a105_r_en = ST1_47d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a105_r_en )
		jpeg_out_a105_r <= rl_RD2 ;
assign	jpeg_out_a106_r_en = ST1_47d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a106_r_en )
		jpeg_out_a106_r <= rl_RD3 ;
assign	jpeg_out_a107_r_en = ST1_47d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a107_r_en )
		jpeg_out_a107_r <= rl_RD1 ;
assign	jpeg_out_a108_r_en = ST1_48d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a108_r_en )
		jpeg_out_a108_r <= rl_RD2 ;
assign	jpeg_out_a109_r_en = ST1_48d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a109_r_en )
		jpeg_out_a109_r <= rl_RD3 ;
assign	jpeg_out_a110_r_en = ST1_48d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a110_r_en )
		jpeg_out_a110_r <= rl_RD1 ;
assign	jpeg_out_a111_r_en = ST1_49d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a111_r_en )
		jpeg_out_a111_r <= rl_RD2 ;
assign	jpeg_out_a112_r_en = ST1_49d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a112_r_en )
		jpeg_out_a112_r <= rl_RD3 ;
assign	jpeg_out_a113_r_en = ST1_49d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a113_r_en )
		jpeg_out_a113_r <= rl_RD1 ;
assign	jpeg_out_a114_r_en = ST1_50d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a114_r_en )
		jpeg_out_a114_r <= rl_RD2 ;
assign	jpeg_out_a115_r_en = ST1_50d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a115_r_en )
		jpeg_out_a115_r <= rl_RD3 ;
assign	jpeg_out_a116_r_en = ST1_50d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a116_r_en )
		jpeg_out_a116_r <= rl_RD1 ;
assign	jpeg_out_a117_r_en = ST1_51d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a117_r_en )
		jpeg_out_a117_r <= rl_RD2 ;
assign	jpeg_out_a118_r_en = ST1_51d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a118_r_en )
		jpeg_out_a118_r <= rl_RD3 ;
assign	jpeg_out_a119_r_en = ST1_51d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a119_r_en )
		jpeg_out_a119_r <= rl_RD1 ;
assign	jpeg_out_a120_r_en = ST1_52d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a120_r_en )
		jpeg_out_a120_r <= rl_RD2 ;
assign	jpeg_out_a121_r_en = ST1_52d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a121_r_en )
		jpeg_out_a121_r <= rl_RD3 ;
assign	jpeg_out_a122_r_en = ST1_52d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a122_r_en )
		jpeg_out_a122_r <= rl_RD1 ;
assign	jpeg_out_a123_r_en = ST1_53d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a123_r_en )
		jpeg_out_a123_r <= rl_RD2 ;
assign	jpeg_out_a124_r_en = ST1_53d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a124_r_en )
		jpeg_out_a124_r <= rl_RD3 ;
assign	jpeg_out_a125_r_en = ST1_53d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a125_r_en )
		jpeg_out_a125_r <= rl_RD1 ;
assign	jpeg_out_a126_r_en = ST1_54d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a126_r_en )
		jpeg_out_a126_r <= rl_RD1 ;
assign	jpeg_out_a127_r_en = ST1_54d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a127_r_en )
		jpeg_out_a127_r <= rl_RD2 ;
assign	jpeg_len_out_r_en = ST1_12d ;
always @ ( posedge clk )	// line#=../rle.cpp:93
	if ( jpeg_len_out_r_en )
		jpeg_len_out_r <= { 4'h0 , RG_len_03 } ;
always @ ( ST1_54d )
	valid_r_t = ( { 1{ ST1_54d } } & 1'h1 )	// line#=../rle.cpp:95
		 ;	// line#=../rle.cpp:30
assign	valid_r_en = ( ST1_01d | ST1_54d ) ;
always @ ( posedge clk )
	if ( valid_r_en )
		valid_r <= valid_r_t ;	// line#=../rle.cpp:30,95
assign	incr8u1i1 = RG_len_01_1 ;	// line#=../rle.cpp:68,73,79
always @ ( RG_k_01 or U_87 or RG_k or U_05 )
	TR_03 = ( ( { 6{ U_05 } } & RG_k )		// line#=../rle.cpp:111
		| ( { 6{ U_87 } } & RG_k_01 [5:0] )	// line#=../rle.cpp:142
		) ;
always @ ( TR_03 or U_87 or U_05 or incr8u1ot or M_189 )
	begin
	incr8u2i1_c1 = ( U_05 | U_87 ) ;	// line#=../rle.cpp:111,142
	incr8u2i1 = ( ( { 8{ M_189 } } & incr8u1ot )		// line#=../rle.cpp:68,69,73,74,79,80
		| ( { 8{ incr8u2i1_c1 } } & { 2'h0 , TR_03 } )	// line#=../rle.cpp:111,142
		) ;
	end
assign	incr32s1i1 = RG_j_k ;	// line#=../rle.cpp:64,114,125,145,156
assign	incr32s2i1 = RG_i ;	// line#=../rle.cpp:63,74,119,129,150,160
assign	decr32s1i1 = RG_i ;	// line#=../rle.cpp:124,155
assign	decr32s2i1 = RG_j_k ;	// line#=../rle.cpp:130,161
always @ ( incr8u2ot or CT_35 or ST1_07d or RG_len_01_1 or U_252 )	// line#=../rle.cpp:57,58
	begin
	sub8u_7_11i1_c1 = ( ST1_07d & ( ~CT_35 ) ) ;	// line#=../rle.cpp:69,74,77,78
	sub8u_7_11i1 = ( ( { 7{ U_252 } } & RG_len_01_1 [6:0] )		// line#=../rle.cpp:83,84
		| ( { 7{ sub8u_7_11i1_c1 } } & incr8u2ot [6:0] )	// line#=../rle.cpp:69,74,77,78
		) ;
	end
assign	sub8u_7_11i2 = { 1'h1 , U_252 } ;	// line#=../rle.cpp:77,78,83,84
assign	M_193 = ( U_88 | ST1_12d ) ;
always @ ( ST1_13d )
	M_220 = ( { 2{ ST1_13d } } & 2'h3 )
		 ;	// line#=../rle.cpp:52
always @ ( ST1_15d )
	TR_17 = ( { 2{ ST1_15d } } & 2'h3 )
		 ;
assign	M_197 = ( ST1_14d | ST1_15d ) ;
always @ ( ST1_16d or TR_17 or M_197 )
	TR_18 = ( ( { 3{ M_197 } } & { 1'h0 , TR_17 } )
		| ( { 3{ ST1_16d } } & 3'h6 ) ) ;
assign	M_194 = ( M_193 | ST1_13d ) ;
always @ ( TR_18 or ST1_16d or M_197 or M_220 or M_194 )
	begin
	TR_05_c1 = ( M_197 | ST1_16d ) ;
	TR_05 = ( ( { 4{ M_194 } } & { 1'h0 , M_220 [1] , 1'h0 , M_220 [0] } )	// line#=../rle.cpp:52
		| ( { 4{ TR_05_c1 } } & { 1'h1 , TR_18 } ) ) ;
	end
always @ ( ST1_19d or ST1_18d or ST1_17d )
	TR_19 = ( ( { 3{ ST1_17d } } & 3'h1 )
		| ( { 3{ ST1_18d } } & 3'h4 )
		| ( { 3{ ST1_19d } } & 3'h7 ) ) ;
always @ ( ST1_21d or ST1_20d )
	TR_32 = ( ( { 3{ ST1_20d } } & 3'h2 )
		| ( { 3{ ST1_21d } } & 3'h5 ) ) ;
assign	M_199 = ( ( ST1_17d | ST1_18d ) | ST1_19d ) ;
always @ ( TR_32 or ST1_21d or ST1_20d or TR_19 or M_199 )
	begin
	TR_20_c1 = ( ST1_20d | ST1_21d ) ;
	TR_20 = ( ( { 4{ M_199 } } & { 1'h0 , TR_19 } )
		| ( { 4{ TR_20_c1 } } & { 1'h1 , TR_32 } ) ) ;
	end
assign	M_196 = ( ( ( M_194 | ST1_14d ) | ST1_15d ) | ST1_16d ) ;
always @ ( TR_20 or ST1_21d or ST1_20d or M_199 or TR_05 or M_196 )
	begin
	TR_06_c1 = ( ( M_199 | ST1_20d ) | ST1_21d ) ;
	TR_06 = ( ( { 5{ M_196 } } & { 1'h0 , TR_05 } )	// line#=../rle.cpp:52
		| ( { 5{ TR_06_c1 } } & { 1'h1 , TR_20 } ) ) ;
	end
always @ ( ST1_23d )
	TR_21 = ( { 2{ ST1_23d } } & 2'h3 )
		 ;
assign	M_200 = ( ST1_22d | ST1_23d ) ;
always @ ( ST1_24d or TR_21 or M_200 )
	TR_22 = ( ( { 3{ M_200 } } & { 1'h0 , TR_21 } )
		| ( { 3{ ST1_24d } } & 3'h6 ) ) ;
always @ ( ST1_27d or ST1_26d or ST1_25d )
	TR_33 = ( ( { 3{ ST1_25d } } & 3'h1 )
		| ( { 3{ ST1_26d } } & 3'h4 )
		| ( { 3{ ST1_27d } } & 3'h7 ) ) ;
assign	M_201 = ( M_200 | ST1_24d ) ;
always @ ( TR_33 or ST1_27d or ST1_26d or ST1_25d or TR_22 or M_201 )
	begin
	TR_23_c1 = ( ( ST1_25d | ST1_26d ) | ST1_27d ) ;
	TR_23 = ( ( { 4{ M_201 } } & { 1'h0 , TR_22 } )
		| ( { 4{ TR_23_c1 } } & { 1'h1 , TR_33 } ) ) ;
	end
always @ ( ST1_29d or ST1_28d )
	TR_34 = ( ( { 3{ ST1_28d } } & 3'h2 )
		| ( { 3{ ST1_29d } } & 3'h5 ) ) ;
always @ ( ST1_31d )
	TR_41 = ( { 2{ ST1_31d } } & 2'h3 )
		 ;
assign	M_204 = ( ST1_30d | ST1_31d ) ;
always @ ( ST1_32d or TR_41 or M_204 )
	TR_42 = ( ( { 3{ M_204 } } & { 1'h0 , TR_41 } )
		| ( { 3{ ST1_32d } } & 3'h6 ) ) ;
assign	M_203 = ( ST1_28d | ST1_29d ) ;
always @ ( TR_42 or ST1_32d or M_204 or TR_34 or M_203 )
	begin
	TR_35_c1 = ( M_204 | ST1_32d ) ;
	TR_35 = ( ( { 4{ M_203 } } & { 1'h0 , TR_34 } )
		| ( { 4{ TR_35_c1 } } & { 1'h1 , TR_42 } ) ) ;
	end
assign	M_202 = ( ( ( M_201 | ST1_25d ) | ST1_26d ) | ST1_27d ) ;
always @ ( TR_35 or ST1_32d or ST1_31d or ST1_30d or M_203 or TR_23 or M_202 )
	begin
	TR_24_c1 = ( ( ( M_203 | ST1_30d ) | ST1_31d ) | ST1_32d ) ;
	TR_24 = ( ( { 5{ M_202 } } & { 1'h0 , TR_23 } )
		| ( { 5{ TR_24_c1 } } & { 1'h1 , TR_35 } ) ) ;
	end
assign	M_198 = ( ( ( ( ( M_196 | ST1_17d ) | ST1_18d ) | ST1_19d ) | ST1_20d ) | 
	ST1_21d ) ;
always @ ( TR_24 or ST1_32d or ST1_31d or ST1_30d or ST1_29d or ST1_28d or M_202 or 
	TR_06 or M_198 )
	begin
	TR_07_c1 = ( ( ( ( ( M_202 | ST1_28d ) | ST1_29d ) | ST1_30d ) | ST1_31d ) | 
		ST1_32d ) ;
	TR_07 = ( ( { 6{ M_198 } } & { 1'h0 , TR_06 } )	// line#=../rle.cpp:52
		| ( { 6{ TR_07_c1 } } & { 1'h1 , TR_24 } ) ) ;
	end
always @ ( ST1_35d or ST1_34d or ST1_33d )
	TR_08 = ( ( { 3{ ST1_33d } } & 3'h1 )
		| ( { 3{ ST1_34d } } & 3'h4 )
		| ( { 3{ ST1_35d } } & 3'h7 ) ) ;
always @ ( ST1_37d or ST1_36d )
	TR_25 = ( ( { 3{ ST1_36d } } & 3'h2 )
		| ( { 3{ ST1_37d } } & 3'h5 ) ) ;
assign	M_205 = ( ( ST1_33d | ST1_34d ) | ST1_35d ) ;
always @ ( TR_25 or ST1_37d or ST1_36d or TR_08 or M_205 )
	begin
	TR_09_c1 = ( ST1_36d | ST1_37d ) ;
	TR_09 = ( ( { 4{ M_205 } } & { 1'h0 , TR_08 } )
		| ( { 4{ TR_09_c1 } } & { 1'h1 , TR_25 } ) ) ;
	end
always @ ( ST1_39d )
	TR_26 = ( { 2{ ST1_39d } } & 2'h3 )
		 ;
assign	M_208 = ( ST1_38d | ST1_39d ) ;
always @ ( ST1_40d or TR_26 or M_208 )
	TR_27 = ( ( { 3{ M_208 } } & { 1'h0 , TR_26 } )
		| ( { 3{ ST1_40d } } & 3'h6 ) ) ;
always @ ( ST1_43d or ST1_42d or ST1_41d )
	TR_36 = ( ( { 3{ ST1_41d } } & 3'h1 )
		| ( { 3{ ST1_42d } } & 3'h4 )
		| ( { 3{ ST1_43d } } & 3'h7 ) ) ;
assign	M_209 = ( M_208 | ST1_40d ) ;
always @ ( TR_36 or ST1_43d or ST1_42d or ST1_41d or TR_27 or M_209 )
	begin
	TR_28_c1 = ( ( ST1_41d | ST1_42d ) | ST1_43d ) ;
	TR_28 = ( ( { 4{ M_209 } } & { 1'h0 , TR_27 } )
		| ( { 4{ TR_28_c1 } } & { 1'h1 , TR_36 } ) ) ;
	end
assign	M_206 = ( ( M_205 | ST1_36d ) | ST1_37d ) ;
always @ ( TR_28 or ST1_43d or ST1_42d or ST1_41d or M_209 or TR_09 or M_206 )
	begin
	TR_10_c1 = ( ( ( M_209 | ST1_41d ) | ST1_42d ) | ST1_43d ) ;
	TR_10 = ( ( { 5{ M_206 } } & { 1'h0 , TR_09 } )
		| ( { 5{ TR_10_c1 } } & { 1'h1 , TR_28 } ) ) ;
	end
always @ ( ST1_45d or ST1_44d )
	TR_29 = ( ( { 3{ ST1_44d } } & 3'h2 )
		| ( { 3{ ST1_45d } } & 3'h5 ) ) ;
always @ ( ST1_47d )
	TR_37 = ( { 2{ ST1_47d } } & 2'h3 )
		 ;
assign	M_212 = ( ST1_46d | ST1_47d ) ;
always @ ( ST1_48d or TR_37 or M_212 )
	TR_38 = ( ( { 3{ M_212 } } & { 1'h0 , TR_37 } )
		| ( { 3{ ST1_48d } } & 3'h6 ) ) ;
assign	M_210 = ( ST1_44d | ST1_45d ) ;
always @ ( TR_38 or ST1_48d or M_212 or TR_29 or M_210 )
	begin
	TR_30_c1 = ( M_212 | ST1_48d ) ;
	TR_30 = ( ( { 4{ M_210 } } & { 1'h0 , TR_29 } )
		| ( { 4{ TR_30_c1 } } & { 1'h1 , TR_38 } ) ) ;
	end
always @ ( ST1_51d or ST1_50d or ST1_49d )
	TR_39 = ( ( { 3{ ST1_49d } } & 3'h1 )
		| ( { 3{ ST1_50d } } & 3'h4 )
		| ( { 3{ ST1_51d } } & 3'h7 ) ) ;
always @ ( ST1_54d or ST1_53d or ST1_52d )
	TR_43 = ( ( { 3{ ST1_52d } } & 3'h2 )
		| ( { 3{ ST1_53d } } & 3'h5 )
		| ( { 3{ ST1_54d } } & 3'h6 ) ) ;
assign	M_213 = ( ( ST1_49d | ST1_50d ) | ST1_51d ) ;
always @ ( TR_43 or ST1_54d or ST1_53d or ST1_52d or TR_39 or M_213 )
	begin
	TR_40_c1 = ( ( ST1_52d | ST1_53d ) | ST1_54d ) ;
	TR_40 = ( ( { 4{ M_213 } } & { 1'h0 , TR_39 } )
		| ( { 4{ TR_40_c1 } } & { 1'h1 , TR_43 } ) ) ;
	end
assign	M_211 = ( ( ( M_210 | ST1_46d ) | ST1_47d ) | ST1_48d ) ;
always @ ( TR_40 or ST1_54d or ST1_53d or ST1_52d or M_213 or TR_30 or M_211 )
	begin
	TR_31_c1 = ( ( ( M_213 | ST1_52d ) | ST1_53d ) | ST1_54d ) ;
	TR_31 = ( ( { 5{ M_211 } } & { 1'h0 , TR_30 } )
		| ( { 5{ TR_31_c1 } } & { 1'h1 , TR_40 } ) ) ;
	end
assign	M_207 = ( ( ( ( ( ( M_206 | ST1_38d ) | ST1_39d ) | ST1_40d ) | ST1_41d ) | 
	ST1_42d ) | ST1_43d ) ;
always @ ( TR_31 or ST1_54d or ST1_53d or ST1_52d or ST1_51d or ST1_50d or ST1_49d or 
	M_211 or TR_10 or M_207 )
	begin
	TR_11_c1 = ( ( ( ( ( ( M_211 | ST1_49d ) | ST1_50d ) | ST1_51d ) | ST1_52d ) | 
		ST1_53d ) | ST1_54d ) ;
	TR_11 = ( ( { 6{ M_207 } } & { 1'h0 , TR_10 } )
		| ( { 6{ TR_11_c1 } } & { 1'h1 , TR_31 } ) ) ;
	end
assign	M_189 = ( ST1_07d | ST1_10d ) ;
always @ ( TR_11 or ST1_54d or ST1_53d or ST1_52d or ST1_51d or ST1_50d or ST1_49d or 
	ST1_48d or ST1_47d or ST1_46d or ST1_45d or ST1_44d or M_207 or RG_140_02 or 
	U_257 or incr8u1ot or M_189 or RG_len_01_1 or U_248 or U_175 or TR_07 or 
	ST1_32d or ST1_31d or ST1_30d or ST1_29d or ST1_28d or ST1_27d or ST1_26d or 
	ST1_25d or ST1_24d or ST1_23d or ST1_22d or M_198 )
	begin
	rl_AD1_c1 = ( ( ( ( ( ( ( ( ( ( ( M_198 | ST1_22d ) | ST1_23d ) | ST1_24d ) | 
		ST1_25d ) | ST1_26d ) | ST1_27d ) | ST1_28d ) | ST1_29d ) | ST1_30d ) | 
		ST1_31d ) | ST1_32d ) ;	// line#=../rle.cpp:52
	rl_AD1_c2 = ( U_175 | U_248 ) ;	// line#=../rle.cpp:68,73,79
	rl_AD1_c3 = ( ( ( ( ( ( ( ( ( ( ( M_207 | ST1_44d ) | ST1_45d ) | ST1_46d ) | 
		ST1_47d ) | ST1_48d ) | ST1_49d ) | ST1_50d ) | ST1_51d ) | ST1_52d ) | 
		ST1_53d ) | ST1_54d ) ;
	rl_AD1 = ( ( { 7{ rl_AD1_c1 } } & { 1'h0 , TR_07 } )	// line#=../rle.cpp:52
		| ( { 7{ rl_AD1_c2 } } & RG_len_01_1 [6:0] )	// line#=../rle.cpp:68,73,79
		| ( { 7{ M_189 } } & incr8u1ot [6:0] )		// line#=../rle.cpp:68,69,73,74,79,80
		| ( { 7{ U_257 } } & RG_140_02 )		// line#=../rle.cpp:85
		| ( { 7{ rl_AD1_c3 } } & { 1'h1 , TR_11 } ) ) ;
	end
always @ ( RG_zz_62 or RG_zz_61 or RG_zz_60 or RG_zz_59 or RG_zz_58 or RG_zz_57 or 
	RG_zz_56 or RG_zz_55 or RG_zz_54 or RG_zz_53 or RG_zz_52 or RG_zz_51 or 
	RG_zz_50 or RG_zz_49 or RG_zz_48 or RG_zz_47 or RG_zz_46 or RG_zz_45 or 
	RG_zz_44 or RG_zz_43 or RG_zz_42 or RG_zz_41 or RG_zz_40 or RG_zz_39 or 
	RG_zz_38 or RG_zz_37 or RG_zz_36 or RG_zz_35 or RG_zz_34 or RG_zz_33 or 
	RG_zz_32 or RG_zz_31 or RG_zz_30 or RG_zz_29 or RG_zz_28 or RG_zz_27 or 
	RG_zz_26 or RG_zz_25 or RG_zz_24 or RG_zz_23 or RG_zz_22 or RG_zz_21 or 
	RG_zz_20 or RG_zz_19 or RG_zz_18 or RG_zz_17 or RG_zz_16 or RG_zz_15 or 
	RG_zz_14 or RG_zz_13 or RG_zz_12 or RG_zz_11 or RG_zz_10 or RG_zz_9 or RG_zz_8 or 
	RG_zz_7 or RG_zz_6 or RG_zz_5 or RG_zz_4 or RG_zz_3 or RG_zz_2 or RG_zz_1 or 
	RG_zz or RG_quantized_block_zz or RG_k )	// line#=../rle.cpp:74
	case ( RG_k )
	6'h00 :
		rl_WD1_t1 = RG_quantized_block_zz ;	// line#=../rle.cpp:74
	6'h01 :
		rl_WD1_t1 = RG_zz ;	// line#=../rle.cpp:74
	6'h02 :
		rl_WD1_t1 = RG_zz_1 ;	// line#=../rle.cpp:74
	6'h03 :
		rl_WD1_t1 = RG_zz_2 ;	// line#=../rle.cpp:74
	6'h04 :
		rl_WD1_t1 = RG_zz_3 ;	// line#=../rle.cpp:74
	6'h05 :
		rl_WD1_t1 = RG_zz_4 ;	// line#=../rle.cpp:74
	6'h06 :
		rl_WD1_t1 = RG_zz_5 ;	// line#=../rle.cpp:74
	6'h07 :
		rl_WD1_t1 = RG_zz_6 ;	// line#=../rle.cpp:74
	6'h08 :
		rl_WD1_t1 = RG_zz_7 ;	// line#=../rle.cpp:74
	6'h09 :
		rl_WD1_t1 = RG_zz_8 ;	// line#=../rle.cpp:74
	6'h0a :
		rl_WD1_t1 = RG_zz_9 ;	// line#=../rle.cpp:74
	6'h0b :
		rl_WD1_t1 = RG_zz_10 ;	// line#=../rle.cpp:74
	6'h0c :
		rl_WD1_t1 = RG_zz_11 ;	// line#=../rle.cpp:74
	6'h0d :
		rl_WD1_t1 = RG_zz_12 ;	// line#=../rle.cpp:74
	6'h0e :
		rl_WD1_t1 = RG_zz_13 ;	// line#=../rle.cpp:74
	6'h0f :
		rl_WD1_t1 = RG_zz_14 ;	// line#=../rle.cpp:74
	6'h10 :
		rl_WD1_t1 = RG_zz_15 ;	// line#=../rle.cpp:74
	6'h11 :
		rl_WD1_t1 = RG_zz_16 ;	// line#=../rle.cpp:74
	6'h12 :
		rl_WD1_t1 = RG_zz_17 ;	// line#=../rle.cpp:74
	6'h13 :
		rl_WD1_t1 = RG_zz_18 ;	// line#=../rle.cpp:74
	6'h14 :
		rl_WD1_t1 = RG_zz_19 ;	// line#=../rle.cpp:74
	6'h15 :
		rl_WD1_t1 = RG_zz_20 ;	// line#=../rle.cpp:74
	6'h16 :
		rl_WD1_t1 = RG_zz_21 ;	// line#=../rle.cpp:74
	6'h17 :
		rl_WD1_t1 = RG_zz_22 ;	// line#=../rle.cpp:74
	6'h18 :
		rl_WD1_t1 = RG_zz_23 ;	// line#=../rle.cpp:74
	6'h19 :
		rl_WD1_t1 = RG_zz_24 ;	// line#=../rle.cpp:74
	6'h1a :
		rl_WD1_t1 = RG_zz_25 ;	// line#=../rle.cpp:74
	6'h1b :
		rl_WD1_t1 = RG_zz_26 ;	// line#=../rle.cpp:74
	6'h1c :
		rl_WD1_t1 = RG_zz_27 ;	// line#=../rle.cpp:74
	6'h1d :
		rl_WD1_t1 = RG_zz_28 ;	// line#=../rle.cpp:74
	6'h1e :
		rl_WD1_t1 = RG_zz_29 ;	// line#=../rle.cpp:74
	6'h1f :
		rl_WD1_t1 = RG_zz_30 ;	// line#=../rle.cpp:74
	6'h20 :
		rl_WD1_t1 = RG_zz_31 ;	// line#=../rle.cpp:74
	6'h21 :
		rl_WD1_t1 = RG_zz_32 ;	// line#=../rle.cpp:74
	6'h22 :
		rl_WD1_t1 = RG_zz_33 ;	// line#=../rle.cpp:74
	6'h23 :
		rl_WD1_t1 = RG_zz_34 ;	// line#=../rle.cpp:74
	6'h24 :
		rl_WD1_t1 = RG_zz_35 ;	// line#=../rle.cpp:74
	6'h25 :
		rl_WD1_t1 = RG_zz_36 ;	// line#=../rle.cpp:74
	6'h26 :
		rl_WD1_t1 = RG_zz_37 ;	// line#=../rle.cpp:74
	6'h27 :
		rl_WD1_t1 = RG_zz_38 ;	// line#=../rle.cpp:74
	6'h28 :
		rl_WD1_t1 = RG_zz_39 ;	// line#=../rle.cpp:74
	6'h29 :
		rl_WD1_t1 = RG_zz_40 ;	// line#=../rle.cpp:74
	6'h2a :
		rl_WD1_t1 = RG_zz_41 ;	// line#=../rle.cpp:74
	6'h2b :
		rl_WD1_t1 = RG_zz_42 ;	// line#=../rle.cpp:74
	6'h2c :
		rl_WD1_t1 = RG_zz_43 ;	// line#=../rle.cpp:74
	6'h2d :
		rl_WD1_t1 = RG_zz_44 ;	// line#=../rle.cpp:74
	6'h2e :
		rl_WD1_t1 = RG_zz_45 ;	// line#=../rle.cpp:74
	6'h2f :
		rl_WD1_t1 = RG_zz_46 ;	// line#=../rle.cpp:74
	6'h30 :
		rl_WD1_t1 = RG_zz_47 ;	// line#=../rle.cpp:74
	6'h31 :
		rl_WD1_t1 = RG_zz_48 ;	// line#=../rle.cpp:74
	6'h32 :
		rl_WD1_t1 = RG_zz_49 ;	// line#=../rle.cpp:74
	6'h33 :
		rl_WD1_t1 = RG_zz_50 ;	// line#=../rle.cpp:74
	6'h34 :
		rl_WD1_t1 = RG_zz_51 ;	// line#=../rle.cpp:74
	6'h35 :
		rl_WD1_t1 = RG_zz_52 ;	// line#=../rle.cpp:74
	6'h36 :
		rl_WD1_t1 = RG_zz_53 ;	// line#=../rle.cpp:74
	6'h37 :
		rl_WD1_t1 = RG_zz_54 ;	// line#=../rle.cpp:74
	6'h38 :
		rl_WD1_t1 = RG_zz_55 ;	// line#=../rle.cpp:74
	6'h39 :
		rl_WD1_t1 = RG_zz_56 ;	// line#=../rle.cpp:74
	6'h3a :
		rl_WD1_t1 = RG_zz_57 ;	// line#=../rle.cpp:74
	6'h3b :
		rl_WD1_t1 = RG_zz_58 ;	// line#=../rle.cpp:74
	6'h3c :
		rl_WD1_t1 = RG_zz_59 ;	// line#=../rle.cpp:74
	6'h3d :
		rl_WD1_t1 = RG_zz_60 ;	// line#=../rle.cpp:74
	6'h3e :
		rl_WD1_t1 = RG_zz_61 ;	// line#=../rle.cpp:74
	6'h3f :
		rl_WD1_t1 = RG_zz_62 ;	// line#=../rle.cpp:74
	default :
		rl_WD1_t1 = 9'hx ;
	endcase
always @ ( rl_WD1_t1 or U_179 or RG_j_k or U_177 or sub12s_91ot or U_88 )
	rl_WD1 = ( ( { 9{ U_88 } } & sub12s_91ot )	// line#=../rle.cpp:52
		| ( { 9{ U_177 } } & RG_j_k [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ U_179 } } & rl_WD1_t1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:68,69,79,80,85
assign	M_107 = ~|( RG_k ^ 6'h01 ) ;	// line#=../rle.cpp:74,111,142
assign	M_110 = ~|RG_k ;	// line#=../rle.cpp:74,111,142
assign	M_114 = ~|( RG_k ^ 6'h08 ) ;	// line#=../rle.cpp:74,111,142
assign	M_115 = ~|( RG_k ^ 6'h24 ) ;	// line#=../rle.cpp:74,111,142
assign	M_116 = ~|( RG_k ^ 6'h02 ) ;	// line#=../rle.cpp:74,111,142
assign	M_118 = ~|( RG_k ^ 6'h07 ) ;	// line#=../rle.cpp:74,111,142
assign	M_120 = ~|( RG_k ^ 6'h0f ) ;	// line#=../rle.cpp:74,111,142
assign	M_122 = ~|( RG_k ^ 6'h04 ) ;	// line#=../rle.cpp:74,111,142
assign	M_124 = ~|( RG_k ^ 6'h03 ) ;	// line#=../rle.cpp:74,111,142
assign	M_126 = ~|( RG_k ^ 6'h05 ) ;	// line#=../rle.cpp:74,111,142
assign	M_128 = ~|( RG_k ^ 6'h06 ) ;	// line#=../rle.cpp:74,111,142
assign	M_130 = ~|( RG_k ^ 6'h3f ) ;	// line#=../rle.cpp:74,111,142
assign	M_131 = ~|( RG_k ^ 6'h3e ) ;	// line#=../rle.cpp:74,111,142
assign	M_132 = ~|( RG_k ^ 6'h3d ) ;	// line#=../rle.cpp:74,111,142
assign	M_133 = ~|( RG_k ^ 6'h3c ) ;	// line#=../rle.cpp:74,111,142
assign	M_134 = ~|( RG_k ^ 6'h3b ) ;	// line#=../rle.cpp:74,111,142
assign	M_135 = ~|( RG_k ^ 6'h3a ) ;	// line#=../rle.cpp:74,111,142
assign	M_136 = ~|( RG_k ^ 6'h39 ) ;	// line#=../rle.cpp:74,111,142
assign	M_137 = ~|( RG_k ^ 6'h38 ) ;	// line#=../rle.cpp:74,111,142
assign	M_138 = ~|( RG_k ^ 6'h37 ) ;	// line#=../rle.cpp:74,111,142
assign	M_139 = ~|( RG_k ^ 6'h36 ) ;	// line#=../rle.cpp:74,111,142
assign	M_140 = ~|( RG_k ^ 6'h35 ) ;	// line#=../rle.cpp:74,111,142
assign	M_141 = ~|( RG_k ^ 6'h34 ) ;	// line#=../rle.cpp:74,111,142
assign	M_142 = ~|( RG_k ^ 6'h33 ) ;	// line#=../rle.cpp:74,111,142
assign	M_143 = ~|( RG_k ^ 6'h32 ) ;	// line#=../rle.cpp:74,111,142
assign	M_144 = ~|( RG_k ^ 6'h31 ) ;	// line#=../rle.cpp:74,111,142
assign	M_145 = ~|( RG_k ^ 6'h30 ) ;	// line#=../rle.cpp:74,111,142
assign	M_146 = ~|( RG_k ^ 6'h2f ) ;	// line#=../rle.cpp:74,111,142
assign	M_147 = ~|( RG_k ^ 6'h2e ) ;	// line#=../rle.cpp:74,111,142
assign	M_148 = ~|( RG_k ^ 6'h2d ) ;	// line#=../rle.cpp:74,111,142
assign	M_149 = ~|( RG_k ^ 6'h2c ) ;	// line#=../rle.cpp:74,111,142
assign	M_150 = ~|( RG_k ^ 6'h2b ) ;	// line#=../rle.cpp:74,111,142
assign	M_151 = ~|( RG_k ^ 6'h2a ) ;	// line#=../rle.cpp:74,111,142
assign	M_152 = ~|( RG_k ^ 6'h29 ) ;	// line#=../rle.cpp:74,111,142
assign	M_153 = ~|( RG_k ^ 6'h28 ) ;	// line#=../rle.cpp:74,111,142
assign	M_154 = ~|( RG_k ^ 6'h27 ) ;	// line#=../rle.cpp:74,111,142
assign	M_155 = ~|( RG_k ^ 6'h26 ) ;	// line#=../rle.cpp:74,111,142
assign	M_156 = ~|( RG_k ^ 6'h25 ) ;	// line#=../rle.cpp:74,111,142
assign	M_157 = ~|( RG_k ^ 6'h23 ) ;	// line#=../rle.cpp:74,111,142
assign	M_158 = ~|( RG_k ^ 6'h22 ) ;	// line#=../rle.cpp:74,111,142
assign	M_159 = ~|( RG_k ^ 6'h21 ) ;	// line#=../rle.cpp:74,111,142
assign	M_160 = ~|( RG_k ^ 6'h20 ) ;	// line#=../rle.cpp:74,111,142
assign	M_161 = ~|( RG_k ^ 6'h1f ) ;	// line#=../rle.cpp:74,111,142
assign	M_162 = ~|( RG_k ^ 6'h1e ) ;	// line#=../rle.cpp:74,111,142
assign	M_163 = ~|( RG_k ^ 6'h1d ) ;	// line#=../rle.cpp:74,111,142
assign	M_164 = ~|( RG_k ^ 6'h1c ) ;	// line#=../rle.cpp:74,111,142
assign	M_165 = ~|( RG_k ^ 6'h1b ) ;	// line#=../rle.cpp:74,111,142
assign	M_166 = ~|( RG_k ^ 6'h1a ) ;	// line#=../rle.cpp:74,111,142
assign	M_167 = ~|( RG_k ^ 6'h19 ) ;	// line#=../rle.cpp:74,111,142
assign	M_168 = ~|( RG_k ^ 6'h18 ) ;	// line#=../rle.cpp:74,111,142
assign	M_169 = ~|( RG_k ^ 6'h17 ) ;	// line#=../rle.cpp:74,111,142
assign	M_170 = ~|( RG_k ^ 6'h16 ) ;	// line#=../rle.cpp:74,111,142
assign	M_171 = ~|( RG_k ^ 6'h15 ) ;	// line#=../rle.cpp:74,111,142
assign	M_172 = ~|( RG_k ^ 6'h14 ) ;	// line#=../rle.cpp:74,111,142
assign	M_173 = ~|( RG_k ^ 6'h13 ) ;	// line#=../rle.cpp:74,111,142
assign	M_174 = ~|( RG_k ^ 6'h12 ) ;	// line#=../rle.cpp:74,111,142
assign	M_175 = ~|( RG_k ^ 6'h11 ) ;	// line#=../rle.cpp:74,111,142
assign	M_176 = ~|( RG_k ^ 6'h10 ) ;	// line#=../rle.cpp:74,111,142
assign	M_177 = ~|( RG_k ^ 6'h0e ) ;	// line#=../rle.cpp:74,111,142
assign	M_178 = ~|( RG_k ^ 6'h0d ) ;	// line#=../rle.cpp:74,111,142
assign	M_179 = ~|( RG_k ^ 6'h0c ) ;	// line#=../rle.cpp:74,111,142
assign	M_180 = ~|( RG_k ^ 6'h0b ) ;	// line#=../rle.cpp:74,111,142
assign	M_181 = ~|( RG_k ^ 6'h0a ) ;	// line#=../rle.cpp:74,111,142
assign	M_182 = ~|( RG_k ^ 6'h09 ) ;	// line#=../rle.cpp:74,111,142
assign	rl_WE1 = ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	U_88 | U_175 ) | ( U_179 & M_130 ) ) | ( U_179 & M_131 ) ) | ( U_179 & M_132 ) ) | 
	( U_179 & M_133 ) ) | ( U_179 & M_134 ) ) | ( U_179 & M_135 ) ) | ( U_179 & 
	M_136 ) ) | ( U_179 & M_137 ) ) | ( U_179 & M_138 ) ) | ( U_179 & M_139 ) ) | 
	( U_179 & M_140 ) ) | ( U_179 & M_141 ) ) | ( U_179 & M_142 ) ) | ( U_179 & 
	M_143 ) ) | ( U_179 & M_144 ) ) | ( U_179 & M_145 ) ) | ( U_179 & M_146 ) ) | 
	( U_179 & M_147 ) ) | ( U_179 & M_148 ) ) | ( U_179 & M_149 ) ) | ( U_179 & 
	M_150 ) ) | ( U_179 & M_151 ) ) | ( U_179 & M_152 ) ) | ( U_179 & M_153 ) ) | 
	( U_179 & M_154 ) ) | ( U_179 & M_155 ) ) | ( U_179 & M_156 ) ) | ( U_179 & 
	M_115 ) ) | ( U_179 & M_157 ) ) | ( U_179 & M_158 ) ) | ( U_179 & M_159 ) ) | 
	( U_179 & M_160 ) ) | ( U_179 & M_161 ) ) | ( U_179 & M_162 ) ) | ( U_179 & 
	M_163 ) ) | ( U_179 & M_164 ) ) | ( U_179 & M_165 ) ) | ( U_179 & M_166 ) ) | 
	( U_179 & M_167 ) ) | ( U_179 & M_168 ) ) | ( U_179 & M_169 ) ) | ( U_179 & 
	M_170 ) ) | ( U_179 & M_171 ) ) | ( U_179 & M_172 ) ) | ( U_179 & M_173 ) ) | 
	( U_179 & M_174 ) ) | ( U_179 & M_175 ) ) | ( U_179 & M_176 ) ) | ( U_179 & 
	M_120 ) ) | ( U_179 & M_177 ) ) | ( U_179 & M_178 ) ) | ( U_179 & M_179 ) ) | 
	( U_179 & M_180 ) ) | ( U_179 & M_181 ) ) | ( U_179 & M_182 ) ) | ( U_179 & 
	M_114 ) ) | ( U_179 & M_118 ) ) | ( U_179 & M_128 ) ) | ( U_179 & M_126 ) ) | 
	( U_179 & M_122 ) ) | ( U_179 & M_124 ) ) | ( U_179 & M_116 ) ) | ( U_179 & 
	M_107 ) ) | ( U_179 & M_110 ) ) | U_178 ) | U_248 ) | ST1_10d ) | U_257 ) ;
always @ ( ST1_52d or ST1_50d or ST1_48d or ST1_46d or ST1_44d or ST1_42d or ST1_40d or 
	ST1_38d or ST1_36d or ST1_34d or ST1_31d or ST1_29d or ST1_27d or ST1_25d or 
	ST1_23d or ST1_21d or ST1_19d or ST1_17d or ST1_15d or ST1_13d or ST1_12d )
	TR_12 = ( ( { 6{ ST1_12d } } & 6'h01 )
		| ( { 6{ ST1_13d } } & 6'h02 )
		| ( { 6{ ST1_15d } } & 6'h05 )
		| ( { 6{ ST1_17d } } & 6'h08 )
		| ( { 6{ ST1_19d } } & 6'h0b )
		| ( { 6{ ST1_21d } } & 6'h0e )
		| ( { 6{ ST1_23d } } & 6'h11 )
		| ( { 6{ ST1_25d } } & 6'h14 )
		| ( { 6{ ST1_27d } } & 6'h17 )
		| ( { 6{ ST1_29d } } & 6'h1a )
		| ( { 6{ ST1_31d } } & 6'h1d )
		| ( { 6{ ST1_34d } } & 6'h21 )
		| ( { 6{ ST1_36d } } & 6'h24 )
		| ( { 6{ ST1_38d } } & 6'h27 )
		| ( { 6{ ST1_40d } } & 6'h2a )
		| ( { 6{ ST1_42d } } & 6'h2d )
		| ( { 6{ ST1_44d } } & 6'h30 )
		| ( { 6{ ST1_46d } } & 6'h33 )
		| ( { 6{ ST1_48d } } & 6'h36 )
		| ( { 6{ ST1_50d } } & 6'h39 )
		| ( { 6{ ST1_52d } } & 6'h3c ) ) ;
always @ ( ST1_54d or ST1_53d or ST1_51d or ST1_49d or ST1_47d or ST1_45d or ST1_43d or 
	ST1_41d or ST1_39d or ST1_37d or ST1_35d or ST1_33d or ST1_32d or ST1_30d or 
	ST1_28d or ST1_26d or ST1_24d or ST1_22d or ST1_20d or ST1_18d or ST1_16d or 
	ST1_14d )
	TR_13 = ( ( { 6{ ST1_14d } } & 6'h03 )
		| ( { 6{ ST1_16d } } & 6'h06 )
		| ( { 6{ ST1_18d } } & 6'h09 )
		| ( { 6{ ST1_20d } } & 6'h0c )
		| ( { 6{ ST1_22d } } & 6'h0f )
		| ( { 6{ ST1_24d } } & 6'h12 )
		| ( { 6{ ST1_26d } } & 6'h15 )
		| ( { 6{ ST1_28d } } & 6'h18 )
		| ( { 6{ ST1_30d } } & 6'h1b )
		| ( { 6{ ST1_32d } } & 6'h1e )
		| ( { 6{ ST1_33d } } & 6'h1f )
		| ( { 6{ ST1_35d } } & 6'h22 )
		| ( { 6{ ST1_37d } } & 6'h25 )
		| ( { 6{ ST1_39d } } & 6'h28 )
		| ( { 6{ ST1_41d } } & 6'h2b )
		| ( { 6{ ST1_43d } } & 6'h2e )
		| ( { 6{ ST1_45d } } & 6'h31 )
		| ( { 6{ ST1_47d } } & 6'h34 )
		| ( { 6{ ST1_49d } } & 6'h37 )
		| ( { 6{ ST1_51d } } & 6'h3a )
		| ( { 6{ ST1_53d } } & 6'h3d )
		| ( { 6{ ST1_54d } } & 6'h3f ) ) ;
always @ ( TR_13 or ST1_54d or M_195 or TR_12 or M_192 or RG_142_01 or M_188 )
	begin
	rl_RA2_c1 = ( M_195 | ST1_54d ) ;
	rl_RA2 = ( ( { 7{ M_188 } } & RG_142_01 )
		| ( { 7{ M_192 } } & { TR_12 , 1'h0 } )
		| ( { 7{ rl_RA2_c1 } } & { TR_13 , 1'h1 } ) ) ;
	end
always @ ( ST1_52d or ST1_50d or ST1_48d or ST1_46d or ST1_44d or ST1_42d or ST1_40d or 
	ST1_38d or ST1_36d or ST1_34d or ST1_31d or ST1_29d or ST1_27d or ST1_25d or 
	ST1_23d or ST1_21d or ST1_19d or ST1_17d or ST1_15d or ST1_13d )
	TR_14 = ( ( { 6{ ST1_13d } } & 6'h01 )
		| ( { 6{ ST1_15d } } & 6'h04 )
		| ( { 6{ ST1_17d } } & 6'h07 )
		| ( { 6{ ST1_19d } } & 6'h0a )
		| ( { 6{ ST1_21d } } & 6'h0d )
		| ( { 6{ ST1_23d } } & 6'h10 )
		| ( { 6{ ST1_25d } } & 6'h13 )
		| ( { 6{ ST1_27d } } & 6'h16 )
		| ( { 6{ ST1_29d } } & 6'h19 )
		| ( { 6{ ST1_31d } } & 6'h1c )
		| ( { 6{ ST1_34d } } & 6'h21 )
		| ( { 6{ ST1_36d } } & 6'h24 )
		| ( { 6{ ST1_38d } } & 6'h27 )
		| ( { 6{ ST1_40d } } & 6'h2a )
		| ( { 6{ ST1_42d } } & 6'h2d )
		| ( { 6{ ST1_44d } } & 6'h30 )
		| ( { 6{ ST1_46d } } & 6'h33 )
		| ( { 6{ ST1_48d } } & 6'h36 )
		| ( { 6{ ST1_50d } } & 6'h39 )
		| ( { 6{ ST1_52d } } & 6'h3c ) ) ;
always @ ( ST1_53d or ST1_51d or ST1_49d or ST1_47d or ST1_45d or ST1_43d or ST1_41d or 
	ST1_39d or ST1_37d or ST1_35d or ST1_33d or ST1_32d or ST1_30d or ST1_28d or 
	ST1_26d or ST1_24d or ST1_22d or ST1_20d or ST1_18d or ST1_16d or ST1_14d )
	TR_15 = ( ( { 6{ ST1_14d } } & 6'h03 )
		| ( { 6{ ST1_16d } } & 6'h06 )
		| ( { 6{ ST1_18d } } & 6'h09 )
		| ( { 6{ ST1_20d } } & 6'h0c )
		| ( { 6{ ST1_22d } } & 6'h0f )
		| ( { 6{ ST1_24d } } & 6'h12 )
		| ( { 6{ ST1_26d } } & 6'h15 )
		| ( { 6{ ST1_28d } } & 6'h18 )
		| ( { 6{ ST1_30d } } & 6'h1b )
		| ( { 6{ ST1_32d } } & 6'h1e )
		| ( { 6{ ST1_33d } } & 6'h20 )
		| ( { 6{ ST1_35d } } & 6'h23 )
		| ( { 6{ ST1_37d } } & 6'h26 )
		| ( { 6{ ST1_39d } } & 6'h29 )
		| ( { 6{ ST1_41d } } & 6'h2c )
		| ( { 6{ ST1_43d } } & 6'h2f )
		| ( { 6{ ST1_45d } } & 6'h32 )
		| ( { 6{ ST1_47d } } & 6'h35 )
		| ( { 6{ ST1_49d } } & 6'h38 )
		| ( { 6{ ST1_51d } } & 6'h3b )
		| ( { 6{ ST1_53d } } & 6'h3e ) ) ;
assign	M_192 = ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ST1_12d | ST1_13d ) | ST1_15d ) | 
	ST1_17d ) | ST1_19d ) | ST1_21d ) | ST1_23d ) | ST1_25d ) | ST1_27d ) | ST1_29d ) | 
	ST1_31d ) | ST1_34d ) | ST1_36d ) | ST1_38d ) | ST1_40d ) | ST1_42d ) | ST1_44d ) | 
	ST1_46d ) | ST1_48d ) | ST1_50d ) | ST1_52d ) ;
assign	M_195 = ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ST1_14d | ST1_16d ) | ST1_18d ) | 
	ST1_20d ) | ST1_22d ) | ST1_24d ) | ST1_26d ) | ST1_28d ) | ST1_30d ) | ST1_32d ) | 
	ST1_33d ) | ST1_35d ) | ST1_37d ) | ST1_39d ) | ST1_41d ) | ST1_43d ) | ST1_45d ) | 
	ST1_47d ) | ST1_49d ) | ST1_51d ) | ST1_53d ) ;
always @ ( TR_15 or M_195 or TR_14 or M_192 or RG_k_01 or M_188 )
	rl_RA3 = ( ( { 7{ M_188 } } & RG_k_01 )	// line#=../rle.cpp:77,78,83,84
		| ( { 7{ M_192 } } & { TR_14 , 1'h1 } )
		| ( { 7{ M_195 } } & { TR_15 , 1'h0 } ) ) ;

endmodule

module jpeg_sub8u_7_1 ( i1 ,i2 ,o1 );
input	[6:0]	i1 ;
input	[1:0]	i2 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - { 5'h00 , i2 } ) ;

endmodule

module jpeg_sub8u_7 ( i1 ,i2 ,o1 );
input	[6:0]	i1 ;
input	[2:0]	i2 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - { 4'h0 , i2 } ) ;

endmodule

module jpeg_decr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_decr8u_7 ( i1 ,o1 );
input	[6:0]	i1 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_incr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr8u ( i1 ,o1 );
input	[7:0]	i1 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr4s ( i1 ,o1 );
input	[3:0]	i1 ;
output	[3:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_lop8u_1 ( i1 ,i2 ,o1 );
input	[5:0]	i1 ;
input	[5:0]	i2 ;
output		o1 ;
wire		M_01 ;

assign	M_01 = ( i1 < i2 ) ;
assign	o1 = M_01 ;

endmodule

module jpeg_sub12s_9 ( i1 ,i2 ,o1 );
input	[8:0]	i1 ;
input	[8:0]	i2 ;
output	[8:0]	o1 ;

assign	o1 = ( i1 - i2 ) ;

endmodule

module jpeg_sub8u ( i1 ,i2 ,o1 );
input	[7:0]	i1 ;
input	[1:0]	i2 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 - { 6'h00 , i2 } ) ;

endmodule

module jpeg_MEM_rl ( AD1 ,RD1 ,WD1 ,WE1 ,CLK1 ,RA2 ,RD2 ,RA3 ,RD3 );
input	[6:0]	AD1 ;
output	[8:0]	RD1 ;
input	[8:0]	WD1 ;
input		WE1 ;
input		CLK1 ;
input	[6:0]	RA2 ;
output	[8:0]	RD2 ;
input	[6:0]	RA3 ;
output	[8:0]	RD3 ;

jpeg_MEM_rl_subD INST_MEM_rl_subD_1 ( .RD1(RD1) ,.AD1(AD1) ,.WE1(WE1) ,.WD1(WD1) ,
	.CLK1(CLK1) ,.RD2(RD2) ,.RA2(RA2) );
jpeg_MEM_rl_subD INST_MEM_rl_subD_2 ( .RD1() ,.AD1(AD1) ,.WE1(WE1) ,.WD1(WD1) ,.CLK1(CLK1) ,
	.RD2(RD3) ,.RA2(RA3) );

endmodule

(* ram_extract = "yes" *)
module jpeg_MEM_rl_subD ( RD1 ,AD1 ,WE1 ,WD1 ,CLK1 ,RD2 ,RA2 );
output	[8:0]	RD1 ;
input	[6:0]	AD1 ;
input		WE1 ;
input	[8:0]	WD1 ;
input		CLK1 ;
output	[8:0]	RD2 ;
input	[6:0]	RA2 ;
(* ram_style = "distributed" *)reg	[8:0]	rl_r	[0:127] ;

assign	RD1 = rl_r[AD1] ;
assign	RD2 = rl_r[RA2] ;

always @ ( posedge CLK1 )
	begin
	if ( WE1 )
		rl_r [AD1] = WD1 ;
	end

endmodule
