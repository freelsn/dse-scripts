// verilog_out version 6.79.2
// options:  veriloggen jpeg_E.IFF
// bdlpars options:  -DDSE ../rle.cpp
// bdltran options:  -c1000 -s -Zresource_fcnt=GENERATE -Zresource_mcnt=GENERATE -lb /home/shuangnan/share/packages/zynq-1.BLIB -lfl /home/shuangnan/share/packages/zynq-1.FLIB jpeg.IFF -OX -a8196 -Zfu_cnt_incr_rate=0 -tcio 
// timestamp_0: 20180213184527_31358_33285
// timestamp_5: 20180213184531_32298_73001
// timestamp_9: 20180213184836_32298_37333
// timestamp_C: 20180213184830_32298_74311
// timestamp_E: 20180213184844_32298_15814
// timestamp_V: 20180213184912_26970_83364

module jpeg ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,jpeg_in_a04 ,
	jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,jpeg_in_a10 ,
	jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,jpeg_in_a16 ,
	jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,jpeg_in_a22 ,
	jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,jpeg_in_a28 ,
	jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,jpeg_in_a34 ,
	jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,jpeg_in_a40 ,
	jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,jpeg_in_a46 ,
	jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,jpeg_in_a52 ,
	jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,jpeg_in_a58 ,
	jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,jpeg_in_a64 ,
	jpeg_in_a65 ,jpeg_in_a66 ,jpeg_in_a67 ,jpeg_in_a68 ,jpeg_in_a69 ,jpeg_in_a70 ,
	jpeg_in_a71 ,jpeg_in_a72 ,jpeg_in_a73 ,jpeg_in_a74 ,jpeg_in_a75 ,jpeg_in_a76 ,
	jpeg_in_a77 ,jpeg_in_a78 ,jpeg_in_a79 ,jpeg_in_a80 ,jpeg_in_a81 ,jpeg_in_a82 ,
	jpeg_in_a83 ,jpeg_in_a84 ,jpeg_in_a85 ,jpeg_in_a86 ,jpeg_in_a87 ,jpeg_in_a88 ,
	jpeg_in_a89 ,jpeg_in_a90 ,jpeg_in_a91 ,jpeg_in_a92 ,jpeg_in_a93 ,jpeg_in_a94 ,
	jpeg_in_a95 ,jpeg_in_a96 ,jpeg_in_a97 ,jpeg_in_a98 ,jpeg_in_a99 ,jpeg_in_a100 ,
	jpeg_in_a101 ,jpeg_in_a102 ,jpeg_in_a103 ,jpeg_in_a104 ,jpeg_in_a105 ,jpeg_in_a106 ,
	jpeg_in_a107 ,jpeg_in_a108 ,jpeg_in_a109 ,jpeg_in_a110 ,jpeg_in_a111 ,jpeg_in_a112 ,
	jpeg_in_a113 ,jpeg_in_a114 ,jpeg_in_a115 ,jpeg_in_a116 ,jpeg_in_a117 ,jpeg_in_a118 ,
	jpeg_in_a119 ,jpeg_in_a120 ,jpeg_in_a121 ,jpeg_in_a122 ,jpeg_in_a123 ,jpeg_in_a124 ,
	jpeg_in_a125 ,jpeg_in_a126 ,jpeg_in_a127 ,jpeg_len_in ,jpeg_out_a00 ,jpeg_out_a01 ,
	jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,jpeg_out_a06 ,jpeg_out_a07 ,
	jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,jpeg_out_a12 ,jpeg_out_a13 ,
	jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,jpeg_out_a18 ,jpeg_out_a19 ,
	jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,jpeg_out_a24 ,jpeg_out_a25 ,
	jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,jpeg_out_a30 ,jpeg_out_a31 ,
	jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,jpeg_out_a36 ,jpeg_out_a37 ,
	jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,jpeg_out_a42 ,jpeg_out_a43 ,
	jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,jpeg_out_a48 ,jpeg_out_a49 ,
	jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,jpeg_out_a54 ,jpeg_out_a55 ,
	jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,jpeg_out_a60 ,jpeg_out_a61 ,
	jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,jpeg_out_a66 ,jpeg_out_a67 ,
	jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,jpeg_out_a72 ,jpeg_out_a73 ,
	jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,jpeg_out_a78 ,jpeg_out_a79 ,
	jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,jpeg_out_a84 ,jpeg_out_a85 ,
	jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,jpeg_out_a90 ,jpeg_out_a91 ,
	jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,jpeg_out_a96 ,jpeg_out_a97 ,
	jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,jpeg_out_a102 ,
	jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,jpeg_out_a107 ,
	jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,jpeg_out_a112 ,
	jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,jpeg_out_a117 ,
	jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,jpeg_out_a122 ,
	jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,jpeg_out_a127 ,
	jpeg_len_out ,valid );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a64 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a65 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a66 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a67 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a68 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a69 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a70 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a71 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a72 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a73 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a74 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a75 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a76 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a77 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a78 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a79 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a80 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a81 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a82 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a83 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a84 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a85 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a86 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a87 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a88 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a89 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a90 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a91 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a92 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a93 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a94 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a95 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a96 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a97 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a98 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a99 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a100 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a101 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a102 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a103 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a104 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a105 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a106 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a107 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a108 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a109 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a110 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a111 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a112 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a113 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a114 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a115 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a116 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a117 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a118 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a119 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a120 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a121 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a122 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a123 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a124 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a125 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a126 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a127 ;	// line#=../rle.h:56
input	[11:0]	jpeg_len_in ;	// line#=../rle.h:57
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
wire		ST1_01d ;
wire		ST1_02d ;
wire		ST1_03d ;
wire		ST1_04d ;
wire		ST1_05d ;
wire		ST1_06d ;
wire		ST1_07d ;
wire		ST1_08d ;
wire		JF_01 ;
wire		lop8u_11ot ;
wire		JF_03 ;
wire		C_07 ;
wire		C_08 ;
wire		JF_06 ;

jpeg_fsm INST_fsm ( .clk(clk) ,.rst(rst) ,.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,
	.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,
	.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,.JF_01(JF_01) ,.lop8u_11ot(lop8u_11ot) ,
	.JF_03(JF_03) ,.C_07(C_07) ,.C_08(C_08) ,.JF_06(JF_06) );
jpeg_dat INST_dat ( .clk(clk) ,.rst(rst) ,.jpeg_in_a00(jpeg_in_a00) ,.jpeg_in_a01(jpeg_in_a01) ,
	.jpeg_in_a02(jpeg_in_a02) ,.jpeg_in_a03(jpeg_in_a03) ,.jpeg_in_a04(jpeg_in_a04) ,
	.jpeg_in_a05(jpeg_in_a05) ,.jpeg_in_a06(jpeg_in_a06) ,.jpeg_in_a07(jpeg_in_a07) ,
	.jpeg_in_a08(jpeg_in_a08) ,.jpeg_in_a09(jpeg_in_a09) ,.jpeg_in_a10(jpeg_in_a10) ,
	.jpeg_in_a11(jpeg_in_a11) ,.jpeg_in_a12(jpeg_in_a12) ,.jpeg_in_a13(jpeg_in_a13) ,
	.jpeg_in_a14(jpeg_in_a14) ,.jpeg_in_a15(jpeg_in_a15) ,.jpeg_in_a16(jpeg_in_a16) ,
	.jpeg_in_a17(jpeg_in_a17) ,.jpeg_in_a18(jpeg_in_a18) ,.jpeg_in_a19(jpeg_in_a19) ,
	.jpeg_in_a20(jpeg_in_a20) ,.jpeg_in_a21(jpeg_in_a21) ,.jpeg_in_a22(jpeg_in_a22) ,
	.jpeg_in_a23(jpeg_in_a23) ,.jpeg_in_a24(jpeg_in_a24) ,.jpeg_in_a25(jpeg_in_a25) ,
	.jpeg_in_a26(jpeg_in_a26) ,.jpeg_in_a27(jpeg_in_a27) ,.jpeg_in_a28(jpeg_in_a28) ,
	.jpeg_in_a29(jpeg_in_a29) ,.jpeg_in_a30(jpeg_in_a30) ,.jpeg_in_a31(jpeg_in_a31) ,
	.jpeg_in_a32(jpeg_in_a32) ,.jpeg_in_a33(jpeg_in_a33) ,.jpeg_in_a34(jpeg_in_a34) ,
	.jpeg_in_a35(jpeg_in_a35) ,.jpeg_in_a36(jpeg_in_a36) ,.jpeg_in_a37(jpeg_in_a37) ,
	.jpeg_in_a38(jpeg_in_a38) ,.jpeg_in_a39(jpeg_in_a39) ,.jpeg_in_a40(jpeg_in_a40) ,
	.jpeg_in_a41(jpeg_in_a41) ,.jpeg_in_a42(jpeg_in_a42) ,.jpeg_in_a43(jpeg_in_a43) ,
	.jpeg_in_a44(jpeg_in_a44) ,.jpeg_in_a45(jpeg_in_a45) ,.jpeg_in_a46(jpeg_in_a46) ,
	.jpeg_in_a47(jpeg_in_a47) ,.jpeg_in_a48(jpeg_in_a48) ,.jpeg_in_a49(jpeg_in_a49) ,
	.jpeg_in_a50(jpeg_in_a50) ,.jpeg_in_a51(jpeg_in_a51) ,.jpeg_in_a52(jpeg_in_a52) ,
	.jpeg_in_a53(jpeg_in_a53) ,.jpeg_in_a54(jpeg_in_a54) ,.jpeg_in_a55(jpeg_in_a55) ,
	.jpeg_in_a56(jpeg_in_a56) ,.jpeg_in_a57(jpeg_in_a57) ,.jpeg_in_a58(jpeg_in_a58) ,
	.jpeg_in_a59(jpeg_in_a59) ,.jpeg_in_a60(jpeg_in_a60) ,.jpeg_in_a61(jpeg_in_a61) ,
	.jpeg_in_a62(jpeg_in_a62) ,.jpeg_in_a63(jpeg_in_a63) ,.jpeg_out_a00(jpeg_out_a00) ,
	.jpeg_out_a01(jpeg_out_a01) ,.jpeg_out_a02(jpeg_out_a02) ,.jpeg_out_a03(jpeg_out_a03) ,
	.jpeg_out_a04(jpeg_out_a04) ,.jpeg_out_a05(jpeg_out_a05) ,.jpeg_out_a06(jpeg_out_a06) ,
	.jpeg_out_a07(jpeg_out_a07) ,.jpeg_out_a08(jpeg_out_a08) ,.jpeg_out_a09(jpeg_out_a09) ,
	.jpeg_out_a10(jpeg_out_a10) ,.jpeg_out_a11(jpeg_out_a11) ,.jpeg_out_a12(jpeg_out_a12) ,
	.jpeg_out_a13(jpeg_out_a13) ,.jpeg_out_a14(jpeg_out_a14) ,.jpeg_out_a15(jpeg_out_a15) ,
	.jpeg_out_a16(jpeg_out_a16) ,.jpeg_out_a17(jpeg_out_a17) ,.jpeg_out_a18(jpeg_out_a18) ,
	.jpeg_out_a19(jpeg_out_a19) ,.jpeg_out_a20(jpeg_out_a20) ,.jpeg_out_a21(jpeg_out_a21) ,
	.jpeg_out_a22(jpeg_out_a22) ,.jpeg_out_a23(jpeg_out_a23) ,.jpeg_out_a24(jpeg_out_a24) ,
	.jpeg_out_a25(jpeg_out_a25) ,.jpeg_out_a26(jpeg_out_a26) ,.jpeg_out_a27(jpeg_out_a27) ,
	.jpeg_out_a28(jpeg_out_a28) ,.jpeg_out_a29(jpeg_out_a29) ,.jpeg_out_a30(jpeg_out_a30) ,
	.jpeg_out_a31(jpeg_out_a31) ,.jpeg_out_a32(jpeg_out_a32) ,.jpeg_out_a33(jpeg_out_a33) ,
	.jpeg_out_a34(jpeg_out_a34) ,.jpeg_out_a35(jpeg_out_a35) ,.jpeg_out_a36(jpeg_out_a36) ,
	.jpeg_out_a37(jpeg_out_a37) ,.jpeg_out_a38(jpeg_out_a38) ,.jpeg_out_a39(jpeg_out_a39) ,
	.jpeg_out_a40(jpeg_out_a40) ,.jpeg_out_a41(jpeg_out_a41) ,.jpeg_out_a42(jpeg_out_a42) ,
	.jpeg_out_a43(jpeg_out_a43) ,.jpeg_out_a44(jpeg_out_a44) ,.jpeg_out_a45(jpeg_out_a45) ,
	.jpeg_out_a46(jpeg_out_a46) ,.jpeg_out_a47(jpeg_out_a47) ,.jpeg_out_a48(jpeg_out_a48) ,
	.jpeg_out_a49(jpeg_out_a49) ,.jpeg_out_a50(jpeg_out_a50) ,.jpeg_out_a51(jpeg_out_a51) ,
	.jpeg_out_a52(jpeg_out_a52) ,.jpeg_out_a53(jpeg_out_a53) ,.jpeg_out_a54(jpeg_out_a54) ,
	.jpeg_out_a55(jpeg_out_a55) ,.jpeg_out_a56(jpeg_out_a56) ,.jpeg_out_a57(jpeg_out_a57) ,
	.jpeg_out_a58(jpeg_out_a58) ,.jpeg_out_a59(jpeg_out_a59) ,.jpeg_out_a60(jpeg_out_a60) ,
	.jpeg_out_a61(jpeg_out_a61) ,.jpeg_out_a62(jpeg_out_a62) ,.jpeg_out_a63(jpeg_out_a63) ,
	.jpeg_out_a64(jpeg_out_a64) ,.jpeg_out_a65(jpeg_out_a65) ,.jpeg_out_a66(jpeg_out_a66) ,
	.jpeg_out_a67(jpeg_out_a67) ,.jpeg_out_a68(jpeg_out_a68) ,.jpeg_out_a69(jpeg_out_a69) ,
	.jpeg_out_a70(jpeg_out_a70) ,.jpeg_out_a71(jpeg_out_a71) ,.jpeg_out_a72(jpeg_out_a72) ,
	.jpeg_out_a73(jpeg_out_a73) ,.jpeg_out_a74(jpeg_out_a74) ,.jpeg_out_a75(jpeg_out_a75) ,
	.jpeg_out_a76(jpeg_out_a76) ,.jpeg_out_a77(jpeg_out_a77) ,.jpeg_out_a78(jpeg_out_a78) ,
	.jpeg_out_a79(jpeg_out_a79) ,.jpeg_out_a80(jpeg_out_a80) ,.jpeg_out_a81(jpeg_out_a81) ,
	.jpeg_out_a82(jpeg_out_a82) ,.jpeg_out_a83(jpeg_out_a83) ,.jpeg_out_a84(jpeg_out_a84) ,
	.jpeg_out_a85(jpeg_out_a85) ,.jpeg_out_a86(jpeg_out_a86) ,.jpeg_out_a87(jpeg_out_a87) ,
	.jpeg_out_a88(jpeg_out_a88) ,.jpeg_out_a89(jpeg_out_a89) ,.jpeg_out_a90(jpeg_out_a90) ,
	.jpeg_out_a91(jpeg_out_a91) ,.jpeg_out_a92(jpeg_out_a92) ,.jpeg_out_a93(jpeg_out_a93) ,
	.jpeg_out_a94(jpeg_out_a94) ,.jpeg_out_a95(jpeg_out_a95) ,.jpeg_out_a96(jpeg_out_a96) ,
	.jpeg_out_a97(jpeg_out_a97) ,.jpeg_out_a98(jpeg_out_a98) ,.jpeg_out_a99(jpeg_out_a99) ,
	.jpeg_out_a100(jpeg_out_a100) ,.jpeg_out_a101(jpeg_out_a101) ,.jpeg_out_a102(jpeg_out_a102) ,
	.jpeg_out_a103(jpeg_out_a103) ,.jpeg_out_a104(jpeg_out_a104) ,.jpeg_out_a105(jpeg_out_a105) ,
	.jpeg_out_a106(jpeg_out_a106) ,.jpeg_out_a107(jpeg_out_a107) ,.jpeg_out_a108(jpeg_out_a108) ,
	.jpeg_out_a109(jpeg_out_a109) ,.jpeg_out_a110(jpeg_out_a110) ,.jpeg_out_a111(jpeg_out_a111) ,
	.jpeg_out_a112(jpeg_out_a112) ,.jpeg_out_a113(jpeg_out_a113) ,.jpeg_out_a114(jpeg_out_a114) ,
	.jpeg_out_a115(jpeg_out_a115) ,.jpeg_out_a116(jpeg_out_a116) ,.jpeg_out_a117(jpeg_out_a117) ,
	.jpeg_out_a118(jpeg_out_a118) ,.jpeg_out_a119(jpeg_out_a119) ,.jpeg_out_a120(jpeg_out_a120) ,
	.jpeg_out_a121(jpeg_out_a121) ,.jpeg_out_a122(jpeg_out_a122) ,.jpeg_out_a123(jpeg_out_a123) ,
	.jpeg_out_a124(jpeg_out_a124) ,.jpeg_out_a125(jpeg_out_a125) ,.jpeg_out_a126(jpeg_out_a126) ,
	.jpeg_out_a127(jpeg_out_a127) ,.jpeg_len_out(jpeg_len_out) ,.valid(valid) ,
	.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,
	.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,
	.JF_01(JF_01) ,.lop8u_11ot_port(lop8u_11ot) ,.JF_03(JF_03) ,.C_07_port(C_07) ,
	.C_08_port(C_08) ,.JF_06(JF_06) );

endmodule

module jpeg_fsm ( clk ,rst ,ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,
	ST1_02d ,ST1_01d ,JF_01 ,lop8u_11ot ,JF_03 ,C_07 ,C_08 ,JF_06 );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
output		ST1_08d ;
output		ST1_07d ;
output		ST1_06d ;
output		ST1_05d ;
output		ST1_04d ;
output		ST1_03d ;
output		ST1_02d ;
output		ST1_01d ;
input		JF_01 ;
input		lop8u_11ot ;
input		JF_03 ;
input		C_07 ;
input		C_08 ;
input		JF_06 ;
reg	[2:0]	B01_streg ;

parameter	ST1_01 = 3'h0 ;
parameter	ST1_02 = 3'h1 ;
parameter	ST1_03 = 3'h2 ;
parameter	ST1_04 = 3'h3 ;
parameter	ST1_05 = 3'h4 ;
parameter	ST1_06 = 3'h5 ;
parameter	ST1_07 = 3'h6 ;
parameter	ST1_08 = 3'h7 ;

assign	ST1_01d = ( ( B01_streg == ST1_01 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_02d = ( ( B01_streg == ST1_02 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_03d = ( ( B01_streg == ST1_03 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_04d = ( ( B01_streg == ST1_04 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_05d = ( ( B01_streg == ST1_05 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_06d = ( ( B01_streg == ST1_06 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_07d = ( ( B01_streg == ST1_07 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_08d = ( ( B01_streg == ST1_08 ) ? 1'h1 : 1'h0 ) ;
always @ ( posedge clk )
	if ( !rst )
		B01_streg <= ST1_01 ;
	else
		case ( B01_streg )
		ST1_01 :
			B01_streg <= ST1_02 ;
		ST1_02 :
			if ( ( JF_01 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_03 ;
		ST1_03 :
			if ( ( lop8u_11ot != 1'h0 ) )
				B01_streg <= ST1_03 ;
			else
				B01_streg <= ST1_04 ;
		ST1_04 :
			if ( ( JF_03 != 1'h0 ) )
				B01_streg <= ST1_04 ;
			else
				B01_streg <= ST1_05 ;
		ST1_05 :
			if ( ( C_07 != 1'h0 ) )
				B01_streg <= ST1_06 ;
			else
				B01_streg <= ST1_07 ;
		ST1_06 :
			if ( ( C_08 != 1'h0 ) )
				B01_streg <= ST1_06 ;
			else
				B01_streg <= ST1_08 ;
		ST1_07 :
			if ( ( JF_06 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_07 ;
		ST1_08 :
			B01_streg <= ST1_05 ;
		default :
			B01_streg <= ST1_01 ;
		endcase

endmodule

module jpeg_dat ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,
	jpeg_in_a04 ,jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,
	jpeg_in_a10 ,jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,
	jpeg_in_a16 ,jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,
	jpeg_in_a22 ,jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,
	jpeg_in_a28 ,jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,
	jpeg_in_a34 ,jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,
	jpeg_in_a40 ,jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,
	jpeg_in_a46 ,jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,
	jpeg_in_a52 ,jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,
	jpeg_in_a58 ,jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,
	jpeg_out_a00 ,jpeg_out_a01 ,jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,
	jpeg_out_a06 ,jpeg_out_a07 ,jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,
	jpeg_out_a12 ,jpeg_out_a13 ,jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,
	jpeg_out_a18 ,jpeg_out_a19 ,jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,
	jpeg_out_a24 ,jpeg_out_a25 ,jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,
	jpeg_out_a30 ,jpeg_out_a31 ,jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,
	jpeg_out_a36 ,jpeg_out_a37 ,jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,
	jpeg_out_a42 ,jpeg_out_a43 ,jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,
	jpeg_out_a48 ,jpeg_out_a49 ,jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,
	jpeg_out_a54 ,jpeg_out_a55 ,jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,
	jpeg_out_a60 ,jpeg_out_a61 ,jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,
	jpeg_out_a66 ,jpeg_out_a67 ,jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,
	jpeg_out_a72 ,jpeg_out_a73 ,jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,
	jpeg_out_a78 ,jpeg_out_a79 ,jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,
	jpeg_out_a84 ,jpeg_out_a85 ,jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,
	jpeg_out_a90 ,jpeg_out_a91 ,jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,
	jpeg_out_a96 ,jpeg_out_a97 ,jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,
	jpeg_out_a102 ,jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,
	jpeg_out_a107 ,jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,
	jpeg_out_a112 ,jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,
	jpeg_out_a117 ,jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,
	jpeg_out_a122 ,jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,
	jpeg_out_a127 ,jpeg_len_out ,valid ,ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,
	ST1_04d ,ST1_03d ,ST1_02d ,ST1_01d ,JF_01 ,lop8u_11ot_port ,JF_03 ,C_07_port ,
	C_08_port ,JF_06 );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
input		ST1_08d ;
input		ST1_07d ;
input		ST1_06d ;
input		ST1_05d ;
input		ST1_04d ;
input		ST1_03d ;
input		ST1_02d ;
input		ST1_01d ;
output		JF_01 ;
output		lop8u_11ot_port ;
output		JF_03 ;
output		C_07_port ;
output		C_08_port ;
output		JF_06 ;
wire		M_183 ;
wire		M_182 ;
wire		M_181 ;
wire		M_180 ;
wire		M_179 ;
wire		M_178 ;
wire		M_177 ;
wire		M_176 ;
wire		M_175 ;
wire		M_174 ;
wire		M_173 ;
wire		M_172 ;
wire		M_171 ;
wire		M_170 ;
wire		M_169 ;
wire		M_168 ;
wire		M_167 ;
wire		M_166 ;
wire		M_165 ;
wire		M_164 ;
wire		M_163 ;
wire		M_162 ;
wire		M_161 ;
wire		M_160 ;
wire		M_159 ;
wire		M_158 ;
wire		M_157 ;
wire		M_156 ;
wire		M_155 ;
wire		M_154 ;
wire		M_153 ;
wire		M_152 ;
wire		M_151 ;
wire		M_150 ;
wire		M_149 ;
wire		M_148 ;
wire		M_147 ;
wire		M_146 ;
wire		M_145 ;
wire		M_144 ;
wire		M_143 ;
wire		M_142 ;
wire		M_141 ;
wire		M_140 ;
wire		M_139 ;
wire		M_138 ;
wire		M_137 ;
wire		M_136 ;
wire		M_135 ;
wire		M_134 ;
wire		M_133 ;
wire		M_132 ;
wire		M_131 ;
wire		M_130 ;
wire		M_129 ;
wire		M_128 ;
wire		M_127 ;
wire		M_126 ;
wire		M_125 ;
wire		M_124 ;
wire		M_123 ;
wire		M_122 ;
wire		M_120 ;
wire		M_119 ;
wire		M_118 ;
wire		M_117 ;
wire		M_116 ;
wire		M_115 ;
wire		M_114 ;
wire		M_113 ;
wire		M_112 ;
wire		M_110 ;
wire		M_109 ;
wire		M_108 ;
wire		M_107 ;
wire		M_106 ;
wire		M_105 ;
wire		M_104 ;
wire		M_103 ;
wire		M_102 ;
wire		M_100 ;
wire		M_99 ;
wire		M_98 ;
wire		M_97 ;
wire		M_96 ;
wire		M_95 ;
wire		M_94 ;
wire		M_93 ;
wire		M_92 ;
wire		M_91 ;
wire		M_90 ;
wire		M_89 ;
wire		M_88 ;
wire		M_87 ;
wire		M_86 ;
wire		M_85 ;
wire		M_84 ;
wire		M_83 ;
wire		M_82 ;
wire		M_81 ;
wire		M_80 ;
wire		M_79 ;
wire		M_78 ;
wire		M_77 ;
wire		M_76 ;
wire		M_75 ;
wire		M_74 ;
wire		M_73 ;
wire		M_72 ;
wire		M_71 ;
wire		M_70 ;
wire		M_69 ;
wire		M_68 ;
wire		M_67 ;
wire		M_66 ;
wire		M_65 ;
wire		M_64 ;
wire		M_63 ;
wire		M_62 ;
wire		M_61 ;
wire		M_60 ;
wire		M_59 ;
wire		M_58 ;
wire		M_57 ;
wire		M_56 ;
wire		M_55 ;
wire		M_54 ;
wire		M_53 ;
wire		M_52 ;
wire		M_51 ;
wire		M_50 ;
wire		M_49 ;
wire		M_48 ;
wire		M_39 ;
wire		U_318 ;
wire		C_09 ;
wire		U_317 ;
wire		U_184 ;
wire		U_183 ;
wire		C_08 ;
wire		U_174 ;
wire		U_173 ;
wire		U_170 ;
wire		C_07 ;
wire		U_166 ;
wire		U_165 ;
wire		U_164 ;
wire		U_163 ;
wire		U_162 ;
wire		C_05 ;
wire		U_161 ;
wire		U_88 ;
wire		U_87 ;
wire		U_84 ;
wire		U_83 ;
wire		U_82 ;
wire		U_81 ;
wire		U_80 ;
wire		C_02 ;
wire		U_79 ;
wire		U_06 ;
wire		U_05 ;
wire		C_01 ;
wire		U_01 ;
wire	[1:0]	sub8u_7_11i2 ;
wire	[6:0]	sub8u_7_11ot ;
wire	[2:0]	sub8u_71i2 ;
wire	[6:0]	sub8u_71i1 ;
wire	[6:0]	sub8u_71ot ;
wire	[31:0]	decr32s2i1 ;
wire	[31:0]	decr32s2ot ;
wire	[31:0]	decr32s1i1 ;
wire	[31:0]	decr32s1ot ;
wire	[6:0]	decr8u_71i1 ;
wire	[6:0]	decr8u_71ot ;
wire	[31:0]	incr32s2i1 ;
wire	[31:0]	incr32s2ot ;
wire	[31:0]	incr32s1i1 ;
wire	[31:0]	incr32s1ot ;
wire	[7:0]	incr8u4i1 ;
wire	[7:0]	incr8u4ot ;
wire	[7:0]	incr8u3ot ;
wire	[7:0]	incr8u2i1 ;
wire	[7:0]	incr8u2ot ;
wire	[7:0]	incr8u1i1 ;
wire	[7:0]	incr8u1ot ;
wire	[3:0]	incr4s1i1 ;
wire	[3:0]	incr4s1ot ;
wire	[5:0]	lop8u_11i2 ;
wire	[5:0]	lop8u_11i1 ;
wire		lop8u_11ot ;
wire	[8:0]	sub12s_91i2 ;
wire	[8:0]	sub12s_91i1 ;
wire	[8:0]	sub12s_91ot ;
wire	[1:0]	sub8u1i2 ;
wire	[7:0]	sub8u1i1 ;
wire	[7:0]	sub8u1ot ;
wire		JF_06 ;
wire		CT_18 ;
wire		JF_03 ;
wire		CT_03 ;
wire		JF_01 ;
wire		FF_j_en ;
wire		FF_i_en ;
wire		jpeg_out_a00_r_en ;
wire		jpeg_out_a01_r_en ;
wire		jpeg_out_a02_r_en ;
wire		jpeg_out_a03_r_en ;
wire		jpeg_out_a04_r_en ;
wire		jpeg_out_a05_r_en ;
wire		jpeg_out_a06_r_en ;
wire		jpeg_out_a07_r_en ;
wire		jpeg_out_a08_r_en ;
wire		jpeg_out_a09_r_en ;
wire		jpeg_out_a10_r_en ;
wire		jpeg_out_a11_r_en ;
wire		jpeg_out_a12_r_en ;
wire		jpeg_out_a13_r_en ;
wire		jpeg_out_a14_r_en ;
wire		jpeg_out_a15_r_en ;
wire		jpeg_out_a16_r_en ;
wire		jpeg_out_a17_r_en ;
wire		jpeg_out_a18_r_en ;
wire		jpeg_out_a19_r_en ;
wire		jpeg_out_a20_r_en ;
wire		jpeg_out_a21_r_en ;
wire		jpeg_out_a22_r_en ;
wire		jpeg_out_a23_r_en ;
wire		jpeg_out_a24_r_en ;
wire		jpeg_out_a25_r_en ;
wire		jpeg_out_a26_r_en ;
wire		jpeg_out_a27_r_en ;
wire		jpeg_out_a28_r_en ;
wire		jpeg_out_a29_r_en ;
wire		jpeg_out_a30_r_en ;
wire		jpeg_out_a31_r_en ;
wire		jpeg_out_a32_r_en ;
wire		jpeg_out_a33_r_en ;
wire		jpeg_out_a34_r_en ;
wire		jpeg_out_a35_r_en ;
wire		jpeg_out_a36_r_en ;
wire		jpeg_out_a37_r_en ;
wire		jpeg_out_a38_r_en ;
wire		jpeg_out_a39_r_en ;
wire		jpeg_out_a40_r_en ;
wire		jpeg_out_a41_r_en ;
wire		jpeg_out_a42_r_en ;
wire		jpeg_out_a43_r_en ;
wire		jpeg_out_a44_r_en ;
wire		jpeg_out_a45_r_en ;
wire		jpeg_out_a46_r_en ;
wire		jpeg_out_a47_r_en ;
wire		jpeg_out_a48_r_en ;
wire		jpeg_out_a49_r_en ;
wire		jpeg_out_a50_r_en ;
wire		jpeg_out_a51_r_en ;
wire		jpeg_out_a52_r_en ;
wire		jpeg_out_a53_r_en ;
wire		jpeg_out_a54_r_en ;
wire		jpeg_out_a55_r_en ;
wire		jpeg_out_a56_r_en ;
wire		jpeg_out_a57_r_en ;
wire		jpeg_out_a58_r_en ;
wire		jpeg_out_a59_r_en ;
wire		jpeg_out_a60_r_en ;
wire		jpeg_out_a61_r_en ;
wire		jpeg_out_a62_r_en ;
wire		jpeg_out_a63_r_en ;
wire		jpeg_out_a64_r_en ;
wire		jpeg_out_a65_r_en ;
wire		jpeg_out_a66_r_en ;
wire		jpeg_out_a67_r_en ;
wire		jpeg_out_a68_r_en ;
wire		jpeg_out_a69_r_en ;
wire		jpeg_out_a70_r_en ;
wire		jpeg_out_a71_r_en ;
wire		jpeg_out_a72_r_en ;
wire		jpeg_out_a73_r_en ;
wire		jpeg_out_a74_r_en ;
wire		jpeg_out_a75_r_en ;
wire		jpeg_out_a76_r_en ;
wire		jpeg_out_a77_r_en ;
wire		jpeg_out_a78_r_en ;
wire		jpeg_out_a79_r_en ;
wire		jpeg_out_a80_r_en ;
wire		jpeg_out_a81_r_en ;
wire		jpeg_out_a82_r_en ;
wire		jpeg_out_a83_r_en ;
wire		jpeg_out_a84_r_en ;
wire		jpeg_out_a85_r_en ;
wire		jpeg_out_a86_r_en ;
wire		jpeg_out_a87_r_en ;
wire		jpeg_out_a88_r_en ;
wire		jpeg_out_a89_r_en ;
wire		jpeg_out_a90_r_en ;
wire		jpeg_out_a91_r_en ;
wire		jpeg_out_a92_r_en ;
wire		jpeg_out_a93_r_en ;
wire		jpeg_out_a94_r_en ;
wire		jpeg_out_a95_r_en ;
wire		jpeg_out_a96_r_en ;
wire		jpeg_out_a97_r_en ;
wire		jpeg_out_a98_r_en ;
wire		jpeg_out_a99_r_en ;
wire		jpeg_out_a100_r_en ;
wire		jpeg_out_a101_r_en ;
wire		jpeg_out_a102_r_en ;
wire		jpeg_out_a103_r_en ;
wire		jpeg_out_a104_r_en ;
wire		jpeg_out_a105_r_en ;
wire		jpeg_out_a106_r_en ;
wire		jpeg_out_a107_r_en ;
wire		jpeg_out_a108_r_en ;
wire		jpeg_out_a109_r_en ;
wire		jpeg_out_a110_r_en ;
wire		jpeg_out_a111_r_en ;
wire		jpeg_out_a112_r_en ;
wire		jpeg_out_a113_r_en ;
wire		jpeg_out_a114_r_en ;
wire		jpeg_out_a115_r_en ;
wire		jpeg_out_a116_r_en ;
wire		jpeg_out_a117_r_en ;
wire		jpeg_out_a118_r_en ;
wire		jpeg_out_a119_r_en ;
wire		jpeg_out_a120_r_en ;
wire		jpeg_out_a121_r_en ;
wire		jpeg_out_a122_r_en ;
wire		jpeg_out_a123_r_en ;
wire		jpeg_out_a124_r_en ;
wire		jpeg_out_a125_r_en ;
wire		jpeg_out_a126_r_en ;
wire		jpeg_out_a127_r_en ;
wire		jpeg_len_out_r_en ;
wire		RG_rl_en ;
wire		RG_previous_dc_zz_en ;
wire		RG_rl_1_en ;
wire		RG_rl_2_en ;
wire		RG_rl_3_en ;
wire		RG_rl_4_en ;
wire		RG_rl_5_en ;
wire		RG_rl_6_en ;
wire		RG_rl_7_en ;
wire		RG_rl_8_en ;
wire		RG_rl_9_en ;
wire		RG_rl_10_en ;
wire		RG_rl_11_en ;
wire		RG_rl_12_en ;
wire		RG_rl_13_en ;
wire		RG_rl_14_en ;
wire		RG_rl_15_en ;
wire		RG_rl_16_en ;
wire		RG_rl_17_en ;
wire		RG_rl_18_en ;
wire		RG_rl_19_en ;
wire		RG_rl_20_en ;
wire		RG_rl_21_en ;
wire		RG_rl_22_en ;
wire		RG_rl_23_en ;
wire		RG_rl_24_en ;
wire		RG_rl_25_en ;
wire		RG_rl_26_en ;
wire		RG_rl_27_en ;
wire		RG_rl_28_en ;
wire		RG_rl_29_en ;
wire		RG_rl_30_en ;
wire		RG_rl_31_en ;
wire		RG_rl_32_en ;
wire		RG_rl_33_en ;
wire		RG_rl_34_en ;
wire		RG_rl_35_en ;
wire		RG_rl_36_en ;
wire		RG_rl_37_en ;
wire		RG_rl_38_en ;
wire		RG_rl_39_en ;
wire		RG_rl_40_en ;
wire		RG_rl_41_en ;
wire		RG_rl_42_en ;
wire		RG_rl_43_en ;
wire		RG_rl_44_en ;
wire		RG_rl_45_en ;
wire		RG_rl_46_en ;
wire		RG_rl_47_en ;
wire		RG_rl_48_en ;
wire		RG_rl_49_en ;
wire		RG_rl_50_en ;
wire		RG_rl_51_en ;
wire		RG_rl_52_en ;
wire		RG_rl_53_en ;
wire		RG_rl_54_en ;
wire		RG_rl_55_en ;
wire		RG_rl_56_en ;
wire		RG_rl_57_en ;
wire		RG_rl_58_en ;
wire		RG_rl_59_en ;
wire		RG_rl_60_en ;
wire		RG_rl_61_en ;
wire		RG_rl_62_en ;
wire		RG_rl_63_en ;
wire		RG_rl_64_en ;
wire		RG_rl_65_en ;
wire		RG_rl_66_en ;
wire		RG_rl_67_en ;
wire		RG_rl_68_en ;
wire		RG_rl_69_en ;
wire		RG_rl_70_en ;
wire		RG_rl_71_en ;
wire		RG_rl_72_en ;
wire		RG_rl_73_en ;
wire		RG_rl_74_en ;
wire		RG_rl_75_en ;
wire		RG_rl_76_en ;
wire		RG_rl_77_en ;
wire		RG_rl_78_en ;
wire		RG_rl_79_en ;
wire		RG_rl_80_en ;
wire		RG_rl_81_en ;
wire		RG_rl_82_en ;
wire		RG_rl_83_en ;
wire		RG_rl_84_en ;
wire		RG_rl_85_en ;
wire		RG_rl_86_en ;
wire		RG_rl_87_en ;
wire		RG_rl_88_en ;
wire		RG_rl_89_en ;
wire		RG_rl_90_en ;
wire		RG_rl_91_en ;
wire		RG_rl_92_en ;
wire		RG_rl_93_en ;
wire		RG_rl_94_en ;
wire		RG_rl_95_en ;
wire		RG_rl_96_en ;
wire		RG_rl_97_en ;
wire		RG_rl_98_en ;
wire		RG_rl_99_en ;
wire		RG_rl_100_en ;
wire		RG_rl_101_en ;
wire		RG_rl_102_en ;
wire		RG_rl_103_en ;
wire		RG_rl_104_en ;
wire		RG_rl_105_en ;
wire		RG_rl_106_en ;
wire		RG_rl_107_en ;
wire		RG_rl_108_en ;
wire		RG_rl_109_en ;
wire		RG_rl_110_en ;
wire		RG_rl_111_en ;
wire		RG_rl_112_en ;
wire		RG_rl_113_en ;
wire		RG_rl_114_en ;
wire		RG_rl_115_en ;
wire		RG_rl_116_en ;
wire		RG_rl_117_en ;
wire		RG_rl_118_en ;
wire		RG_rl_119_en ;
wire		RG_rl_120_en ;
wire		RG_rl_121_en ;
wire		RG_rl_122_en ;
wire		RG_rl_123_en ;
wire		RG_rl_124_en ;
wire		RG_rl_125_en ;
wire		RG_rl_126_en ;
wire		RG_rl_127_en ;
wire		RG_zz_en ;
wire		RG_zz_1_en ;
wire		RG_zz_2_en ;
wire		RG_zz_3_en ;
wire		RG_zz_4_en ;
wire		RG_zz_5_en ;
wire		RG_zz_6_en ;
wire		RG_zz_7_en ;
wire		RG_zz_8_en ;
wire		RG_zz_9_en ;
wire		RG_zz_10_en ;
wire		RG_zz_11_en ;
wire		RG_zz_12_en ;
wire		RG_zz_13_en ;
wire		RG_zz_14_en ;
wire		RG_zz_15_en ;
wire		RG_zz_16_en ;
wire		RG_zz_17_en ;
wire		RG_zz_18_en ;
wire		RG_zz_19_en ;
wire		RG_zz_20_en ;
wire		RG_zz_21_en ;
wire		RG_zz_22_en ;
wire		RG_zz_23_en ;
wire		RG_zz_24_en ;
wire		RG_zz_25_en ;
wire		RG_zz_26_en ;
wire		RG_zz_27_en ;
wire		RG_zz_28_en ;
wire		RG_zz_29_en ;
wire		RG_zz_30_en ;
wire		RG_zz_31_en ;
wire		RG_zz_32_en ;
wire		RG_zz_33_en ;
wire		RG_zz_34_en ;
wire		RG_zz_35_en ;
wire		RG_zz_36_en ;
wire		RG_zz_37_en ;
wire		RG_zz_38_en ;
wire		RG_zz_39_en ;
wire		RG_zz_40_en ;
wire		RG_zz_41_en ;
wire		RG_zz_42_en ;
wire		RG_zz_43_en ;
wire		RG_zz_44_en ;
wire		RG_zz_45_en ;
wire		RG_zz_46_en ;
wire		RG_zz_47_en ;
wire		RG_zz_48_en ;
wire		RG_zz_49_en ;
wire		RG_zz_50_en ;
wire		RG_zz_51_en ;
wire		RG_zz_52_en ;
wire		RG_zz_53_en ;
wire		RG_zz_54_en ;
wire		RG_zz_55_en ;
wire		RG_zz_56_en ;
wire		RG_zz_57_en ;
wire		RG_zz_58_en ;
wire		RG_zz_59_en ;
wire		RG_zz_60_en ;
wire		RG_zz_61_en ;
wire		RG_zz_62_en ;
wire		RG_i_k_01_en ;
wire		RG_i_j_01_en ;
wire		RG_quantized_block_rl_en ;
wire		RG_quantized_block_rl_1_en ;
wire		RG_quantized_block_rl_2_en ;
wire		RG_quantized_block_rl_3_en ;
wire		RG_quantized_block_rl_4_en ;
wire		RG_quantized_block_rl_5_en ;
wire		RG_quantized_block_rl_6_en ;
wire		RG_quantized_block_rl_7_en ;
wire		RG_quantized_block_rl_8_en ;
wire		RG_quantized_block_rl_9_en ;
wire		RG_quantized_block_rl_10_en ;
wire		RG_quantized_block_rl_11_en ;
wire		RG_quantized_block_rl_12_en ;
wire		RG_quantized_block_rl_13_en ;
wire		RG_quantized_block_rl_14_en ;
wire		RG_quantized_block_rl_15_en ;
wire		RG_quantized_block_rl_16_en ;
wire		RG_quantized_block_rl_17_en ;
wire		RG_quantized_block_rl_18_en ;
wire		RG_quantized_block_rl_19_en ;
wire		RG_quantized_block_rl_20_en ;
wire		RG_quantized_block_rl_21_en ;
wire		RG_quantized_block_rl_22_en ;
wire		RG_quantized_block_rl_23_en ;
wire		RG_quantized_block_rl_24_en ;
wire		RG_quantized_block_rl_25_en ;
wire		RG_quantized_block_rl_26_en ;
wire		RG_quantized_block_rl_27_en ;
wire		RG_quantized_block_rl_28_en ;
wire		RG_quantized_block_rl_29_en ;
wire		RG_quantized_block_rl_30_en ;
wire		RG_quantized_block_rl_31_en ;
wire		RG_quantized_block_rl_32_en ;
wire		RG_quantized_block_rl_33_en ;
wire		RG_quantized_block_rl_34_en ;
wire		RG_quantized_block_rl_35_en ;
wire		RG_quantized_block_rl_36_en ;
wire		RG_quantized_block_rl_37_en ;
wire		RG_quantized_block_rl_38_en ;
wire		RG_quantized_block_rl_39_en ;
wire		RG_quantized_block_rl_40_en ;
wire		RG_quantized_block_rl_41_en ;
wire		RG_quantized_block_rl_42_en ;
wire		RG_quantized_block_rl_43_en ;
wire		RG_quantized_block_rl_44_en ;
wire		RG_quantized_block_rl_45_en ;
wire		RG_quantized_block_rl_46_en ;
wire		RG_quantized_block_rl_47_en ;
wire		RG_quantized_block_rl_48_en ;
wire		RG_quantized_block_rl_49_en ;
wire		RG_quantized_block_rl_50_en ;
wire		RG_quantized_block_rl_51_en ;
wire		RG_quantized_block_rl_52_en ;
wire		RG_quantized_block_rl_53_en ;
wire		RG_quantized_block_rl_54_en ;
wire		RG_quantized_block_rl_55_en ;
wire		RG_quantized_block_rl_56_en ;
wire		RG_quantized_block_rl_57_en ;
wire		RG_quantized_block_rl_58_en ;
wire		RG_quantized_block_rl_59_en ;
wire		RG_quantized_block_rl_60_en ;
wire		RG_quantized_block_rl_61_en ;
wire		RG_k_quantized_block_rl_01_en ;
wire		RG_quantized_block_rl_zz_en ;
wire		FF_d_en ;
wire		RG_previous_dc_rl_en ;
wire		RG_rl_128_en ;
wire		RG_rl_129_en ;
wire		RG_rl_130_en ;
wire		RG_rl_131_en ;
wire		RG_rl_132_en ;
wire		RG_rl_133_en ;
wire		RG_rl_134_en ;
wire		RG_rl_135_en ;
wire		RG_rl_136_en ;
wire		RG_rl_137_en ;
wire		RG_rl_138_en ;
wire		RG_rl_139_en ;
wire		RG_rl_140_en ;
wire		RG_rl_141_en ;
wire		RG_rl_142_en ;
wire		RG_rl_143_en ;
wire		RG_rl_144_en ;
wire		RG_rl_145_en ;
wire		RG_rl_146_en ;
wire		RG_rl_147_en ;
wire		RG_rl_148_en ;
wire		RG_rl_149_en ;
wire		RG_rl_150_en ;
wire		RG_rl_151_en ;
wire		RG_rl_152_en ;
wire		RG_rl_153_en ;
wire		RG_rl_154_en ;
wire		RG_rl_155_en ;
wire		RG_rl_156_en ;
wire		RG_rl_157_en ;
wire		RG_rl_158_en ;
wire		RG_rl_159_en ;
wire		RG_rl_160_en ;
wire		RG_rl_161_en ;
wire		RG_rl_162_en ;
wire		RG_rl_163_en ;
wire		RG_rl_164_en ;
wire		RG_rl_165_en ;
wire		RG_rl_166_en ;
wire		RG_rl_167_en ;
wire		RG_rl_168_en ;
wire		RG_rl_169_en ;
wire		RG_rl_170_en ;
wire		RG_rl_171_en ;
wire		RG_rl_172_en ;
wire		RG_rl_173_en ;
wire		RG_rl_174_en ;
wire		RG_rl_175_en ;
wire		RG_rl_176_en ;
wire		RG_rl_177_en ;
wire		RG_rl_178_en ;
wire		RG_rl_179_en ;
wire		RG_rl_180_en ;
wire		RG_rl_181_en ;
wire		RG_rl_182_en ;
wire		RG_rl_183_en ;
wire		RG_rl_184_en ;
wire		RG_rl_185_en ;
wire		RG_rl_186_en ;
wire		RG_rl_187_en ;
wire		RG_rl_188_en ;
wire		RG_rl_189_en ;
wire		RG_rl_190_en ;
wire		RG_rl_191_en ;
wire		RG_len_en ;
wire		valid_r_en ;
reg	[8:0]	RG_rl ;	// line#=../rle.cpp:23
reg	[8:0]	RG_previous_dc_zz ;	// line#=../rle.h:65,66
reg	[8:0]	RG_rl_1 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_2 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_3 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_4 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_5 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_6 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_7 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_8 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_9 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_10 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_11 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_12 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_13 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_14 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_15 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_16 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_17 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_18 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_19 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_20 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_21 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_22 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_23 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_24 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_25 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_26 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_27 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_28 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_29 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_30 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_31 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_32 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_33 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_34 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_35 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_36 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_37 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_38 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_39 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_40 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_41 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_42 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_43 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_44 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_45 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_46 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_47 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_48 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_49 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_50 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_51 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_52 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_53 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_54 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_55 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_56 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_57 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_58 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_59 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_60 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_61 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_62 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_63 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_64 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_65 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_66 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_67 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_68 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_69 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_70 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_71 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_72 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_73 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_74 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_75 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_76 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_77 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_78 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_79 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_80 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_81 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_82 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_83 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_84 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_85 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_86 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_87 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_88 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_89 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_90 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_91 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_92 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_93 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_94 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_95 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_96 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_97 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_98 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_99 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_100 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_101 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_102 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_103 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_104 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_105 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_106 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_107 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_108 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_109 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_110 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_111 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_112 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_113 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_114 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_115 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_116 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_117 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_118 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_119 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_120 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_121 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_122 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_123 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_124 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_125 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_126 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_127 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_zz ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_1 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_2 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_3 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_4 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_5 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_6 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_7 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_8 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_9 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_10 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_11 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_12 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_13 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_14 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_15 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_16 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_17 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_18 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_19 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_20 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_21 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_22 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_23 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_24 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_25 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_26 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_27 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_28 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_29 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_30 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_31 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_32 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_33 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_34 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_35 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_36 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_37 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_38 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_39 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_40 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_41 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_42 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_43 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_44 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_45 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_46 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_47 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_48 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_49 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_50 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_51 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_52 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_53 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_54 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_55 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_56 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_57 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_58 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_59 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_60 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_61 ;	// line#=../rle.h:65
reg	[8:0]	RG_zz_62 ;	// line#=../rle.h:65
reg	[3:0]	RG_j ;	// line#=../rle.cpp:27
reg	[31:0]	RG_i_k_01 ;	// line#=../rle.cpp:25,105
reg	[31:0]	RG_i_j_01 ;	// line#=../rle.cpp:25,105
reg	[8:0]	RG_quantized_block_rl ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_1 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_2 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_3 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_4 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_5 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_6 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_7 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_8 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_9 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_10 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_11 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_12 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_13 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_14 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_15 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_16 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_17 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_18 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_19 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_20 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_21 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_22 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_23 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_24 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_25 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_26 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_27 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_28 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_29 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_30 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_31 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_32 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_33 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_34 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_35 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_36 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_37 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_38 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_39 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_40 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_41 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_42 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_43 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_44 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_45 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_46 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_47 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_48 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_49 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_50 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_51 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_52 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_53 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_54 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_55 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_56 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_57 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_58 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_59 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_60 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_61 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:22,23,25
reg	[8:0]	RG_quantized_block_rl_zz ;	// line#=../rle.cpp:22,23 ../rle.h:65
reg	[5:0]	RG_k ;	// line#=../rle.cpp:105
reg	FF_d ;	// line#=../rle.cpp:105
reg	FF_j ;	// line#=../rle.cpp:27
reg	FF_i ;	// line#=../rle.cpp:24,25
reg	[8:0]	RG_previous_dc_rl ;	// line#=../rle.h:66 ../rle.cpp:23
reg	[8:0]	RG_rl_128 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_129 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_130 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_131 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_132 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_133 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_134 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_135 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_136 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_137 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_138 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_139 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_140 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_141 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_142 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_143 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_144 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_145 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_146 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_147 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_148 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_149 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_150 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_151 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_152 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_153 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_154 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_155 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_156 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_157 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_158 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_159 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_160 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_161 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_162 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_163 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_164 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_165 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_166 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_167 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_168 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_169 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_170 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_171 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_172 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_173 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_174 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_175 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_176 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_177 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_178 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_179 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_180 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_181 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_182 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_183 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_184 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_185 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_186 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_187 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_188 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_189 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_190 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_191 ;	// line#=../rle.cpp:23
reg	[7:0]	RG_len ;	// line#=../rle.cpp:24
reg	[7:0]	RG_len_1 ;	// line#=../rle.cpp:24
reg	[6:0]	RG_k_1 ;	// line#=../rle.cpp:105
reg	[8:0]	jpeg_out_a00_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a01_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a02_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a03_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a04_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a05_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a06_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a07_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a08_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a09_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a10_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a11_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a12_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a13_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a14_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a15_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a16_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a17_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a18_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a19_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a20_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a21_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a22_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a23_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a24_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a25_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a26_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a27_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a28_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a29_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a30_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a31_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a32_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a33_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a34_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a35_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a36_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a37_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a38_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a39_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a40_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a41_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a42_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a43_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a44_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a45_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a46_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a47_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a48_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a49_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a50_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a51_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a52_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a53_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a54_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a55_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a56_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a57_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a58_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a59_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a60_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a61_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a62_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a63_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a64_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a65_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a66_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a67_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a68_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a69_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a70_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a71_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a72_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a73_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a74_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a75_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a76_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a77_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a78_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a79_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a80_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a81_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a82_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a83_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a84_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a85_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a86_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a87_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a88_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a89_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a90_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a91_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a92_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a93_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a94_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a95_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a96_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a97_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a98_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a99_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a100_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a101_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a102_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a103_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a104_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a105_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a106_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a107_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a108_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a109_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a110_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a111_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a112_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a113_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a114_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a115_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a116_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a117_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a118_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a119_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a120_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a121_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a122_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a123_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a124_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a125_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a126_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a127_r ;	// line#=../rle.h:60
reg	[11:0]	jpeg_len_out_r ;	// line#=../rle.h:61
reg	valid_r ;	// line#=../rle.h:62
reg	M_14_t128 ;
reg	[8:0]	TR_12 ;
reg	[8:0]	TR_13 ;
reg	[8:0]	TR_14 ;
reg	[8:0]	TR_15 ;
reg	[8:0]	TR_16 ;
reg	[8:0]	TR_17 ;
reg	[8:0]	TR_18 ;
reg	[8:0]	TR_19 ;
reg	[8:0]	TR_20 ;
reg	[8:0]	TR_21 ;
reg	[8:0]	TR_22 ;
reg	[8:0]	TR_23 ;
reg	[8:0]	TR_24 ;
reg	[8:0]	TR_25 ;
reg	[8:0]	TR_26 ;
reg	[8:0]	TR_27 ;
reg	[8:0]	TR_28 ;
reg	[8:0]	TR_29 ;
reg	[8:0]	TR_30 ;
reg	[8:0]	TR_31 ;
reg	[8:0]	TR_32 ;
reg	[8:0]	TR_33 ;
reg	[8:0]	TR_34 ;
reg	[8:0]	TR_35 ;
reg	[8:0]	TR_36 ;
reg	[8:0]	TR_37 ;
reg	[8:0]	TR_38 ;
reg	[8:0]	TR_39 ;
reg	[8:0]	TR_40 ;
reg	[8:0]	TR_41 ;
reg	[8:0]	TR_42 ;
reg	[8:0]	TR_43 ;
reg	[8:0]	TR_44 ;
reg	[8:0]	TR_45 ;
reg	[8:0]	TR_46 ;
reg	[8:0]	TR_47 ;
reg	[8:0]	TR_48 ;
reg	[8:0]	TR_49 ;
reg	[8:0]	TR_50 ;
reg	[8:0]	TR_51 ;
reg	[8:0]	TR_52 ;
reg	[8:0]	TR_53 ;
reg	[8:0]	TR_54 ;
reg	[8:0]	TR_55 ;
reg	[8:0]	TR_56 ;
reg	[8:0]	TR_57 ;
reg	[8:0]	TR_58 ;
reg	[8:0]	TR_59 ;
reg	[8:0]	TR_60 ;
reg	[8:0]	TR_61 ;
reg	[8:0]	TR_62 ;
reg	[8:0]	TR_63 ;
reg	[8:0]	TR_64 ;
reg	[8:0]	TR_65 ;
reg	[8:0]	TR_66 ;
reg	[8:0]	TR_67 ;
reg	[8:0]	TR_68 ;
reg	[8:0]	TR_69 ;
reg	[8:0]	TR_70 ;
reg	[8:0]	TR_71 ;
reg	[8:0]	TR_72 ;
reg	[8:0]	TR_73 ;
reg	[8:0]	TR_74 ;
reg	[8:0]	TR_75 ;
reg	[8:0]	TR_76 ;
reg	[8:0]	TR_77 ;
reg	[8:0]	TR_78 ;
reg	[8:0]	TR_79 ;
reg	[8:0]	TR_80 ;
reg	[8:0]	TR_81 ;
reg	[8:0]	TR_82 ;
reg	[8:0]	TR_83 ;
reg	[8:0]	TR_84 ;
reg	[8:0]	TR_85 ;
reg	[8:0]	TR_86 ;
reg	[8:0]	TR_87 ;
reg	[8:0]	TR_88 ;
reg	[8:0]	TR_89 ;
reg	[8:0]	TR_90 ;
reg	[8:0]	TR_91 ;
reg	[8:0]	TR_92 ;
reg	[8:0]	TR_93 ;
reg	[8:0]	TR_94 ;
reg	[8:0]	TR_95 ;
reg	[8:0]	TR_96 ;
reg	[8:0]	TR_97 ;
reg	[8:0]	TR_98 ;
reg	[8:0]	TR_99 ;
reg	[8:0]	TR_100 ;
reg	[8:0]	TR_101 ;
reg	[8:0]	TR_102 ;
reg	[8:0]	TR_103 ;
reg	[8:0]	TR_104 ;
reg	[8:0]	TR_105 ;
reg	[8:0]	TR_106 ;
reg	[8:0]	TR_107 ;
reg	[8:0]	TR_108 ;
reg	[8:0]	TR_109 ;
reg	[8:0]	TR_110 ;
reg	[8:0]	TR_111 ;
reg	[8:0]	TR_112 ;
reg	[8:0]	TR_113 ;
reg	[8:0]	TR_114 ;
reg	[8:0]	TR_115 ;
reg	[8:0]	TR_116 ;
reg	[8:0]	TR_117 ;
reg	[8:0]	TR_118 ;
reg	[8:0]	TR_119 ;
reg	[8:0]	TR_120 ;
reg	[8:0]	TR_121 ;
reg	[8:0]	TR_122 ;
reg	[8:0]	TR_123 ;
reg	[8:0]	TR_124 ;
reg	[8:0]	TR_125 ;
reg	[8:0]	TR_126 ;
reg	[8:0]	TR_127 ;
reg	[8:0]	TR_128 ;
reg	[8:0]	TR_129 ;
reg	[8:0]	TR_130 ;
reg	[8:0]	TR_131 ;
reg	[8:0]	TR_132 ;
reg	[8:0]	TR_133 ;
reg	[8:0]	TR_134 ;
reg	[8:0]	TR_135 ;
reg	[8:0]	TR_136 ;
reg	[8:0]	TR_137 ;
reg	[8:0]	TR_138 ;
reg	[8:0]	rl_a127_t2 ;
reg	M_15_t128 ;
reg	[8:0]	M_16_t ;
reg	[8:0]	rl_a00_t8 ;
reg	[8:0]	rl_a01_t8 ;
reg	[8:0]	rl_a02_t8 ;
reg	[8:0]	rl_a03_t8 ;
reg	[8:0]	rl_a04_t8 ;
reg	[8:0]	rl_a05_t8 ;
reg	[8:0]	rl_a06_t8 ;
reg	[8:0]	rl_a07_t8 ;
reg	[8:0]	rl_a08_t8 ;
reg	[8:0]	rl_a09_t8 ;
reg	[8:0]	rl_a10_t8 ;
reg	[8:0]	rl_a11_t8 ;
reg	[8:0]	rl_a12_t8 ;
reg	[8:0]	rl_a13_t8 ;
reg	[8:0]	rl_a14_t8 ;
reg	[8:0]	rl_a15_t8 ;
reg	[8:0]	rl_a16_t8 ;
reg	[8:0]	rl_a17_t8 ;
reg	[8:0]	rl_a18_t8 ;
reg	[8:0]	rl_a19_t8 ;
reg	[8:0]	rl_a20_t8 ;
reg	[8:0]	rl_a21_t8 ;
reg	[8:0]	rl_a22_t8 ;
reg	[8:0]	rl_a23_t8 ;
reg	[8:0]	rl_a24_t8 ;
reg	[8:0]	rl_a25_t8 ;
reg	[8:0]	rl_a26_t8 ;
reg	[8:0]	rl_a27_t8 ;
reg	[8:0]	rl_a28_t8 ;
reg	[8:0]	rl_a29_t8 ;
reg	[8:0]	rl_a30_t8 ;
reg	[8:0]	rl_a31_t8 ;
reg	[8:0]	rl_a32_t8 ;
reg	[8:0]	rl_a33_t8 ;
reg	[8:0]	rl_a34_t8 ;
reg	[8:0]	rl_a35_t8 ;
reg	[8:0]	rl_a36_t8 ;
reg	[8:0]	rl_a37_t8 ;
reg	[8:0]	rl_a38_t8 ;
reg	[8:0]	rl_a39_t8 ;
reg	[8:0]	rl_a40_t8 ;
reg	[8:0]	rl_a41_t8 ;
reg	[8:0]	rl_a42_t8 ;
reg	[8:0]	rl_a43_t8 ;
reg	[8:0]	rl_a44_t8 ;
reg	[8:0]	rl_a45_t8 ;
reg	[8:0]	rl_a46_t8 ;
reg	[8:0]	rl_a47_t8 ;
reg	[8:0]	rl_a48_t8 ;
reg	[8:0]	rl_a49_t8 ;
reg	[8:0]	rl_a50_t8 ;
reg	[8:0]	rl_a51_t8 ;
reg	[8:0]	rl_a52_t8 ;
reg	[8:0]	rl_a53_t8 ;
reg	[8:0]	rl_a54_t8 ;
reg	[8:0]	rl_a55_t8 ;
reg	[8:0]	rl_a56_t8 ;
reg	[8:0]	rl_a57_t8 ;
reg	[8:0]	rl_a58_t8 ;
reg	[8:0]	rl_a59_t8 ;
reg	[8:0]	rl_a60_t8 ;
reg	[8:0]	rl_a61_t8 ;
reg	[8:0]	rl_a62_t8 ;
reg	[8:0]	rl_a63_t8 ;
reg	[8:0]	rl_a64_t8 ;
reg	[8:0]	rl_a65_t8 ;
reg	[8:0]	rl_a66_t8 ;
reg	[8:0]	rl_a67_t8 ;
reg	[8:0]	rl_a68_t8 ;
reg	[8:0]	rl_a69_t8 ;
reg	[8:0]	rl_a70_t8 ;
reg	[8:0]	rl_a71_t8 ;
reg	[8:0]	rl_a72_t8 ;
reg	[8:0]	rl_a73_t8 ;
reg	[8:0]	rl_a74_t8 ;
reg	[8:0]	rl_a75_t8 ;
reg	[8:0]	rl_a76_t8 ;
reg	[8:0]	rl_a77_t8 ;
reg	[8:0]	rl_a78_t8 ;
reg	[8:0]	rl_a79_t8 ;
reg	[8:0]	rl_a80_t8 ;
reg	[8:0]	rl_a81_t8 ;
reg	[8:0]	rl_a82_t8 ;
reg	[8:0]	rl_a83_t8 ;
reg	[8:0]	rl_a84_t8 ;
reg	[8:0]	rl_a85_t8 ;
reg	[8:0]	rl_a86_t8 ;
reg	[8:0]	rl_a87_t8 ;
reg	[8:0]	rl_a88_t8 ;
reg	[8:0]	rl_a89_t8 ;
reg	[8:0]	rl_a90_t8 ;
reg	[8:0]	rl_a91_t8 ;
reg	[8:0]	rl_a92_t8 ;
reg	[8:0]	rl_a93_t8 ;
reg	[8:0]	rl_a94_t8 ;
reg	[8:0]	rl_a95_t8 ;
reg	[8:0]	rl_a96_t8 ;
reg	[8:0]	rl_a97_t8 ;
reg	[8:0]	rl_a98_t8 ;
reg	[8:0]	rl_a99_t8 ;
reg	[8:0]	rl_a100_t8 ;
reg	[8:0]	rl_a101_t8 ;
reg	[8:0]	rl_a102_t8 ;
reg	[8:0]	rl_a103_t8 ;
reg	[8:0]	rl_a104_t8 ;
reg	[8:0]	rl_a105_t8 ;
reg	[8:0]	rl_a106_t8 ;
reg	[8:0]	rl_a107_t8 ;
reg	[8:0]	rl_a108_t8 ;
reg	[8:0]	rl_a109_t8 ;
reg	[8:0]	rl_a110_t8 ;
reg	[8:0]	rl_a111_t8 ;
reg	[8:0]	rl_a112_t8 ;
reg	[8:0]	rl_a113_t8 ;
reg	[8:0]	rl_a114_t8 ;
reg	[8:0]	rl_a115_t8 ;
reg	[8:0]	rl_a116_t8 ;
reg	[8:0]	rl_a117_t8 ;
reg	[8:0]	rl_a118_t8 ;
reg	[8:0]	rl_a119_t8 ;
reg	[8:0]	rl_a120_t8 ;
reg	[8:0]	rl_a121_t8 ;
reg	[8:0]	rl_a122_t8 ;
reg	[8:0]	rl_a123_t8 ;
reg	[8:0]	rl_a124_t8 ;
reg	[8:0]	rl_a125_t8 ;
reg	[8:0]	rl_a126_t8 ;
reg	[8:0]	rl_a127_t7 ;
reg	[8:0]	rl_a127_t8 ;
reg	[8:0]	TR_265 ;
reg	[8:0]	RG_rl_t ;
reg	RG_rl_t_c1 ;
reg	[8:0]	RG_previous_dc_zz_t ;
reg	RG_previous_dc_zz_t_c1 ;
reg	RG_previous_dc_zz_t_c2 ;
reg	[8:0]	TR_264 ;
reg	[8:0]	RG_rl_1_t ;
reg	RG_rl_1_t_c1 ;
reg	[8:0]	TR_263 ;
reg	[8:0]	RG_rl_2_t ;
reg	RG_rl_2_t_c1 ;
reg	[8:0]	TR_262 ;
reg	[8:0]	RG_rl_3_t ;
reg	RG_rl_3_t_c1 ;
reg	[8:0]	TR_261 ;
reg	[8:0]	RG_rl_4_t ;
reg	RG_rl_4_t_c1 ;
reg	[8:0]	TR_260 ;
reg	[8:0]	RG_rl_5_t ;
reg	RG_rl_5_t_c1 ;
reg	[8:0]	TR_259 ;
reg	[8:0]	RG_rl_6_t ;
reg	RG_rl_6_t_c1 ;
reg	[8:0]	TR_258 ;
reg	[8:0]	RG_rl_7_t ;
reg	RG_rl_7_t_c1 ;
reg	[8:0]	TR_257 ;
reg	[8:0]	RG_rl_8_t ;
reg	RG_rl_8_t_c1 ;
reg	[8:0]	TR_256 ;
reg	[8:0]	RG_rl_9_t ;
reg	RG_rl_9_t_c1 ;
reg	[8:0]	TR_255 ;
reg	[8:0]	RG_rl_10_t ;
reg	RG_rl_10_t_c1 ;
reg	[8:0]	TR_254 ;
reg	[8:0]	RG_rl_11_t ;
reg	RG_rl_11_t_c1 ;
reg	[8:0]	TR_253 ;
reg	[8:0]	RG_rl_12_t ;
reg	RG_rl_12_t_c1 ;
reg	[8:0]	TR_252 ;
reg	[8:0]	RG_rl_13_t ;
reg	RG_rl_13_t_c1 ;
reg	[8:0]	TR_251 ;
reg	[8:0]	RG_rl_14_t ;
reg	RG_rl_14_t_c1 ;
reg	[8:0]	TR_250 ;
reg	[8:0]	RG_rl_15_t ;
reg	RG_rl_15_t_c1 ;
reg	[8:0]	TR_249 ;
reg	[8:0]	RG_rl_16_t ;
reg	RG_rl_16_t_c1 ;
reg	[8:0]	TR_248 ;
reg	[8:0]	RG_rl_17_t ;
reg	RG_rl_17_t_c1 ;
reg	[8:0]	TR_247 ;
reg	[8:0]	RG_rl_18_t ;
reg	RG_rl_18_t_c1 ;
reg	[8:0]	TR_246 ;
reg	[8:0]	RG_rl_19_t ;
reg	RG_rl_19_t_c1 ;
reg	[8:0]	TR_245 ;
reg	[8:0]	RG_rl_20_t ;
reg	RG_rl_20_t_c1 ;
reg	[8:0]	TR_244 ;
reg	[8:0]	RG_rl_21_t ;
reg	RG_rl_21_t_c1 ;
reg	[8:0]	TR_243 ;
reg	[8:0]	RG_rl_22_t ;
reg	RG_rl_22_t_c1 ;
reg	[8:0]	TR_242 ;
reg	[8:0]	RG_rl_23_t ;
reg	RG_rl_23_t_c1 ;
reg	[8:0]	TR_241 ;
reg	[8:0]	RG_rl_24_t ;
reg	RG_rl_24_t_c1 ;
reg	[8:0]	TR_240 ;
reg	[8:0]	RG_rl_25_t ;
reg	RG_rl_25_t_c1 ;
reg	[8:0]	TR_239 ;
reg	[8:0]	RG_rl_26_t ;
reg	RG_rl_26_t_c1 ;
reg	[8:0]	TR_238 ;
reg	[8:0]	RG_rl_27_t ;
reg	RG_rl_27_t_c1 ;
reg	[8:0]	TR_237 ;
reg	[8:0]	RG_rl_28_t ;
reg	RG_rl_28_t_c1 ;
reg	[8:0]	TR_236 ;
reg	[8:0]	RG_rl_29_t ;
reg	RG_rl_29_t_c1 ;
reg	[8:0]	TR_235 ;
reg	[8:0]	RG_rl_30_t ;
reg	RG_rl_30_t_c1 ;
reg	[8:0]	TR_234 ;
reg	[8:0]	RG_rl_31_t ;
reg	RG_rl_31_t_c1 ;
reg	[8:0]	TR_233 ;
reg	[8:0]	RG_rl_32_t ;
reg	RG_rl_32_t_c1 ;
reg	[8:0]	TR_232 ;
reg	[8:0]	RG_rl_33_t ;
reg	RG_rl_33_t_c1 ;
reg	[8:0]	TR_231 ;
reg	[8:0]	RG_rl_34_t ;
reg	RG_rl_34_t_c1 ;
reg	[8:0]	TR_230 ;
reg	[8:0]	RG_rl_35_t ;
reg	RG_rl_35_t_c1 ;
reg	[8:0]	TR_229 ;
reg	[8:0]	RG_rl_36_t ;
reg	RG_rl_36_t_c1 ;
reg	[8:0]	TR_228 ;
reg	[8:0]	RG_rl_37_t ;
reg	RG_rl_37_t_c1 ;
reg	[8:0]	TR_227 ;
reg	[8:0]	RG_rl_38_t ;
reg	RG_rl_38_t_c1 ;
reg	[8:0]	TR_226 ;
reg	[8:0]	RG_rl_39_t ;
reg	RG_rl_39_t_c1 ;
reg	[8:0]	TR_225 ;
reg	[8:0]	RG_rl_40_t ;
reg	RG_rl_40_t_c1 ;
reg	[8:0]	TR_224 ;
reg	[8:0]	RG_rl_41_t ;
reg	RG_rl_41_t_c1 ;
reg	[8:0]	TR_223 ;
reg	[8:0]	RG_rl_42_t ;
reg	RG_rl_42_t_c1 ;
reg	[8:0]	TR_222 ;
reg	[8:0]	RG_rl_43_t ;
reg	RG_rl_43_t_c1 ;
reg	[8:0]	TR_221 ;
reg	[8:0]	RG_rl_44_t ;
reg	RG_rl_44_t_c1 ;
reg	[8:0]	TR_220 ;
reg	[8:0]	RG_rl_45_t ;
reg	RG_rl_45_t_c1 ;
reg	[8:0]	TR_219 ;
reg	[8:0]	RG_rl_46_t ;
reg	RG_rl_46_t_c1 ;
reg	[8:0]	TR_218 ;
reg	[8:0]	RG_rl_47_t ;
reg	RG_rl_47_t_c1 ;
reg	[8:0]	TR_217 ;
reg	[8:0]	RG_rl_48_t ;
reg	RG_rl_48_t_c1 ;
reg	[8:0]	TR_216 ;
reg	[8:0]	RG_rl_49_t ;
reg	RG_rl_49_t_c1 ;
reg	[8:0]	TR_215 ;
reg	[8:0]	RG_rl_50_t ;
reg	RG_rl_50_t_c1 ;
reg	[8:0]	TR_214 ;
reg	[8:0]	RG_rl_51_t ;
reg	RG_rl_51_t_c1 ;
reg	[8:0]	TR_213 ;
reg	[8:0]	RG_rl_52_t ;
reg	RG_rl_52_t_c1 ;
reg	[8:0]	TR_212 ;
reg	[8:0]	RG_rl_53_t ;
reg	RG_rl_53_t_c1 ;
reg	[8:0]	TR_211 ;
reg	[8:0]	RG_rl_54_t ;
reg	RG_rl_54_t_c1 ;
reg	[8:0]	TR_210 ;
reg	[8:0]	RG_rl_55_t ;
reg	RG_rl_55_t_c1 ;
reg	[8:0]	TR_209 ;
reg	[8:0]	RG_rl_56_t ;
reg	RG_rl_56_t_c1 ;
reg	[8:0]	TR_208 ;
reg	[8:0]	RG_rl_57_t ;
reg	RG_rl_57_t_c1 ;
reg	[8:0]	TR_207 ;
reg	[8:0]	RG_rl_58_t ;
reg	RG_rl_58_t_c1 ;
reg	[8:0]	TR_206 ;
reg	[8:0]	RG_rl_59_t ;
reg	RG_rl_59_t_c1 ;
reg	[8:0]	TR_205 ;
reg	[8:0]	RG_rl_60_t ;
reg	RG_rl_60_t_c1 ;
reg	[8:0]	TR_204 ;
reg	[8:0]	RG_rl_61_t ;
reg	RG_rl_61_t_c1 ;
reg	[8:0]	TR_203 ;
reg	[8:0]	RG_rl_62_t ;
reg	RG_rl_62_t_c1 ;
reg	[8:0]	TR_202 ;
reg	[8:0]	RG_rl_63_t ;
reg	RG_rl_63_t_c1 ;
reg	[8:0]	TR_201 ;
reg	[8:0]	RG_rl_64_t ;
reg	RG_rl_64_t_c1 ;
reg	[8:0]	TR_200 ;
reg	[8:0]	RG_rl_65_t ;
reg	RG_rl_65_t_c1 ;
reg	[8:0]	TR_199 ;
reg	[8:0]	RG_rl_66_t ;
reg	RG_rl_66_t_c1 ;
reg	[8:0]	TR_198 ;
reg	[8:0]	RG_rl_67_t ;
reg	RG_rl_67_t_c1 ;
reg	[8:0]	TR_197 ;
reg	[8:0]	RG_rl_68_t ;
reg	RG_rl_68_t_c1 ;
reg	[8:0]	TR_196 ;
reg	[8:0]	RG_rl_69_t ;
reg	RG_rl_69_t_c1 ;
reg	[8:0]	TR_195 ;
reg	[8:0]	RG_rl_70_t ;
reg	RG_rl_70_t_c1 ;
reg	[8:0]	TR_194 ;
reg	[8:0]	RG_rl_71_t ;
reg	RG_rl_71_t_c1 ;
reg	[8:0]	TR_193 ;
reg	[8:0]	RG_rl_72_t ;
reg	RG_rl_72_t_c1 ;
reg	[8:0]	TR_192 ;
reg	[8:0]	RG_rl_73_t ;
reg	RG_rl_73_t_c1 ;
reg	[8:0]	TR_191 ;
reg	[8:0]	RG_rl_74_t ;
reg	RG_rl_74_t_c1 ;
reg	[8:0]	TR_190 ;
reg	[8:0]	RG_rl_75_t ;
reg	RG_rl_75_t_c1 ;
reg	[8:0]	TR_189 ;
reg	[8:0]	RG_rl_76_t ;
reg	RG_rl_76_t_c1 ;
reg	[8:0]	TR_188 ;
reg	[8:0]	RG_rl_77_t ;
reg	RG_rl_77_t_c1 ;
reg	[8:0]	TR_187 ;
reg	[8:0]	RG_rl_78_t ;
reg	RG_rl_78_t_c1 ;
reg	[8:0]	TR_186 ;
reg	[8:0]	RG_rl_79_t ;
reg	RG_rl_79_t_c1 ;
reg	[8:0]	TR_185 ;
reg	[8:0]	RG_rl_80_t ;
reg	RG_rl_80_t_c1 ;
reg	[8:0]	TR_184 ;
reg	[8:0]	RG_rl_81_t ;
reg	RG_rl_81_t_c1 ;
reg	[8:0]	TR_183 ;
reg	[8:0]	RG_rl_82_t ;
reg	RG_rl_82_t_c1 ;
reg	[8:0]	TR_182 ;
reg	[8:0]	RG_rl_83_t ;
reg	RG_rl_83_t_c1 ;
reg	[8:0]	TR_181 ;
reg	[8:0]	RG_rl_84_t ;
reg	RG_rl_84_t_c1 ;
reg	[8:0]	TR_180 ;
reg	[8:0]	RG_rl_85_t ;
reg	RG_rl_85_t_c1 ;
reg	[8:0]	TR_179 ;
reg	[8:0]	RG_rl_86_t ;
reg	RG_rl_86_t_c1 ;
reg	[8:0]	TR_178 ;
reg	[8:0]	RG_rl_87_t ;
reg	RG_rl_87_t_c1 ;
reg	[8:0]	TR_177 ;
reg	[8:0]	RG_rl_88_t ;
reg	RG_rl_88_t_c1 ;
reg	[8:0]	TR_176 ;
reg	[8:0]	RG_rl_89_t ;
reg	RG_rl_89_t_c1 ;
reg	[8:0]	TR_175 ;
reg	[8:0]	RG_rl_90_t ;
reg	RG_rl_90_t_c1 ;
reg	[8:0]	TR_174 ;
reg	[8:0]	RG_rl_91_t ;
reg	RG_rl_91_t_c1 ;
reg	[8:0]	TR_173 ;
reg	[8:0]	RG_rl_92_t ;
reg	RG_rl_92_t_c1 ;
reg	[8:0]	TR_172 ;
reg	[8:0]	RG_rl_93_t ;
reg	RG_rl_93_t_c1 ;
reg	[8:0]	TR_171 ;
reg	[8:0]	RG_rl_94_t ;
reg	RG_rl_94_t_c1 ;
reg	[8:0]	TR_170 ;
reg	[8:0]	RG_rl_95_t ;
reg	RG_rl_95_t_c1 ;
reg	[8:0]	TR_169 ;
reg	[8:0]	RG_rl_96_t ;
reg	RG_rl_96_t_c1 ;
reg	[8:0]	TR_168 ;
reg	[8:0]	RG_rl_97_t ;
reg	RG_rl_97_t_c1 ;
reg	[8:0]	TR_167 ;
reg	[8:0]	RG_rl_98_t ;
reg	RG_rl_98_t_c1 ;
reg	[8:0]	TR_166 ;
reg	[8:0]	RG_rl_99_t ;
reg	RG_rl_99_t_c1 ;
reg	[8:0]	TR_165 ;
reg	[8:0]	RG_rl_100_t ;
reg	RG_rl_100_t_c1 ;
reg	[8:0]	TR_164 ;
reg	[8:0]	RG_rl_101_t ;
reg	RG_rl_101_t_c1 ;
reg	[8:0]	TR_163 ;
reg	[8:0]	RG_rl_102_t ;
reg	RG_rl_102_t_c1 ;
reg	[8:0]	TR_162 ;
reg	[8:0]	RG_rl_103_t ;
reg	RG_rl_103_t_c1 ;
reg	[8:0]	TR_161 ;
reg	[8:0]	RG_rl_104_t ;
reg	RG_rl_104_t_c1 ;
reg	[8:0]	TR_160 ;
reg	[8:0]	RG_rl_105_t ;
reg	RG_rl_105_t_c1 ;
reg	[8:0]	TR_159 ;
reg	[8:0]	RG_rl_106_t ;
reg	RG_rl_106_t_c1 ;
reg	[8:0]	TR_158 ;
reg	[8:0]	RG_rl_107_t ;
reg	RG_rl_107_t_c1 ;
reg	[8:0]	TR_157 ;
reg	[8:0]	RG_rl_108_t ;
reg	RG_rl_108_t_c1 ;
reg	[8:0]	TR_156 ;
reg	[8:0]	RG_rl_109_t ;
reg	RG_rl_109_t_c1 ;
reg	[8:0]	TR_155 ;
reg	[8:0]	RG_rl_110_t ;
reg	RG_rl_110_t_c1 ;
reg	[8:0]	TR_154 ;
reg	[8:0]	RG_rl_111_t ;
reg	RG_rl_111_t_c1 ;
reg	[8:0]	TR_153 ;
reg	[8:0]	RG_rl_112_t ;
reg	RG_rl_112_t_c1 ;
reg	[8:0]	TR_152 ;
reg	[8:0]	RG_rl_113_t ;
reg	RG_rl_113_t_c1 ;
reg	[8:0]	TR_151 ;
reg	[8:0]	RG_rl_114_t ;
reg	RG_rl_114_t_c1 ;
reg	[8:0]	TR_150 ;
reg	[8:0]	RG_rl_115_t ;
reg	RG_rl_115_t_c1 ;
reg	[8:0]	TR_149 ;
reg	[8:0]	RG_rl_116_t ;
reg	RG_rl_116_t_c1 ;
reg	[8:0]	TR_148 ;
reg	[8:0]	RG_rl_117_t ;
reg	RG_rl_117_t_c1 ;
reg	[8:0]	TR_147 ;
reg	[8:0]	RG_rl_118_t ;
reg	RG_rl_118_t_c1 ;
reg	[8:0]	TR_146 ;
reg	[8:0]	RG_rl_119_t ;
reg	RG_rl_119_t_c1 ;
reg	[8:0]	TR_145 ;
reg	[8:0]	RG_rl_120_t ;
reg	RG_rl_120_t_c1 ;
reg	[8:0]	TR_144 ;
reg	[8:0]	RG_rl_121_t ;
reg	RG_rl_121_t_c1 ;
reg	[8:0]	TR_143 ;
reg	[8:0]	RG_rl_122_t ;
reg	RG_rl_122_t_c1 ;
reg	[8:0]	TR_142 ;
reg	[8:0]	RG_rl_123_t ;
reg	RG_rl_123_t_c1 ;
reg	[8:0]	TR_141 ;
reg	[8:0]	RG_rl_124_t ;
reg	RG_rl_124_t_c1 ;
reg	[8:0]	TR_140 ;
reg	[8:0]	RG_rl_125_t ;
reg	RG_rl_125_t_c1 ;
reg	[8:0]	TR_139 ;
reg	[8:0]	RG_rl_126_t ;
reg	RG_rl_126_t_c1 ;
reg	RG_rl_126_t_c2 ;
reg	[8:0]	RG_rl_127_t ;
reg	RG_rl_127_t_c1 ;
reg	RG_rl_127_t_c2 ;
reg	[8:0]	RG_rl_127_t1 ;
reg	[8:0]	RG_zz_t ;
reg	RG_zz_t_c1 ;
reg	RG_zz_t_c2 ;
reg	[8:0]	RG_zz_1_t ;
reg	RG_zz_1_t_c1 ;
reg	RG_zz_1_t_c2 ;
reg	[8:0]	RG_zz_2_t ;
reg	RG_zz_2_t_c1 ;
reg	RG_zz_2_t_c2 ;
reg	[8:0]	RG_zz_3_t ;
reg	RG_zz_3_t_c1 ;
reg	RG_zz_3_t_c2 ;
reg	[8:0]	RG_zz_4_t ;
reg	RG_zz_4_t_c1 ;
reg	RG_zz_4_t_c2 ;
reg	[8:0]	RG_zz_5_t ;
reg	RG_zz_5_t_c1 ;
reg	RG_zz_5_t_c2 ;
reg	[8:0]	RG_zz_6_t ;
reg	RG_zz_6_t_c1 ;
reg	RG_zz_6_t_c2 ;
reg	[8:0]	RG_zz_7_t ;
reg	RG_zz_7_t_c1 ;
reg	RG_zz_7_t_c2 ;
reg	[8:0]	RG_zz_8_t ;
reg	RG_zz_8_t_c1 ;
reg	RG_zz_8_t_c2 ;
reg	[8:0]	RG_zz_9_t ;
reg	RG_zz_9_t_c1 ;
reg	RG_zz_9_t_c2 ;
reg	[8:0]	RG_zz_10_t ;
reg	RG_zz_10_t_c1 ;
reg	RG_zz_10_t_c2 ;
reg	[8:0]	RG_zz_11_t ;
reg	RG_zz_11_t_c1 ;
reg	RG_zz_11_t_c2 ;
reg	[8:0]	RG_zz_12_t ;
reg	RG_zz_12_t_c1 ;
reg	RG_zz_12_t_c2 ;
reg	[8:0]	RG_zz_13_t ;
reg	RG_zz_13_t_c1 ;
reg	RG_zz_13_t_c2 ;
reg	[8:0]	RG_zz_14_t ;
reg	RG_zz_14_t_c1 ;
reg	RG_zz_14_t_c2 ;
reg	[8:0]	RG_zz_15_t ;
reg	RG_zz_15_t_c1 ;
reg	RG_zz_15_t_c2 ;
reg	[8:0]	RG_zz_16_t ;
reg	RG_zz_16_t_c1 ;
reg	RG_zz_16_t_c2 ;
reg	[8:0]	RG_zz_17_t ;
reg	RG_zz_17_t_c1 ;
reg	RG_zz_17_t_c2 ;
reg	[8:0]	RG_zz_18_t ;
reg	RG_zz_18_t_c1 ;
reg	RG_zz_18_t_c2 ;
reg	[8:0]	RG_zz_19_t ;
reg	RG_zz_19_t_c1 ;
reg	RG_zz_19_t_c2 ;
reg	[8:0]	RG_zz_20_t ;
reg	RG_zz_20_t_c1 ;
reg	RG_zz_20_t_c2 ;
reg	[8:0]	RG_zz_21_t ;
reg	RG_zz_21_t_c1 ;
reg	RG_zz_21_t_c2 ;
reg	[8:0]	RG_zz_22_t ;
reg	RG_zz_22_t_c1 ;
reg	RG_zz_22_t_c2 ;
reg	[8:0]	RG_zz_23_t ;
reg	RG_zz_23_t_c1 ;
reg	RG_zz_23_t_c2 ;
reg	[8:0]	RG_zz_24_t ;
reg	RG_zz_24_t_c1 ;
reg	RG_zz_24_t_c2 ;
reg	[8:0]	RG_zz_25_t ;
reg	RG_zz_25_t_c1 ;
reg	RG_zz_25_t_c2 ;
reg	[8:0]	RG_zz_26_t ;
reg	RG_zz_26_t_c1 ;
reg	RG_zz_26_t_c2 ;
reg	[8:0]	RG_zz_27_t ;
reg	RG_zz_27_t_c1 ;
reg	RG_zz_27_t_c2 ;
reg	[8:0]	RG_zz_28_t ;
reg	RG_zz_28_t_c1 ;
reg	RG_zz_28_t_c2 ;
reg	[8:0]	RG_zz_29_t ;
reg	RG_zz_29_t_c1 ;
reg	RG_zz_29_t_c2 ;
reg	[8:0]	RG_zz_30_t ;
reg	RG_zz_30_t_c1 ;
reg	RG_zz_30_t_c2 ;
reg	[8:0]	RG_zz_31_t ;
reg	RG_zz_31_t_c1 ;
reg	RG_zz_31_t_c2 ;
reg	[8:0]	RG_zz_32_t ;
reg	RG_zz_32_t_c1 ;
reg	RG_zz_32_t_c2 ;
reg	[8:0]	RG_zz_33_t ;
reg	RG_zz_33_t_c1 ;
reg	RG_zz_33_t_c2 ;
reg	[8:0]	RG_zz_34_t ;
reg	RG_zz_34_t_c1 ;
reg	RG_zz_34_t_c2 ;
reg	[8:0]	RG_zz_35_t ;
reg	RG_zz_35_t_c1 ;
reg	RG_zz_35_t_c2 ;
reg	[8:0]	RG_zz_36_t ;
reg	RG_zz_36_t_c1 ;
reg	RG_zz_36_t_c2 ;
reg	[8:0]	RG_zz_37_t ;
reg	RG_zz_37_t_c1 ;
reg	RG_zz_37_t_c2 ;
reg	[8:0]	RG_zz_38_t ;
reg	RG_zz_38_t_c1 ;
reg	RG_zz_38_t_c2 ;
reg	[8:0]	RG_zz_39_t ;
reg	RG_zz_39_t_c1 ;
reg	RG_zz_39_t_c2 ;
reg	[8:0]	RG_zz_40_t ;
reg	RG_zz_40_t_c1 ;
reg	RG_zz_40_t_c2 ;
reg	[8:0]	RG_zz_41_t ;
reg	RG_zz_41_t_c1 ;
reg	RG_zz_41_t_c2 ;
reg	[8:0]	RG_zz_42_t ;
reg	RG_zz_42_t_c1 ;
reg	RG_zz_42_t_c2 ;
reg	[8:0]	RG_zz_43_t ;
reg	RG_zz_43_t_c1 ;
reg	RG_zz_43_t_c2 ;
reg	[8:0]	RG_zz_44_t ;
reg	RG_zz_44_t_c1 ;
reg	RG_zz_44_t_c2 ;
reg	[8:0]	RG_zz_45_t ;
reg	RG_zz_45_t_c1 ;
reg	RG_zz_45_t_c2 ;
reg	[8:0]	RG_zz_46_t ;
reg	RG_zz_46_t_c1 ;
reg	RG_zz_46_t_c2 ;
reg	[8:0]	RG_zz_47_t ;
reg	RG_zz_47_t_c1 ;
reg	RG_zz_47_t_c2 ;
reg	[8:0]	RG_zz_48_t ;
reg	RG_zz_48_t_c1 ;
reg	RG_zz_48_t_c2 ;
reg	[8:0]	RG_zz_49_t ;
reg	RG_zz_49_t_c1 ;
reg	RG_zz_49_t_c2 ;
reg	[8:0]	RG_zz_50_t ;
reg	RG_zz_50_t_c1 ;
reg	RG_zz_50_t_c2 ;
reg	[8:0]	RG_zz_51_t ;
reg	RG_zz_51_t_c1 ;
reg	RG_zz_51_t_c2 ;
reg	[8:0]	RG_zz_52_t ;
reg	RG_zz_52_t_c1 ;
reg	RG_zz_52_t_c2 ;
reg	[8:0]	RG_zz_53_t ;
reg	RG_zz_53_t_c1 ;
reg	RG_zz_53_t_c2 ;
reg	[8:0]	RG_zz_54_t ;
reg	RG_zz_54_t_c1 ;
reg	RG_zz_54_t_c2 ;
reg	[8:0]	RG_zz_55_t ;
reg	RG_zz_55_t_c1 ;
reg	RG_zz_55_t_c2 ;
reg	[8:0]	RG_zz_56_t ;
reg	RG_zz_56_t_c1 ;
reg	RG_zz_56_t_c2 ;
reg	[8:0]	RG_zz_57_t ;
reg	RG_zz_57_t_c1 ;
reg	RG_zz_57_t_c2 ;
reg	[8:0]	RG_zz_58_t ;
reg	RG_zz_58_t_c1 ;
reg	RG_zz_58_t_c2 ;
reg	[8:0]	RG_zz_59_t ;
reg	RG_zz_59_t_c1 ;
reg	RG_zz_59_t_c2 ;
reg	[8:0]	RG_zz_60_t ;
reg	RG_zz_60_t_c1 ;
reg	RG_zz_60_t_c2 ;
reg	[8:0]	RG_zz_61_t ;
reg	RG_zz_61_t_c1 ;
reg	RG_zz_61_t_c2 ;
reg	[8:0]	RG_zz_62_t ;
reg	RG_zz_62_t_c1 ;
reg	RG_zz_62_t_c2 ;
reg	[3:0]	RG_j_t ;
reg	[2:0]	TR_01 ;
reg	[31:0]	RG_i_k_01_t ;
reg	RG_i_k_01_t_c1 ;
reg	RG_i_k_01_t_c2 ;
reg	RG_i_k_01_t_c3 ;
reg	TR_02 ;
reg	[31:0]	RG_i_j_01_t ;
reg	RG_i_j_01_t_c1 ;
reg	RG_i_j_01_t_c2 ;
reg	RG_i_j_01_t_c3 ;
reg	[8:0]	RG_quantized_block_rl_t ;
reg	[8:0]	RG_quantized_block_rl_t1 ;
reg	[8:0]	RG_quantized_block_rl_1_t ;
reg	[8:0]	RG_quantized_block_rl_1_t1 ;
reg	[8:0]	RG_quantized_block_rl_2_t ;
reg	[8:0]	RG_quantized_block_rl_2_t1 ;
reg	[8:0]	RG_quantized_block_rl_3_t ;
reg	[8:0]	RG_quantized_block_rl_3_t1 ;
reg	[8:0]	RG_quantized_block_rl_4_t ;
reg	[8:0]	RG_quantized_block_rl_4_t1 ;
reg	[8:0]	RG_quantized_block_rl_5_t ;
reg	[8:0]	RG_quantized_block_rl_5_t1 ;
reg	[8:0]	RG_quantized_block_rl_6_t ;
reg	[8:0]	RG_quantized_block_rl_6_t1 ;
reg	[8:0]	RG_quantized_block_rl_7_t ;
reg	[8:0]	RG_quantized_block_rl_7_t1 ;
reg	[8:0]	RG_quantized_block_rl_8_t ;
reg	[8:0]	RG_quantized_block_rl_8_t1 ;
reg	[8:0]	RG_quantized_block_rl_9_t ;
reg	[8:0]	RG_quantized_block_rl_9_t1 ;
reg	[8:0]	RG_quantized_block_rl_10_t ;
reg	[8:0]	RG_quantized_block_rl_10_t1 ;
reg	[8:0]	RG_quantized_block_rl_11_t ;
reg	[8:0]	RG_quantized_block_rl_11_t1 ;
reg	[8:0]	RG_quantized_block_rl_12_t ;
reg	[8:0]	RG_quantized_block_rl_12_t1 ;
reg	[8:0]	RG_quantized_block_rl_13_t ;
reg	[8:0]	RG_quantized_block_rl_13_t1 ;
reg	[8:0]	RG_quantized_block_rl_14_t ;
reg	[8:0]	RG_quantized_block_rl_14_t1 ;
reg	[8:0]	RG_quantized_block_rl_15_t ;
reg	[8:0]	RG_quantized_block_rl_15_t1 ;
reg	[8:0]	RG_quantized_block_rl_16_t ;
reg	[8:0]	RG_quantized_block_rl_16_t1 ;
reg	[8:0]	RG_quantized_block_rl_17_t ;
reg	[8:0]	RG_quantized_block_rl_17_t1 ;
reg	[8:0]	RG_quantized_block_rl_18_t ;
reg	[8:0]	RG_quantized_block_rl_18_t1 ;
reg	[8:0]	RG_quantized_block_rl_19_t ;
reg	[8:0]	RG_quantized_block_rl_19_t1 ;
reg	[8:0]	RG_quantized_block_rl_20_t ;
reg	[8:0]	RG_quantized_block_rl_20_t1 ;
reg	[8:0]	RG_quantized_block_rl_21_t ;
reg	[8:0]	RG_quantized_block_rl_21_t1 ;
reg	[8:0]	RG_quantized_block_rl_22_t ;
reg	[8:0]	RG_quantized_block_rl_22_t1 ;
reg	[8:0]	RG_quantized_block_rl_23_t ;
reg	[8:0]	RG_quantized_block_rl_23_t1 ;
reg	[8:0]	RG_quantized_block_rl_24_t ;
reg	[8:0]	RG_quantized_block_rl_24_t1 ;
reg	[8:0]	RG_quantized_block_rl_25_t ;
reg	[8:0]	RG_quantized_block_rl_25_t1 ;
reg	[8:0]	RG_quantized_block_rl_26_t ;
reg	[8:0]	RG_quantized_block_rl_26_t1 ;
reg	[8:0]	RG_quantized_block_rl_27_t ;
reg	[8:0]	RG_quantized_block_rl_27_t1 ;
reg	[8:0]	RG_quantized_block_rl_28_t ;
reg	[8:0]	RG_quantized_block_rl_28_t1 ;
reg	[8:0]	RG_quantized_block_rl_29_t ;
reg	[8:0]	RG_quantized_block_rl_29_t1 ;
reg	[8:0]	RG_quantized_block_rl_30_t ;
reg	[8:0]	RG_quantized_block_rl_30_t1 ;
reg	[8:0]	RG_quantized_block_rl_31_t ;
reg	[8:0]	RG_quantized_block_rl_31_t1 ;
reg	[8:0]	RG_quantized_block_rl_32_t ;
reg	[8:0]	RG_quantized_block_rl_32_t1 ;
reg	[8:0]	RG_quantized_block_rl_33_t ;
reg	[8:0]	RG_quantized_block_rl_33_t1 ;
reg	[8:0]	RG_quantized_block_rl_34_t ;
reg	[8:0]	RG_quantized_block_rl_34_t1 ;
reg	[8:0]	RG_quantized_block_rl_35_t ;
reg	[8:0]	RG_quantized_block_rl_35_t1 ;
reg	[8:0]	RG_quantized_block_rl_36_t ;
reg	[8:0]	RG_quantized_block_rl_36_t1 ;
reg	[8:0]	RG_quantized_block_rl_37_t ;
reg	[8:0]	RG_quantized_block_rl_37_t1 ;
reg	[8:0]	RG_quantized_block_rl_38_t ;
reg	[8:0]	RG_quantized_block_rl_38_t1 ;
reg	[8:0]	RG_quantized_block_rl_39_t ;
reg	[8:0]	RG_quantized_block_rl_39_t1 ;
reg	[8:0]	RG_quantized_block_rl_40_t ;
reg	[8:0]	RG_quantized_block_rl_40_t1 ;
reg	[8:0]	RG_quantized_block_rl_41_t ;
reg	[8:0]	RG_quantized_block_rl_41_t1 ;
reg	[8:0]	RG_quantized_block_rl_42_t ;
reg	[8:0]	RG_quantized_block_rl_42_t1 ;
reg	[8:0]	RG_quantized_block_rl_43_t ;
reg	[8:0]	RG_quantized_block_rl_43_t1 ;
reg	[8:0]	RG_quantized_block_rl_44_t ;
reg	[8:0]	RG_quantized_block_rl_44_t1 ;
reg	[8:0]	RG_quantized_block_rl_45_t ;
reg	[8:0]	RG_quantized_block_rl_45_t1 ;
reg	[8:0]	RG_quantized_block_rl_46_t ;
reg	[8:0]	RG_quantized_block_rl_46_t1 ;
reg	[8:0]	RG_quantized_block_rl_47_t ;
reg	[8:0]	RG_quantized_block_rl_47_t1 ;
reg	[8:0]	RG_quantized_block_rl_48_t ;
reg	[8:0]	RG_quantized_block_rl_48_t1 ;
reg	[8:0]	RG_quantized_block_rl_49_t ;
reg	[8:0]	RG_quantized_block_rl_49_t1 ;
reg	[8:0]	RG_quantized_block_rl_50_t ;
reg	[8:0]	RG_quantized_block_rl_50_t1 ;
reg	[8:0]	RG_quantized_block_rl_51_t ;
reg	[8:0]	RG_quantized_block_rl_51_t1 ;
reg	[8:0]	RG_quantized_block_rl_52_t ;
reg	[8:0]	RG_quantized_block_rl_52_t1 ;
reg	[8:0]	RG_quantized_block_rl_53_t ;
reg	[8:0]	RG_quantized_block_rl_53_t1 ;
reg	[8:0]	RG_quantized_block_rl_54_t ;
reg	[8:0]	RG_quantized_block_rl_54_t1 ;
reg	[8:0]	RG_quantized_block_rl_55_t ;
reg	[8:0]	RG_quantized_block_rl_55_t1 ;
reg	[8:0]	RG_quantized_block_rl_56_t ;
reg	[8:0]	RG_quantized_block_rl_56_t1 ;
reg	[8:0]	RG_quantized_block_rl_57_t ;
reg	[8:0]	RG_quantized_block_rl_57_t1 ;
reg	[8:0]	RG_quantized_block_rl_58_t ;
reg	[8:0]	RG_quantized_block_rl_58_t1 ;
reg	[8:0]	RG_quantized_block_rl_59_t ;
reg	[8:0]	RG_quantized_block_rl_59_t1 ;
reg	[8:0]	RG_quantized_block_rl_60_t ;
reg	[8:0]	RG_quantized_block_rl_60_t1 ;
reg	[8:0]	RG_quantized_block_rl_61_t ;
reg	[8:0]	RG_quantized_block_rl_61_t1 ;
reg	[8:0]	RG_k_quantized_block_rl_01_t ;
reg	[8:0]	RG_k_quantized_block_rl_01_t1 ;
reg	[8:0]	RG_k_quantized_block_rl_01_t2 ;
reg	[8:0]	RG_quantized_block_rl_zz_t ;
reg	[5:0]	RG_k_t ;
reg	FF_d_t ;
reg	FF_d_t_c1 ;
reg	FF_d_t_c2 ;
reg	[8:0]	RG_previous_dc_rl_t ;
reg	[8:0]	RG_previous_dc_rl_t1 ;
reg	[8:0]	RG_rl_128_t ;
reg	[8:0]	RG_rl_128_t1 ;
reg	[8:0]	RG_rl_129_t ;
reg	[8:0]	RG_rl_129_t1 ;
reg	[8:0]	RG_rl_130_t ;
reg	[8:0]	RG_rl_130_t1 ;
reg	[8:0]	RG_rl_131_t ;
reg	[8:0]	RG_rl_131_t1 ;
reg	[8:0]	RG_rl_132_t ;
reg	[8:0]	RG_rl_132_t1 ;
reg	[8:0]	RG_rl_133_t ;
reg	[8:0]	RG_rl_133_t1 ;
reg	[8:0]	RG_rl_134_t ;
reg	[8:0]	RG_rl_134_t1 ;
reg	[8:0]	RG_rl_135_t ;
reg	[8:0]	RG_rl_135_t1 ;
reg	[8:0]	RG_rl_136_t ;
reg	[8:0]	RG_rl_136_t1 ;
reg	[8:0]	RG_rl_137_t ;
reg	[8:0]	RG_rl_137_t1 ;
reg	[8:0]	RG_rl_138_t ;
reg	[8:0]	RG_rl_138_t1 ;
reg	[8:0]	RG_rl_139_t ;
reg	[8:0]	RG_rl_139_t1 ;
reg	[8:0]	RG_rl_140_t ;
reg	[8:0]	RG_rl_140_t1 ;
reg	[8:0]	RG_rl_141_t ;
reg	[8:0]	RG_rl_141_t1 ;
reg	[8:0]	RG_rl_142_t ;
reg	[8:0]	RG_rl_142_t1 ;
reg	[8:0]	RG_rl_143_t ;
reg	[8:0]	RG_rl_143_t1 ;
reg	[8:0]	RG_rl_144_t ;
reg	[8:0]	RG_rl_144_t1 ;
reg	[8:0]	RG_rl_145_t ;
reg	[8:0]	RG_rl_145_t1 ;
reg	[8:0]	RG_rl_146_t ;
reg	[8:0]	RG_rl_146_t1 ;
reg	[8:0]	RG_rl_147_t ;
reg	[8:0]	RG_rl_147_t1 ;
reg	[8:0]	RG_rl_148_t ;
reg	[8:0]	RG_rl_148_t1 ;
reg	[8:0]	RG_rl_149_t ;
reg	[8:0]	RG_rl_149_t1 ;
reg	[8:0]	RG_rl_150_t ;
reg	[8:0]	RG_rl_150_t1 ;
reg	[8:0]	RG_rl_151_t ;
reg	[8:0]	RG_rl_151_t1 ;
reg	[8:0]	RG_rl_152_t ;
reg	[8:0]	RG_rl_152_t1 ;
reg	[8:0]	RG_rl_153_t ;
reg	[8:0]	RG_rl_153_t1 ;
reg	[8:0]	RG_rl_154_t ;
reg	[8:0]	RG_rl_154_t1 ;
reg	[8:0]	RG_rl_155_t ;
reg	[8:0]	RG_rl_155_t1 ;
reg	[8:0]	RG_rl_156_t ;
reg	[8:0]	RG_rl_156_t1 ;
reg	[8:0]	RG_rl_157_t ;
reg	[8:0]	RG_rl_157_t1 ;
reg	[8:0]	RG_rl_158_t ;
reg	[8:0]	RG_rl_158_t1 ;
reg	[8:0]	RG_rl_159_t ;
reg	[8:0]	RG_rl_159_t1 ;
reg	[8:0]	RG_rl_160_t ;
reg	[8:0]	RG_rl_160_t1 ;
reg	[8:0]	RG_rl_161_t ;
reg	[8:0]	RG_rl_161_t1 ;
reg	[8:0]	RG_rl_162_t ;
reg	[8:0]	RG_rl_162_t1 ;
reg	[8:0]	RG_rl_163_t ;
reg	[8:0]	RG_rl_163_t1 ;
reg	[8:0]	RG_rl_164_t ;
reg	[8:0]	RG_rl_164_t1 ;
reg	[8:0]	RG_rl_165_t ;
reg	[8:0]	RG_rl_165_t1 ;
reg	[8:0]	RG_rl_166_t ;
reg	[8:0]	RG_rl_166_t1 ;
reg	[8:0]	RG_rl_167_t ;
reg	[8:0]	RG_rl_167_t1 ;
reg	[8:0]	RG_rl_168_t ;
reg	[8:0]	RG_rl_168_t1 ;
reg	[8:0]	RG_rl_169_t ;
reg	[8:0]	RG_rl_169_t1 ;
reg	[8:0]	RG_rl_170_t ;
reg	[8:0]	RG_rl_170_t1 ;
reg	[8:0]	RG_rl_171_t ;
reg	[8:0]	RG_rl_171_t1 ;
reg	[8:0]	RG_rl_172_t ;
reg	[8:0]	RG_rl_172_t1 ;
reg	[8:0]	RG_rl_173_t ;
reg	[8:0]	RG_rl_173_t1 ;
reg	[8:0]	RG_rl_174_t ;
reg	[8:0]	RG_rl_174_t1 ;
reg	[8:0]	RG_rl_175_t ;
reg	[8:0]	RG_rl_175_t1 ;
reg	[8:0]	RG_rl_176_t ;
reg	[8:0]	RG_rl_176_t1 ;
reg	[8:0]	RG_rl_177_t ;
reg	[8:0]	RG_rl_177_t1 ;
reg	[8:0]	RG_rl_178_t ;
reg	[8:0]	RG_rl_178_t1 ;
reg	[8:0]	RG_rl_179_t ;
reg	[8:0]	RG_rl_179_t1 ;
reg	[8:0]	RG_rl_180_t ;
reg	[8:0]	RG_rl_180_t1 ;
reg	[8:0]	RG_rl_181_t ;
reg	[8:0]	RG_rl_181_t1 ;
reg	[8:0]	RG_rl_182_t ;
reg	[8:0]	RG_rl_182_t1 ;
reg	[8:0]	RG_rl_183_t ;
reg	[8:0]	RG_rl_183_t1 ;
reg	[8:0]	RG_rl_184_t ;
reg	[8:0]	RG_rl_184_t1 ;
reg	[8:0]	RG_rl_185_t ;
reg	[8:0]	RG_rl_185_t1 ;
reg	[8:0]	RG_rl_186_t ;
reg	[8:0]	RG_rl_186_t1 ;
reg	[8:0]	RG_rl_187_t ;
reg	[8:0]	RG_rl_187_t1 ;
reg	[8:0]	RG_rl_188_t ;
reg	[8:0]	RG_rl_188_t1 ;
reg	[8:0]	RG_rl_189_t ;
reg	[8:0]	RG_rl_189_t1 ;
reg	[8:0]	RG_rl_190_t ;
reg	[8:0]	RG_rl_190_t1 ;
reg	[8:0]	RG_rl_191_t ;
reg	[8:0]	RG_rl_191_t1 ;
reg	[7:0]	RG_len_t ;
reg	[7:0]	RG_len_1_t ;
reg	[6:0]	RG_k_1_t ;
reg	[8:0]	TR_04 ;
reg	[8:0]	TR_05 ;
reg	[8:0]	TR_06 ;
reg	[8:0]	TR_07 ;
reg	[8:0]	TR_08 ;
reg	[8:0]	TR_09 ;
reg	[8:0]	TR_10 ;
reg	[8:0]	TR_11 ;
reg	[8:0]	M_184 ;
reg	M_184_c1 ;
reg	M_184_c2 ;
reg	M_184_c3 ;
reg	M_184_c4 ;
reg	M_184_c5 ;
reg	M_184_c6 ;
reg	M_184_c7 ;
reg	M_184_c8 ;
reg	M_02_t128 ;
reg	M_02_t128_t1 ;
reg	M_01_t64 ;
reg	M_01_t64_t1 ;
reg	M_03_t128 ;
reg	M_03_t128_t1 ;
reg	valid_r_t ;
reg	[5:0]	TR_03 ;
reg	[7:0]	incr8u3i1 ;
reg	incr8u3i1_c1 ;
reg	[6:0]	sub8u_7_11i1 ;

jpeg_sub8u_7_1 INST_sub8u_7_1_1 ( .i1(sub8u_7_11i1) ,.i2(sub8u_7_11i2) ,.o1(sub8u_7_11ot) );	// line#=../rle.cpp:77,78,83,84
jpeg_sub8u_7 INST_sub8u_7_1 ( .i1(sub8u_71i1) ,.i2(sub8u_71i2) ,.o1(sub8u_71ot) );	// line#=../rle.cpp:83,84
jpeg_decr32s INST_decr32s_1 ( .i1(decr32s1i1) ,.o1(decr32s1ot) );	// line#=../rle.cpp:124,155
jpeg_decr32s INST_decr32s_2 ( .i1(decr32s2i1) ,.o1(decr32s2ot) );	// line#=../rle.cpp:130,161
jpeg_decr8u_7 INST_decr8u_7_1 ( .i1(decr8u_71i1) ,.o1(decr8u_71ot) );	// line#=../rle.cpp:77,78
jpeg_incr32s INST_incr32s_1 ( .i1(incr32s1i1) ,.o1(incr32s1ot) );	// line#=../rle.cpp:61,62,63,74,114,125
									// ,145,156
jpeg_incr32s INST_incr32s_2 ( .i1(incr32s2i1) ,.o1(incr32s2ot) );	// line#=../rle.cpp:64,119,129,150,160
jpeg_incr8u INST_incr8u_1 ( .i1(incr8u1i1) ,.o1(incr8u1ot) );	// line#=../rle.cpp:68,79
jpeg_incr8u INST_incr8u_2 ( .i1(incr8u2i1) ,.o1(incr8u2ot) );	// line#=../rle.cpp:73
jpeg_incr8u INST_incr8u_3 ( .i1(incr8u3i1) ,.o1(incr8u3ot) );	// line#=../rle.cpp:74,111,142
jpeg_incr8u INST_incr8u_4 ( .i1(incr8u4i1) ,.o1(incr8u4ot) );	// line#=../rle.cpp:69,80
jpeg_incr4s INST_incr4s_1 ( .i1(incr4s1i1) ,.o1(incr4s1ot) );	// line#=../rle.cpp:34
jpeg_lop8u_1 INST_lop8u_1_1 ( .i1(lop8u_11i1) ,.i2(lop8u_11i2) ,.o1(lop8u_11ot) );	// line#=../rle.cpp:109,110
assign	lop8u_11ot_port = lop8u_11ot ;
jpeg_sub12s_9 INST_sub12s_9_1 ( .i1(sub12s_91i1) ,.i2(sub12s_91i2) ,.o1(sub12s_91ot) );	// line#=../rle.cpp:52
jpeg_sub8u INST_sub8u_1 ( .i1(sub8u1i1) ,.i2(sub8u1i2) ,.o1(sub8u1ot) );	// line#=../rle.cpp:86
assign	jpeg_out_a00 = jpeg_out_a00_r ;	// line#=../rle.h:60
assign	jpeg_out_a01 = jpeg_out_a01_r ;	// line#=../rle.h:60
assign	jpeg_out_a02 = jpeg_out_a02_r ;	// line#=../rle.h:60
assign	jpeg_out_a03 = jpeg_out_a03_r ;	// line#=../rle.h:60
assign	jpeg_out_a04 = jpeg_out_a04_r ;	// line#=../rle.h:60
assign	jpeg_out_a05 = jpeg_out_a05_r ;	// line#=../rle.h:60
assign	jpeg_out_a06 = jpeg_out_a06_r ;	// line#=../rle.h:60
assign	jpeg_out_a07 = jpeg_out_a07_r ;	// line#=../rle.h:60
assign	jpeg_out_a08 = jpeg_out_a08_r ;	// line#=../rle.h:60
assign	jpeg_out_a09 = jpeg_out_a09_r ;	// line#=../rle.h:60
assign	jpeg_out_a10 = jpeg_out_a10_r ;	// line#=../rle.h:60
assign	jpeg_out_a11 = jpeg_out_a11_r ;	// line#=../rle.h:60
assign	jpeg_out_a12 = jpeg_out_a12_r ;	// line#=../rle.h:60
assign	jpeg_out_a13 = jpeg_out_a13_r ;	// line#=../rle.h:60
assign	jpeg_out_a14 = jpeg_out_a14_r ;	// line#=../rle.h:60
assign	jpeg_out_a15 = jpeg_out_a15_r ;	// line#=../rle.h:60
assign	jpeg_out_a16 = jpeg_out_a16_r ;	// line#=../rle.h:60
assign	jpeg_out_a17 = jpeg_out_a17_r ;	// line#=../rle.h:60
assign	jpeg_out_a18 = jpeg_out_a18_r ;	// line#=../rle.h:60
assign	jpeg_out_a19 = jpeg_out_a19_r ;	// line#=../rle.h:60
assign	jpeg_out_a20 = jpeg_out_a20_r ;	// line#=../rle.h:60
assign	jpeg_out_a21 = jpeg_out_a21_r ;	// line#=../rle.h:60
assign	jpeg_out_a22 = jpeg_out_a22_r ;	// line#=../rle.h:60
assign	jpeg_out_a23 = jpeg_out_a23_r ;	// line#=../rle.h:60
assign	jpeg_out_a24 = jpeg_out_a24_r ;	// line#=../rle.h:60
assign	jpeg_out_a25 = jpeg_out_a25_r ;	// line#=../rle.h:60
assign	jpeg_out_a26 = jpeg_out_a26_r ;	// line#=../rle.h:60
assign	jpeg_out_a27 = jpeg_out_a27_r ;	// line#=../rle.h:60
assign	jpeg_out_a28 = jpeg_out_a28_r ;	// line#=../rle.h:60
assign	jpeg_out_a29 = jpeg_out_a29_r ;	// line#=../rle.h:60
assign	jpeg_out_a30 = jpeg_out_a30_r ;	// line#=../rle.h:60
assign	jpeg_out_a31 = jpeg_out_a31_r ;	// line#=../rle.h:60
assign	jpeg_out_a32 = jpeg_out_a32_r ;	// line#=../rle.h:60
assign	jpeg_out_a33 = jpeg_out_a33_r ;	// line#=../rle.h:60
assign	jpeg_out_a34 = jpeg_out_a34_r ;	// line#=../rle.h:60
assign	jpeg_out_a35 = jpeg_out_a35_r ;	// line#=../rle.h:60
assign	jpeg_out_a36 = jpeg_out_a36_r ;	// line#=../rle.h:60
assign	jpeg_out_a37 = jpeg_out_a37_r ;	// line#=../rle.h:60
assign	jpeg_out_a38 = jpeg_out_a38_r ;	// line#=../rle.h:60
assign	jpeg_out_a39 = jpeg_out_a39_r ;	// line#=../rle.h:60
assign	jpeg_out_a40 = jpeg_out_a40_r ;	// line#=../rle.h:60
assign	jpeg_out_a41 = jpeg_out_a41_r ;	// line#=../rle.h:60
assign	jpeg_out_a42 = jpeg_out_a42_r ;	// line#=../rle.h:60
assign	jpeg_out_a43 = jpeg_out_a43_r ;	// line#=../rle.h:60
assign	jpeg_out_a44 = jpeg_out_a44_r ;	// line#=../rle.h:60
assign	jpeg_out_a45 = jpeg_out_a45_r ;	// line#=../rle.h:60
assign	jpeg_out_a46 = jpeg_out_a46_r ;	// line#=../rle.h:60
assign	jpeg_out_a47 = jpeg_out_a47_r ;	// line#=../rle.h:60
assign	jpeg_out_a48 = jpeg_out_a48_r ;	// line#=../rle.h:60
assign	jpeg_out_a49 = jpeg_out_a49_r ;	// line#=../rle.h:60
assign	jpeg_out_a50 = jpeg_out_a50_r ;	// line#=../rle.h:60
assign	jpeg_out_a51 = jpeg_out_a51_r ;	// line#=../rle.h:60
assign	jpeg_out_a52 = jpeg_out_a52_r ;	// line#=../rle.h:60
assign	jpeg_out_a53 = jpeg_out_a53_r ;	// line#=../rle.h:60
assign	jpeg_out_a54 = jpeg_out_a54_r ;	// line#=../rle.h:60
assign	jpeg_out_a55 = jpeg_out_a55_r ;	// line#=../rle.h:60
assign	jpeg_out_a56 = jpeg_out_a56_r ;	// line#=../rle.h:60
assign	jpeg_out_a57 = jpeg_out_a57_r ;	// line#=../rle.h:60
assign	jpeg_out_a58 = jpeg_out_a58_r ;	// line#=../rle.h:60
assign	jpeg_out_a59 = jpeg_out_a59_r ;	// line#=../rle.h:60
assign	jpeg_out_a60 = jpeg_out_a60_r ;	// line#=../rle.h:60
assign	jpeg_out_a61 = jpeg_out_a61_r ;	// line#=../rle.h:60
assign	jpeg_out_a62 = jpeg_out_a62_r ;	// line#=../rle.h:60
assign	jpeg_out_a63 = jpeg_out_a63_r ;	// line#=../rle.h:60
assign	jpeg_out_a64 = jpeg_out_a64_r ;	// line#=../rle.h:60
assign	jpeg_out_a65 = jpeg_out_a65_r ;	// line#=../rle.h:60
assign	jpeg_out_a66 = jpeg_out_a66_r ;	// line#=../rle.h:60
assign	jpeg_out_a67 = jpeg_out_a67_r ;	// line#=../rle.h:60
assign	jpeg_out_a68 = jpeg_out_a68_r ;	// line#=../rle.h:60
assign	jpeg_out_a69 = jpeg_out_a69_r ;	// line#=../rle.h:60
assign	jpeg_out_a70 = jpeg_out_a70_r ;	// line#=../rle.h:60
assign	jpeg_out_a71 = jpeg_out_a71_r ;	// line#=../rle.h:60
assign	jpeg_out_a72 = jpeg_out_a72_r ;	// line#=../rle.h:60
assign	jpeg_out_a73 = jpeg_out_a73_r ;	// line#=../rle.h:60
assign	jpeg_out_a74 = jpeg_out_a74_r ;	// line#=../rle.h:60
assign	jpeg_out_a75 = jpeg_out_a75_r ;	// line#=../rle.h:60
assign	jpeg_out_a76 = jpeg_out_a76_r ;	// line#=../rle.h:60
assign	jpeg_out_a77 = jpeg_out_a77_r ;	// line#=../rle.h:60
assign	jpeg_out_a78 = jpeg_out_a78_r ;	// line#=../rle.h:60
assign	jpeg_out_a79 = jpeg_out_a79_r ;	// line#=../rle.h:60
assign	jpeg_out_a80 = jpeg_out_a80_r ;	// line#=../rle.h:60
assign	jpeg_out_a81 = jpeg_out_a81_r ;	// line#=../rle.h:60
assign	jpeg_out_a82 = jpeg_out_a82_r ;	// line#=../rle.h:60
assign	jpeg_out_a83 = jpeg_out_a83_r ;	// line#=../rle.h:60
assign	jpeg_out_a84 = jpeg_out_a84_r ;	// line#=../rle.h:60
assign	jpeg_out_a85 = jpeg_out_a85_r ;	// line#=../rle.h:60
assign	jpeg_out_a86 = jpeg_out_a86_r ;	// line#=../rle.h:60
assign	jpeg_out_a87 = jpeg_out_a87_r ;	// line#=../rle.h:60
assign	jpeg_out_a88 = jpeg_out_a88_r ;	// line#=../rle.h:60
assign	jpeg_out_a89 = jpeg_out_a89_r ;	// line#=../rle.h:60
assign	jpeg_out_a90 = jpeg_out_a90_r ;	// line#=../rle.h:60
assign	jpeg_out_a91 = jpeg_out_a91_r ;	// line#=../rle.h:60
assign	jpeg_out_a92 = jpeg_out_a92_r ;	// line#=../rle.h:60
assign	jpeg_out_a93 = jpeg_out_a93_r ;	// line#=../rle.h:60
assign	jpeg_out_a94 = jpeg_out_a94_r ;	// line#=../rle.h:60
assign	jpeg_out_a95 = jpeg_out_a95_r ;	// line#=../rle.h:60
assign	jpeg_out_a96 = jpeg_out_a96_r ;	// line#=../rle.h:60
assign	jpeg_out_a97 = jpeg_out_a97_r ;	// line#=../rle.h:60
assign	jpeg_out_a98 = jpeg_out_a98_r ;	// line#=../rle.h:60
assign	jpeg_out_a99 = jpeg_out_a99_r ;	// line#=../rle.h:60
assign	jpeg_out_a100 = jpeg_out_a100_r ;	// line#=../rle.h:60
assign	jpeg_out_a101 = jpeg_out_a101_r ;	// line#=../rle.h:60
assign	jpeg_out_a102 = jpeg_out_a102_r ;	// line#=../rle.h:60
assign	jpeg_out_a103 = jpeg_out_a103_r ;	// line#=../rle.h:60
assign	jpeg_out_a104 = jpeg_out_a104_r ;	// line#=../rle.h:60
assign	jpeg_out_a105 = jpeg_out_a105_r ;	// line#=../rle.h:60
assign	jpeg_out_a106 = jpeg_out_a106_r ;	// line#=../rle.h:60
assign	jpeg_out_a107 = jpeg_out_a107_r ;	// line#=../rle.h:60
assign	jpeg_out_a108 = jpeg_out_a108_r ;	// line#=../rle.h:60
assign	jpeg_out_a109 = jpeg_out_a109_r ;	// line#=../rle.h:60
assign	jpeg_out_a110 = jpeg_out_a110_r ;	// line#=../rle.h:60
assign	jpeg_out_a111 = jpeg_out_a111_r ;	// line#=../rle.h:60
assign	jpeg_out_a112 = jpeg_out_a112_r ;	// line#=../rle.h:60
assign	jpeg_out_a113 = jpeg_out_a113_r ;	// line#=../rle.h:60
assign	jpeg_out_a114 = jpeg_out_a114_r ;	// line#=../rle.h:60
assign	jpeg_out_a115 = jpeg_out_a115_r ;	// line#=../rle.h:60
assign	jpeg_out_a116 = jpeg_out_a116_r ;	// line#=../rle.h:60
assign	jpeg_out_a117 = jpeg_out_a117_r ;	// line#=../rle.h:60
assign	jpeg_out_a118 = jpeg_out_a118_r ;	// line#=../rle.h:60
assign	jpeg_out_a119 = jpeg_out_a119_r ;	// line#=../rle.h:60
assign	jpeg_out_a120 = jpeg_out_a120_r ;	// line#=../rle.h:60
assign	jpeg_out_a121 = jpeg_out_a121_r ;	// line#=../rle.h:60
assign	jpeg_out_a122 = jpeg_out_a122_r ;	// line#=../rle.h:60
assign	jpeg_out_a123 = jpeg_out_a123_r ;	// line#=../rle.h:60
assign	jpeg_out_a124 = jpeg_out_a124_r ;	// line#=../rle.h:60
assign	jpeg_out_a125 = jpeg_out_a125_r ;	// line#=../rle.h:60
assign	jpeg_out_a126 = jpeg_out_a126_r ;	// line#=../rle.h:60
assign	jpeg_out_a127 = jpeg_out_a127_r ;	// line#=../rle.h:60
assign	jpeg_len_out = jpeg_len_out_r ;	// line#=../rle.h:61
assign	valid = valid_r ;	// line#=../rle.h:62
assign	CT_03 = ( ( ~|RG_i_j_01 ) & M_39 ) ;	// line#=../rle.cpp:117,118
assign	M_39 = ~|{ ( RG_i_k_01 [31] & RG_i_k_01 [0] ) , ~RG_i_k_01 [0] } ;	// line#=../rle.cpp:117,118,148,149
assign	CT_18 = ( ( ~|{ RG_i_j_01 [31:3] , ~RG_i_j_01 [2:0] } ) & M_39 ) ;	// line#=../rle.cpp:148,149
assign	M_49 = ~|RG_quantized_block_rl ;	// line#=../rle.cpp:77,78
assign	M_50 = ~|RG_quantized_block_rl_1 ;	// line#=../rle.cpp:77,78
assign	M_51 = ~|RG_quantized_block_rl_2 ;	// line#=../rle.cpp:77,78
assign	M_52 = ~|RG_quantized_block_rl_3 ;	// line#=../rle.cpp:77,78
assign	M_53 = ~|RG_quantized_block_rl_4 ;	// line#=../rle.cpp:77,78
assign	M_54 = ~|RG_quantized_block_rl_5 ;	// line#=../rle.cpp:77,78
assign	M_55 = ~|RG_quantized_block_rl_6 ;	// line#=../rle.cpp:77,78
assign	M_56 = ~|RG_quantized_block_rl_7 ;	// line#=../rle.cpp:77,78
assign	M_57 = ~|RG_quantized_block_rl_8 ;	// line#=../rle.cpp:77,78
assign	M_58 = ~|RG_quantized_block_rl_9 ;	// line#=../rle.cpp:77,78
assign	M_59 = ~|RG_quantized_block_rl_10 ;	// line#=../rle.cpp:77,78
assign	M_60 = ~|RG_quantized_block_rl_11 ;	// line#=../rle.cpp:77,78
assign	M_61 = ~|RG_quantized_block_rl_12 ;	// line#=../rle.cpp:77,78
assign	M_62 = ~|RG_quantized_block_rl_13 ;	// line#=../rle.cpp:77,78
assign	M_63 = ~|RG_quantized_block_rl_14 ;	// line#=../rle.cpp:77,78
assign	M_64 = ~|RG_quantized_block_rl_15 ;	// line#=../rle.cpp:77,78
assign	M_65 = ~|RG_quantized_block_rl_16 ;	// line#=../rle.cpp:77,78
assign	M_66 = ~|RG_quantized_block_rl_17 ;	// line#=../rle.cpp:77,78
assign	M_67 = ~|RG_quantized_block_rl_18 ;	// line#=../rle.cpp:77,78
assign	M_68 = ~|RG_quantized_block_rl_19 ;	// line#=../rle.cpp:77,78
assign	M_69 = ~|RG_quantized_block_rl_20 ;	// line#=../rle.cpp:77,78
assign	M_70 = ~|RG_quantized_block_rl_21 ;	// line#=../rle.cpp:77,78
assign	M_71 = ~|RG_quantized_block_rl_22 ;	// line#=../rle.cpp:77,78
assign	M_72 = ~|RG_quantized_block_rl_23 ;	// line#=../rle.cpp:77,78
assign	M_73 = ~|RG_quantized_block_rl_24 ;	// line#=../rle.cpp:77,78
assign	M_74 = ~|RG_quantized_block_rl_25 ;	// line#=../rle.cpp:77,78
assign	M_75 = ~|RG_quantized_block_rl_26 ;	// line#=../rle.cpp:77,78
assign	M_76 = ~|RG_quantized_block_rl_27 ;	// line#=../rle.cpp:77,78
assign	M_77 = ~|RG_quantized_block_rl_28 ;	// line#=../rle.cpp:77,78
assign	M_78 = ~|RG_quantized_block_rl_29 ;	// line#=../rle.cpp:77,78
assign	M_79 = ~|RG_quantized_block_rl_30 ;	// line#=../rle.cpp:77,78
assign	M_80 = ~|RG_quantized_block_rl_31 ;	// line#=../rle.cpp:77,78
assign	M_81 = ~|RG_quantized_block_rl_32 ;	// line#=../rle.cpp:77,78
assign	M_82 = ~|RG_quantized_block_rl_33 ;	// line#=../rle.cpp:77,78
assign	M_83 = ~|RG_quantized_block_rl_34 ;	// line#=../rle.cpp:77,78
assign	M_84 = ~|RG_quantized_block_rl_35 ;	// line#=../rle.cpp:77,78
assign	M_85 = ~|RG_quantized_block_rl_36 ;	// line#=../rle.cpp:77,78
assign	M_86 = ~|RG_quantized_block_rl_37 ;	// line#=../rle.cpp:77,78
assign	M_87 = ~|RG_quantized_block_rl_38 ;	// line#=../rle.cpp:77,78
assign	M_88 = ~|RG_quantized_block_rl_39 ;	// line#=../rle.cpp:77,78
assign	M_89 = ~|RG_quantized_block_rl_40 ;	// line#=../rle.cpp:77,78
assign	M_90 = ~|RG_quantized_block_rl_41 ;	// line#=../rle.cpp:77,78
assign	M_91 = ~|RG_quantized_block_rl_42 ;	// line#=../rle.cpp:77,78
assign	M_92 = ~|RG_quantized_block_rl_43 ;	// line#=../rle.cpp:77,78
assign	M_93 = ~|RG_quantized_block_rl_44 ;	// line#=../rle.cpp:77,78
assign	M_94 = ~|RG_quantized_block_rl_45 ;	// line#=../rle.cpp:77,78
assign	M_95 = ~|RG_quantized_block_rl_46 ;	// line#=../rle.cpp:77,78
assign	M_96 = ~|RG_quantized_block_rl_47 ;	// line#=../rle.cpp:77,78
assign	M_97 = ~|RG_quantized_block_rl_48 ;	// line#=../rle.cpp:77,78
assign	M_98 = ~|RG_quantized_block_rl_49 ;	// line#=../rle.cpp:77,78
assign	M_99 = ~|RG_quantized_block_rl_50 ;	// line#=../rle.cpp:77,78
assign	M_100 = ~|RG_quantized_block_rl_51 ;	// line#=../rle.cpp:77,78
assign	M_102 = ~|RG_quantized_block_rl_52 ;	// line#=../rle.cpp:77,78
assign	M_103 = ~|RG_quantized_block_rl_53 ;	// line#=../rle.cpp:77,78
assign	M_104 = ~|RG_quantized_block_rl_54 ;	// line#=../rle.cpp:77,78
assign	M_105 = ~|RG_quantized_block_rl_55 ;	// line#=../rle.cpp:77,78
assign	M_106 = ~|RG_quantized_block_rl_56 ;	// line#=../rle.cpp:77,78
assign	M_107 = ~|RG_quantized_block_rl_57 ;	// line#=../rle.cpp:77,78
assign	M_108 = ~|RG_quantized_block_rl_58 ;	// line#=../rle.cpp:77,78
assign	M_109 = ~|RG_quantized_block_rl_59 ;	// line#=../rle.cpp:77,78
assign	M_110 = ~|RG_quantized_block_rl_60 ;	// line#=../rle.cpp:77,78
assign	M_112 = ~|RG_quantized_block_rl_61 ;	// line#=../rle.cpp:77,78
assign	M_113 = ~|RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:77,78
assign	M_114 = ~|RG_previous_dc_rl ;	// line#=../rle.cpp:77,78
assign	M_115 = ~|RG_rl_128 ;	// line#=../rle.cpp:77,78
assign	M_116 = ~|RG_rl_129 ;	// line#=../rle.cpp:77,78
assign	M_117 = ~|RG_rl_130 ;	// line#=../rle.cpp:77,78
assign	M_118 = ~|RG_rl_131 ;	// line#=../rle.cpp:77,78
assign	M_119 = ~|RG_rl_132 ;	// line#=../rle.cpp:77,78
assign	M_120 = ~|RG_rl_133 ;	// line#=../rle.cpp:77,78
assign	M_122 = ~|RG_rl_134 ;	// line#=../rle.cpp:77,78
assign	M_123 = ~|RG_rl_135 ;	// line#=../rle.cpp:77,78
assign	M_124 = ~|RG_rl_136 ;	// line#=../rle.cpp:77,78
assign	M_125 = ~|RG_rl_137 ;	// line#=../rle.cpp:77,78
assign	M_126 = ~|RG_rl_138 ;	// line#=../rle.cpp:77,78
assign	M_127 = ~|RG_rl_139 ;	// line#=../rle.cpp:77,78
assign	M_128 = ~|RG_rl_140 ;	// line#=../rle.cpp:77,78
assign	M_129 = ~|RG_rl_141 ;	// line#=../rle.cpp:77,78
assign	M_130 = ~|RG_rl_142 ;	// line#=../rle.cpp:77,78
assign	M_131 = ~|RG_rl_143 ;	// line#=../rle.cpp:77,78
assign	M_132 = ~|RG_rl_144 ;	// line#=../rle.cpp:77,78
assign	M_133 = ~|RG_rl_145 ;	// line#=../rle.cpp:77,78
assign	M_134 = ~|RG_rl_146 ;	// line#=../rle.cpp:77,78
assign	M_135 = ~|RG_rl_147 ;	// line#=../rle.cpp:77,78
assign	M_136 = ~|RG_rl_148 ;	// line#=../rle.cpp:77,78
assign	M_137 = ~|RG_rl_149 ;	// line#=../rle.cpp:77,78
assign	M_138 = ~|RG_rl_150 ;	// line#=../rle.cpp:77,78
assign	M_139 = ~|RG_rl_151 ;	// line#=../rle.cpp:77,78
assign	M_140 = ~|RG_rl_152 ;	// line#=../rle.cpp:77,78
assign	M_141 = ~|RG_rl_153 ;	// line#=../rle.cpp:77,78
assign	M_142 = ~|RG_rl_154 ;	// line#=../rle.cpp:77,78
assign	M_143 = ~|RG_rl_155 ;	// line#=../rle.cpp:77,78
assign	M_144 = ~|RG_rl_156 ;	// line#=../rle.cpp:77,78
assign	M_145 = ~|RG_rl_157 ;	// line#=../rle.cpp:77,78
assign	M_146 = ~|RG_rl_158 ;	// line#=../rle.cpp:77,78
assign	M_147 = ~|RG_rl_159 ;	// line#=../rle.cpp:77,78
assign	M_148 = ~|RG_rl_160 ;	// line#=../rle.cpp:77,78
assign	M_149 = ~|RG_rl_161 ;	// line#=../rle.cpp:77,78
assign	M_150 = ~|RG_rl_162 ;	// line#=../rle.cpp:77,78
assign	M_151 = ~|RG_rl_163 ;	// line#=../rle.cpp:77,78
assign	M_152 = ~|RG_rl_164 ;	// line#=../rle.cpp:77,78
assign	M_153 = ~|RG_rl_165 ;	// line#=../rle.cpp:77,78
assign	M_154 = ~|RG_rl_166 ;	// line#=../rle.cpp:77,78
assign	M_155 = ~|RG_rl_167 ;	// line#=../rle.cpp:77,78
assign	M_156 = ~|RG_rl_168 ;	// line#=../rle.cpp:77,78
assign	M_157 = ~|RG_rl_169 ;	// line#=../rle.cpp:77,78
assign	M_158 = ~|RG_rl_170 ;	// line#=../rle.cpp:77,78
assign	M_159 = ~|RG_rl_171 ;	// line#=../rle.cpp:77,78
assign	M_160 = ~|RG_rl_172 ;	// line#=../rle.cpp:77,78
assign	M_161 = ~|RG_rl_173 ;	// line#=../rle.cpp:77,78
assign	M_162 = ~|RG_rl_174 ;	// line#=../rle.cpp:77,78
assign	M_163 = ~|RG_rl_175 ;	// line#=../rle.cpp:77,78
assign	M_164 = ~|RG_rl_176 ;	// line#=../rle.cpp:77,78
assign	M_165 = ~|RG_rl_177 ;	// line#=../rle.cpp:77,78
assign	M_166 = ~|RG_rl_178 ;	// line#=../rle.cpp:77,78
assign	M_167 = ~|RG_rl_179 ;	// line#=../rle.cpp:77,78
assign	M_168 = ~|RG_rl_180 ;	// line#=../rle.cpp:77,78
assign	M_169 = ~|RG_rl_181 ;	// line#=../rle.cpp:77,78
assign	M_170 = ~|RG_rl_182 ;	// line#=../rle.cpp:77,78
assign	M_171 = ~|RG_rl_183 ;	// line#=../rle.cpp:77,78
assign	M_172 = ~|RG_rl_184 ;	// line#=../rle.cpp:77,78
assign	M_173 = ~|RG_rl_185 ;	// line#=../rle.cpp:77,78
assign	M_174 = ~|RG_rl_186 ;	// line#=../rle.cpp:77,78
assign	M_175 = ~|RG_rl_187 ;	// line#=../rle.cpp:77,78
assign	M_176 = ~|RG_rl_188 ;	// line#=../rle.cpp:77,78
assign	M_177 = ~|RG_rl_189 ;	// line#=../rle.cpp:77,78
assign	M_178 = ~|RG_rl_190 ;	// line#=../rle.cpp:77,78
assign	M_179 = ~|RG_rl_191 ;	// line#=../rle.cpp:77,78
always @ ( M_113 or M_112 or M_110 or M_179 or M_109 or M_178 or M_108 or M_177 or 
	M_107 or M_176 or M_106 or M_175 or M_105 or M_174 or M_104 or M_173 or 
	M_103 or M_172 or M_102 or M_171 or M_100 or M_170 or M_99 or M_169 or M_98 or 
	M_168 or M_97 or M_167 or M_96 or M_166 or M_95 or M_165 or M_94 or M_164 or 
	M_93 or M_163 or M_92 or M_162 or M_91 or M_161 or M_90 or M_160 or M_89 or 
	M_159 or M_88 or M_158 or M_87 or M_157 or M_86 or M_156 or M_85 or M_155 or 
	M_84 or M_154 or M_83 or M_153 or M_82 or M_152 or M_81 or M_151 or M_80 or 
	M_150 or M_79 or M_149 or M_78 or M_148 or M_77 or M_147 or M_76 or M_146 or 
	M_75 or M_145 or M_74 or M_144 or M_73 or M_143 or M_72 or M_142 or M_71 or 
	M_141 or M_70 or M_140 or M_69 or M_139 or M_68 or M_138 or M_67 or M_137 or 
	M_66 or M_136 or M_65 or M_135 or M_64 or M_134 or M_63 or M_133 or M_62 or 
	M_132 or M_61 or M_131 or M_60 or M_130 or M_59 or M_129 or M_58 or M_128 or 
	M_57 or M_127 or M_56 or M_126 or M_55 or M_125 or M_54 or M_124 or M_53 or 
	M_123 or M_52 or M_122 or M_51 or M_120 or M_50 or M_119 or M_49 or M_118 or 
	M_117 or M_116 or M_115 or M_114 or decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot )
	7'h00 :
		M_14_t128 = M_114 ;	// line#=../rle.cpp:77,78
	7'h01 :
		M_14_t128 = M_115 ;	// line#=../rle.cpp:77,78
	7'h02 :
		M_14_t128 = M_116 ;	// line#=../rle.cpp:77,78
	7'h03 :
		M_14_t128 = M_117 ;	// line#=../rle.cpp:77,78
	7'h04 :
		M_14_t128 = M_118 ;	// line#=../rle.cpp:77,78
	7'h05 :
		M_14_t128 = M_49 ;	// line#=../rle.cpp:77,78
	7'h06 :
		M_14_t128 = M_119 ;	// line#=../rle.cpp:77,78
	7'h07 :
		M_14_t128 = M_50 ;	// line#=../rle.cpp:77,78
	7'h08 :
		M_14_t128 = M_120 ;	// line#=../rle.cpp:77,78
	7'h09 :
		M_14_t128 = M_51 ;	// line#=../rle.cpp:77,78
	7'h0a :
		M_14_t128 = M_122 ;	// line#=../rle.cpp:77,78
	7'h0b :
		M_14_t128 = M_52 ;	// line#=../rle.cpp:77,78
	7'h0c :
		M_14_t128 = M_123 ;	// line#=../rle.cpp:77,78
	7'h0d :
		M_14_t128 = M_53 ;	// line#=../rle.cpp:77,78
	7'h0e :
		M_14_t128 = M_124 ;	// line#=../rle.cpp:77,78
	7'h0f :
		M_14_t128 = M_54 ;	// line#=../rle.cpp:77,78
	7'h10 :
		M_14_t128 = M_125 ;	// line#=../rle.cpp:77,78
	7'h11 :
		M_14_t128 = M_55 ;	// line#=../rle.cpp:77,78
	7'h12 :
		M_14_t128 = M_126 ;	// line#=../rle.cpp:77,78
	7'h13 :
		M_14_t128 = M_56 ;	// line#=../rle.cpp:77,78
	7'h14 :
		M_14_t128 = M_127 ;	// line#=../rle.cpp:77,78
	7'h15 :
		M_14_t128 = M_57 ;	// line#=../rle.cpp:77,78
	7'h16 :
		M_14_t128 = M_128 ;	// line#=../rle.cpp:77,78
	7'h17 :
		M_14_t128 = M_58 ;	// line#=../rle.cpp:77,78
	7'h18 :
		M_14_t128 = M_129 ;	// line#=../rle.cpp:77,78
	7'h19 :
		M_14_t128 = M_59 ;	// line#=../rle.cpp:77,78
	7'h1a :
		M_14_t128 = M_130 ;	// line#=../rle.cpp:77,78
	7'h1b :
		M_14_t128 = M_60 ;	// line#=../rle.cpp:77,78
	7'h1c :
		M_14_t128 = M_131 ;	// line#=../rle.cpp:77,78
	7'h1d :
		M_14_t128 = M_61 ;	// line#=../rle.cpp:77,78
	7'h1e :
		M_14_t128 = M_132 ;	// line#=../rle.cpp:77,78
	7'h1f :
		M_14_t128 = M_62 ;	// line#=../rle.cpp:77,78
	7'h20 :
		M_14_t128 = M_133 ;	// line#=../rle.cpp:77,78
	7'h21 :
		M_14_t128 = M_63 ;	// line#=../rle.cpp:77,78
	7'h22 :
		M_14_t128 = M_134 ;	// line#=../rle.cpp:77,78
	7'h23 :
		M_14_t128 = M_64 ;	// line#=../rle.cpp:77,78
	7'h24 :
		M_14_t128 = M_135 ;	// line#=../rle.cpp:77,78
	7'h25 :
		M_14_t128 = M_65 ;	// line#=../rle.cpp:77,78
	7'h26 :
		M_14_t128 = M_136 ;	// line#=../rle.cpp:77,78
	7'h27 :
		M_14_t128 = M_66 ;	// line#=../rle.cpp:77,78
	7'h28 :
		M_14_t128 = M_137 ;	// line#=../rle.cpp:77,78
	7'h29 :
		M_14_t128 = M_67 ;	// line#=../rle.cpp:77,78
	7'h2a :
		M_14_t128 = M_138 ;	// line#=../rle.cpp:77,78
	7'h2b :
		M_14_t128 = M_68 ;	// line#=../rle.cpp:77,78
	7'h2c :
		M_14_t128 = M_139 ;	// line#=../rle.cpp:77,78
	7'h2d :
		M_14_t128 = M_69 ;	// line#=../rle.cpp:77,78
	7'h2e :
		M_14_t128 = M_140 ;	// line#=../rle.cpp:77,78
	7'h2f :
		M_14_t128 = M_70 ;	// line#=../rle.cpp:77,78
	7'h30 :
		M_14_t128 = M_141 ;	// line#=../rle.cpp:77,78
	7'h31 :
		M_14_t128 = M_71 ;	// line#=../rle.cpp:77,78
	7'h32 :
		M_14_t128 = M_142 ;	// line#=../rle.cpp:77,78
	7'h33 :
		M_14_t128 = M_72 ;	// line#=../rle.cpp:77,78
	7'h34 :
		M_14_t128 = M_143 ;	// line#=../rle.cpp:77,78
	7'h35 :
		M_14_t128 = M_73 ;	// line#=../rle.cpp:77,78
	7'h36 :
		M_14_t128 = M_144 ;	// line#=../rle.cpp:77,78
	7'h37 :
		M_14_t128 = M_74 ;	// line#=../rle.cpp:77,78
	7'h38 :
		M_14_t128 = M_145 ;	// line#=../rle.cpp:77,78
	7'h39 :
		M_14_t128 = M_75 ;	// line#=../rle.cpp:77,78
	7'h3a :
		M_14_t128 = M_146 ;	// line#=../rle.cpp:77,78
	7'h3b :
		M_14_t128 = M_76 ;	// line#=../rle.cpp:77,78
	7'h3c :
		M_14_t128 = M_147 ;	// line#=../rle.cpp:77,78
	7'h3d :
		M_14_t128 = M_77 ;	// line#=../rle.cpp:77,78
	7'h3e :
		M_14_t128 = M_148 ;	// line#=../rle.cpp:77,78
	7'h3f :
		M_14_t128 = M_78 ;	// line#=../rle.cpp:77,78
	7'h40 :
		M_14_t128 = M_149 ;	// line#=../rle.cpp:77,78
	7'h41 :
		M_14_t128 = M_79 ;	// line#=../rle.cpp:77,78
	7'h42 :
		M_14_t128 = M_150 ;	// line#=../rle.cpp:77,78
	7'h43 :
		M_14_t128 = M_80 ;	// line#=../rle.cpp:77,78
	7'h44 :
		M_14_t128 = M_151 ;	// line#=../rle.cpp:77,78
	7'h45 :
		M_14_t128 = M_81 ;	// line#=../rle.cpp:77,78
	7'h46 :
		M_14_t128 = M_152 ;	// line#=../rle.cpp:77,78
	7'h47 :
		M_14_t128 = M_82 ;	// line#=../rle.cpp:77,78
	7'h48 :
		M_14_t128 = M_153 ;	// line#=../rle.cpp:77,78
	7'h49 :
		M_14_t128 = M_83 ;	// line#=../rle.cpp:77,78
	7'h4a :
		M_14_t128 = M_154 ;	// line#=../rle.cpp:77,78
	7'h4b :
		M_14_t128 = M_84 ;	// line#=../rle.cpp:77,78
	7'h4c :
		M_14_t128 = M_155 ;	// line#=../rle.cpp:77,78
	7'h4d :
		M_14_t128 = M_85 ;	// line#=../rle.cpp:77,78
	7'h4e :
		M_14_t128 = M_156 ;	// line#=../rle.cpp:77,78
	7'h4f :
		M_14_t128 = M_86 ;	// line#=../rle.cpp:77,78
	7'h50 :
		M_14_t128 = M_157 ;	// line#=../rle.cpp:77,78
	7'h51 :
		M_14_t128 = M_87 ;	// line#=../rle.cpp:77,78
	7'h52 :
		M_14_t128 = M_158 ;	// line#=../rle.cpp:77,78
	7'h53 :
		M_14_t128 = M_88 ;	// line#=../rle.cpp:77,78
	7'h54 :
		M_14_t128 = M_159 ;	// line#=../rle.cpp:77,78
	7'h55 :
		M_14_t128 = M_89 ;	// line#=../rle.cpp:77,78
	7'h56 :
		M_14_t128 = M_160 ;	// line#=../rle.cpp:77,78
	7'h57 :
		M_14_t128 = M_90 ;	// line#=../rle.cpp:77,78
	7'h58 :
		M_14_t128 = M_161 ;	// line#=../rle.cpp:77,78
	7'h59 :
		M_14_t128 = M_91 ;	// line#=../rle.cpp:77,78
	7'h5a :
		M_14_t128 = M_162 ;	// line#=../rle.cpp:77,78
	7'h5b :
		M_14_t128 = M_92 ;	// line#=../rle.cpp:77,78
	7'h5c :
		M_14_t128 = M_163 ;	// line#=../rle.cpp:77,78
	7'h5d :
		M_14_t128 = M_93 ;	// line#=../rle.cpp:77,78
	7'h5e :
		M_14_t128 = M_164 ;	// line#=../rle.cpp:77,78
	7'h5f :
		M_14_t128 = M_94 ;	// line#=../rle.cpp:77,78
	7'h60 :
		M_14_t128 = M_165 ;	// line#=../rle.cpp:77,78
	7'h61 :
		M_14_t128 = M_95 ;	// line#=../rle.cpp:77,78
	7'h62 :
		M_14_t128 = M_166 ;	// line#=../rle.cpp:77,78
	7'h63 :
		M_14_t128 = M_96 ;	// line#=../rle.cpp:77,78
	7'h64 :
		M_14_t128 = M_167 ;	// line#=../rle.cpp:77,78
	7'h65 :
		M_14_t128 = M_97 ;	// line#=../rle.cpp:77,78
	7'h66 :
		M_14_t128 = M_168 ;	// line#=../rle.cpp:77,78
	7'h67 :
		M_14_t128 = M_98 ;	// line#=../rle.cpp:77,78
	7'h68 :
		M_14_t128 = M_169 ;	// line#=../rle.cpp:77,78
	7'h69 :
		M_14_t128 = M_99 ;	// line#=../rle.cpp:77,78
	7'h6a :
		M_14_t128 = M_170 ;	// line#=../rle.cpp:77,78
	7'h6b :
		M_14_t128 = M_100 ;	// line#=../rle.cpp:77,78
	7'h6c :
		M_14_t128 = M_171 ;	// line#=../rle.cpp:77,78
	7'h6d :
		M_14_t128 = M_102 ;	// line#=../rle.cpp:77,78
	7'h6e :
		M_14_t128 = M_172 ;	// line#=../rle.cpp:77,78
	7'h6f :
		M_14_t128 = M_103 ;	// line#=../rle.cpp:77,78
	7'h70 :
		M_14_t128 = M_173 ;	// line#=../rle.cpp:77,78
	7'h71 :
		M_14_t128 = M_104 ;	// line#=../rle.cpp:77,78
	7'h72 :
		M_14_t128 = M_174 ;	// line#=../rle.cpp:77,78
	7'h73 :
		M_14_t128 = M_105 ;	// line#=../rle.cpp:77,78
	7'h74 :
		M_14_t128 = M_175 ;	// line#=../rle.cpp:77,78
	7'h75 :
		M_14_t128 = M_106 ;	// line#=../rle.cpp:77,78
	7'h76 :
		M_14_t128 = M_176 ;	// line#=../rle.cpp:77,78
	7'h77 :
		M_14_t128 = M_107 ;	// line#=../rle.cpp:77,78
	7'h78 :
		M_14_t128 = M_177 ;	// line#=../rle.cpp:77,78
	7'h79 :
		M_14_t128 = M_108 ;	// line#=../rle.cpp:77,78
	7'h7a :
		M_14_t128 = M_178 ;	// line#=../rle.cpp:77,78
	7'h7b :
		M_14_t128 = M_109 ;	// line#=../rle.cpp:77,78
	7'h7c :
		M_14_t128 = M_179 ;	// line#=../rle.cpp:77,78
	7'h7d :
		M_14_t128 = M_110 ;	// line#=../rle.cpp:77,78
	7'h7e :
		M_14_t128 = M_112 ;	// line#=../rle.cpp:77,78
	7'h7f :
		M_14_t128 = M_113 ;	// line#=../rle.cpp:77,78
	default :
		M_14_t128 = 1'hx ;
	endcase
always @ ( RG_previous_dc_rl or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_12 = 9'h000 ;	// line#=../rle.cpp:79
	7'h01 :
		TR_12 = RG_previous_dc_rl ;
	7'h02 :
		TR_12 = RG_previous_dc_rl ;
	7'h03 :
		TR_12 = RG_previous_dc_rl ;
	7'h04 :
		TR_12 = RG_previous_dc_rl ;
	7'h05 :
		TR_12 = RG_previous_dc_rl ;
	7'h06 :
		TR_12 = RG_previous_dc_rl ;
	7'h07 :
		TR_12 = RG_previous_dc_rl ;
	7'h08 :
		TR_12 = RG_previous_dc_rl ;
	7'h09 :
		TR_12 = RG_previous_dc_rl ;
	7'h0a :
		TR_12 = RG_previous_dc_rl ;
	7'h0b :
		TR_12 = RG_previous_dc_rl ;
	7'h0c :
		TR_12 = RG_previous_dc_rl ;
	7'h0d :
		TR_12 = RG_previous_dc_rl ;
	7'h0e :
		TR_12 = RG_previous_dc_rl ;
	7'h0f :
		TR_12 = RG_previous_dc_rl ;
	7'h10 :
		TR_12 = RG_previous_dc_rl ;
	7'h11 :
		TR_12 = RG_previous_dc_rl ;
	7'h12 :
		TR_12 = RG_previous_dc_rl ;
	7'h13 :
		TR_12 = RG_previous_dc_rl ;
	7'h14 :
		TR_12 = RG_previous_dc_rl ;
	7'h15 :
		TR_12 = RG_previous_dc_rl ;
	7'h16 :
		TR_12 = RG_previous_dc_rl ;
	7'h17 :
		TR_12 = RG_previous_dc_rl ;
	7'h18 :
		TR_12 = RG_previous_dc_rl ;
	7'h19 :
		TR_12 = RG_previous_dc_rl ;
	7'h1a :
		TR_12 = RG_previous_dc_rl ;
	7'h1b :
		TR_12 = RG_previous_dc_rl ;
	7'h1c :
		TR_12 = RG_previous_dc_rl ;
	7'h1d :
		TR_12 = RG_previous_dc_rl ;
	7'h1e :
		TR_12 = RG_previous_dc_rl ;
	7'h1f :
		TR_12 = RG_previous_dc_rl ;
	7'h20 :
		TR_12 = RG_previous_dc_rl ;
	7'h21 :
		TR_12 = RG_previous_dc_rl ;
	7'h22 :
		TR_12 = RG_previous_dc_rl ;
	7'h23 :
		TR_12 = RG_previous_dc_rl ;
	7'h24 :
		TR_12 = RG_previous_dc_rl ;
	7'h25 :
		TR_12 = RG_previous_dc_rl ;
	7'h26 :
		TR_12 = RG_previous_dc_rl ;
	7'h27 :
		TR_12 = RG_previous_dc_rl ;
	7'h28 :
		TR_12 = RG_previous_dc_rl ;
	7'h29 :
		TR_12 = RG_previous_dc_rl ;
	7'h2a :
		TR_12 = RG_previous_dc_rl ;
	7'h2b :
		TR_12 = RG_previous_dc_rl ;
	7'h2c :
		TR_12 = RG_previous_dc_rl ;
	7'h2d :
		TR_12 = RG_previous_dc_rl ;
	7'h2e :
		TR_12 = RG_previous_dc_rl ;
	7'h2f :
		TR_12 = RG_previous_dc_rl ;
	7'h30 :
		TR_12 = RG_previous_dc_rl ;
	7'h31 :
		TR_12 = RG_previous_dc_rl ;
	7'h32 :
		TR_12 = RG_previous_dc_rl ;
	7'h33 :
		TR_12 = RG_previous_dc_rl ;
	7'h34 :
		TR_12 = RG_previous_dc_rl ;
	7'h35 :
		TR_12 = RG_previous_dc_rl ;
	7'h36 :
		TR_12 = RG_previous_dc_rl ;
	7'h37 :
		TR_12 = RG_previous_dc_rl ;
	7'h38 :
		TR_12 = RG_previous_dc_rl ;
	7'h39 :
		TR_12 = RG_previous_dc_rl ;
	7'h3a :
		TR_12 = RG_previous_dc_rl ;
	7'h3b :
		TR_12 = RG_previous_dc_rl ;
	7'h3c :
		TR_12 = RG_previous_dc_rl ;
	7'h3d :
		TR_12 = RG_previous_dc_rl ;
	7'h3e :
		TR_12 = RG_previous_dc_rl ;
	7'h3f :
		TR_12 = RG_previous_dc_rl ;
	7'h40 :
		TR_12 = RG_previous_dc_rl ;
	7'h41 :
		TR_12 = RG_previous_dc_rl ;
	7'h42 :
		TR_12 = RG_previous_dc_rl ;
	7'h43 :
		TR_12 = RG_previous_dc_rl ;
	7'h44 :
		TR_12 = RG_previous_dc_rl ;
	7'h45 :
		TR_12 = RG_previous_dc_rl ;
	7'h46 :
		TR_12 = RG_previous_dc_rl ;
	7'h47 :
		TR_12 = RG_previous_dc_rl ;
	7'h48 :
		TR_12 = RG_previous_dc_rl ;
	7'h49 :
		TR_12 = RG_previous_dc_rl ;
	7'h4a :
		TR_12 = RG_previous_dc_rl ;
	7'h4b :
		TR_12 = RG_previous_dc_rl ;
	7'h4c :
		TR_12 = RG_previous_dc_rl ;
	7'h4d :
		TR_12 = RG_previous_dc_rl ;
	7'h4e :
		TR_12 = RG_previous_dc_rl ;
	7'h4f :
		TR_12 = RG_previous_dc_rl ;
	7'h50 :
		TR_12 = RG_previous_dc_rl ;
	7'h51 :
		TR_12 = RG_previous_dc_rl ;
	7'h52 :
		TR_12 = RG_previous_dc_rl ;
	7'h53 :
		TR_12 = RG_previous_dc_rl ;
	7'h54 :
		TR_12 = RG_previous_dc_rl ;
	7'h55 :
		TR_12 = RG_previous_dc_rl ;
	7'h56 :
		TR_12 = RG_previous_dc_rl ;
	7'h57 :
		TR_12 = RG_previous_dc_rl ;
	7'h58 :
		TR_12 = RG_previous_dc_rl ;
	7'h59 :
		TR_12 = RG_previous_dc_rl ;
	7'h5a :
		TR_12 = RG_previous_dc_rl ;
	7'h5b :
		TR_12 = RG_previous_dc_rl ;
	7'h5c :
		TR_12 = RG_previous_dc_rl ;
	7'h5d :
		TR_12 = RG_previous_dc_rl ;
	7'h5e :
		TR_12 = RG_previous_dc_rl ;
	7'h5f :
		TR_12 = RG_previous_dc_rl ;
	7'h60 :
		TR_12 = RG_previous_dc_rl ;
	7'h61 :
		TR_12 = RG_previous_dc_rl ;
	7'h62 :
		TR_12 = RG_previous_dc_rl ;
	7'h63 :
		TR_12 = RG_previous_dc_rl ;
	7'h64 :
		TR_12 = RG_previous_dc_rl ;
	7'h65 :
		TR_12 = RG_previous_dc_rl ;
	7'h66 :
		TR_12 = RG_previous_dc_rl ;
	7'h67 :
		TR_12 = RG_previous_dc_rl ;
	7'h68 :
		TR_12 = RG_previous_dc_rl ;
	7'h69 :
		TR_12 = RG_previous_dc_rl ;
	7'h6a :
		TR_12 = RG_previous_dc_rl ;
	7'h6b :
		TR_12 = RG_previous_dc_rl ;
	7'h6c :
		TR_12 = RG_previous_dc_rl ;
	7'h6d :
		TR_12 = RG_previous_dc_rl ;
	7'h6e :
		TR_12 = RG_previous_dc_rl ;
	7'h6f :
		TR_12 = RG_previous_dc_rl ;
	7'h70 :
		TR_12 = RG_previous_dc_rl ;
	7'h71 :
		TR_12 = RG_previous_dc_rl ;
	7'h72 :
		TR_12 = RG_previous_dc_rl ;
	7'h73 :
		TR_12 = RG_previous_dc_rl ;
	7'h74 :
		TR_12 = RG_previous_dc_rl ;
	7'h75 :
		TR_12 = RG_previous_dc_rl ;
	7'h76 :
		TR_12 = RG_previous_dc_rl ;
	7'h77 :
		TR_12 = RG_previous_dc_rl ;
	7'h78 :
		TR_12 = RG_previous_dc_rl ;
	7'h79 :
		TR_12 = RG_previous_dc_rl ;
	7'h7a :
		TR_12 = RG_previous_dc_rl ;
	7'h7b :
		TR_12 = RG_previous_dc_rl ;
	7'h7c :
		TR_12 = RG_previous_dc_rl ;
	7'h7d :
		TR_12 = RG_previous_dc_rl ;
	7'h7e :
		TR_12 = RG_previous_dc_rl ;
	7'h7f :
		TR_12 = RG_previous_dc_rl ;
	default :
		TR_12 = 9'hx ;
	endcase
always @ ( RG_rl_128 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_13 = RG_rl_128 ;
	7'h01 :
		TR_13 = 9'h000 ;	// line#=../rle.cpp:79
	7'h02 :
		TR_13 = RG_rl_128 ;
	7'h03 :
		TR_13 = RG_rl_128 ;
	7'h04 :
		TR_13 = RG_rl_128 ;
	7'h05 :
		TR_13 = RG_rl_128 ;
	7'h06 :
		TR_13 = RG_rl_128 ;
	7'h07 :
		TR_13 = RG_rl_128 ;
	7'h08 :
		TR_13 = RG_rl_128 ;
	7'h09 :
		TR_13 = RG_rl_128 ;
	7'h0a :
		TR_13 = RG_rl_128 ;
	7'h0b :
		TR_13 = RG_rl_128 ;
	7'h0c :
		TR_13 = RG_rl_128 ;
	7'h0d :
		TR_13 = RG_rl_128 ;
	7'h0e :
		TR_13 = RG_rl_128 ;
	7'h0f :
		TR_13 = RG_rl_128 ;
	7'h10 :
		TR_13 = RG_rl_128 ;
	7'h11 :
		TR_13 = RG_rl_128 ;
	7'h12 :
		TR_13 = RG_rl_128 ;
	7'h13 :
		TR_13 = RG_rl_128 ;
	7'h14 :
		TR_13 = RG_rl_128 ;
	7'h15 :
		TR_13 = RG_rl_128 ;
	7'h16 :
		TR_13 = RG_rl_128 ;
	7'h17 :
		TR_13 = RG_rl_128 ;
	7'h18 :
		TR_13 = RG_rl_128 ;
	7'h19 :
		TR_13 = RG_rl_128 ;
	7'h1a :
		TR_13 = RG_rl_128 ;
	7'h1b :
		TR_13 = RG_rl_128 ;
	7'h1c :
		TR_13 = RG_rl_128 ;
	7'h1d :
		TR_13 = RG_rl_128 ;
	7'h1e :
		TR_13 = RG_rl_128 ;
	7'h1f :
		TR_13 = RG_rl_128 ;
	7'h20 :
		TR_13 = RG_rl_128 ;
	7'h21 :
		TR_13 = RG_rl_128 ;
	7'h22 :
		TR_13 = RG_rl_128 ;
	7'h23 :
		TR_13 = RG_rl_128 ;
	7'h24 :
		TR_13 = RG_rl_128 ;
	7'h25 :
		TR_13 = RG_rl_128 ;
	7'h26 :
		TR_13 = RG_rl_128 ;
	7'h27 :
		TR_13 = RG_rl_128 ;
	7'h28 :
		TR_13 = RG_rl_128 ;
	7'h29 :
		TR_13 = RG_rl_128 ;
	7'h2a :
		TR_13 = RG_rl_128 ;
	7'h2b :
		TR_13 = RG_rl_128 ;
	7'h2c :
		TR_13 = RG_rl_128 ;
	7'h2d :
		TR_13 = RG_rl_128 ;
	7'h2e :
		TR_13 = RG_rl_128 ;
	7'h2f :
		TR_13 = RG_rl_128 ;
	7'h30 :
		TR_13 = RG_rl_128 ;
	7'h31 :
		TR_13 = RG_rl_128 ;
	7'h32 :
		TR_13 = RG_rl_128 ;
	7'h33 :
		TR_13 = RG_rl_128 ;
	7'h34 :
		TR_13 = RG_rl_128 ;
	7'h35 :
		TR_13 = RG_rl_128 ;
	7'h36 :
		TR_13 = RG_rl_128 ;
	7'h37 :
		TR_13 = RG_rl_128 ;
	7'h38 :
		TR_13 = RG_rl_128 ;
	7'h39 :
		TR_13 = RG_rl_128 ;
	7'h3a :
		TR_13 = RG_rl_128 ;
	7'h3b :
		TR_13 = RG_rl_128 ;
	7'h3c :
		TR_13 = RG_rl_128 ;
	7'h3d :
		TR_13 = RG_rl_128 ;
	7'h3e :
		TR_13 = RG_rl_128 ;
	7'h3f :
		TR_13 = RG_rl_128 ;
	7'h40 :
		TR_13 = RG_rl_128 ;
	7'h41 :
		TR_13 = RG_rl_128 ;
	7'h42 :
		TR_13 = RG_rl_128 ;
	7'h43 :
		TR_13 = RG_rl_128 ;
	7'h44 :
		TR_13 = RG_rl_128 ;
	7'h45 :
		TR_13 = RG_rl_128 ;
	7'h46 :
		TR_13 = RG_rl_128 ;
	7'h47 :
		TR_13 = RG_rl_128 ;
	7'h48 :
		TR_13 = RG_rl_128 ;
	7'h49 :
		TR_13 = RG_rl_128 ;
	7'h4a :
		TR_13 = RG_rl_128 ;
	7'h4b :
		TR_13 = RG_rl_128 ;
	7'h4c :
		TR_13 = RG_rl_128 ;
	7'h4d :
		TR_13 = RG_rl_128 ;
	7'h4e :
		TR_13 = RG_rl_128 ;
	7'h4f :
		TR_13 = RG_rl_128 ;
	7'h50 :
		TR_13 = RG_rl_128 ;
	7'h51 :
		TR_13 = RG_rl_128 ;
	7'h52 :
		TR_13 = RG_rl_128 ;
	7'h53 :
		TR_13 = RG_rl_128 ;
	7'h54 :
		TR_13 = RG_rl_128 ;
	7'h55 :
		TR_13 = RG_rl_128 ;
	7'h56 :
		TR_13 = RG_rl_128 ;
	7'h57 :
		TR_13 = RG_rl_128 ;
	7'h58 :
		TR_13 = RG_rl_128 ;
	7'h59 :
		TR_13 = RG_rl_128 ;
	7'h5a :
		TR_13 = RG_rl_128 ;
	7'h5b :
		TR_13 = RG_rl_128 ;
	7'h5c :
		TR_13 = RG_rl_128 ;
	7'h5d :
		TR_13 = RG_rl_128 ;
	7'h5e :
		TR_13 = RG_rl_128 ;
	7'h5f :
		TR_13 = RG_rl_128 ;
	7'h60 :
		TR_13 = RG_rl_128 ;
	7'h61 :
		TR_13 = RG_rl_128 ;
	7'h62 :
		TR_13 = RG_rl_128 ;
	7'h63 :
		TR_13 = RG_rl_128 ;
	7'h64 :
		TR_13 = RG_rl_128 ;
	7'h65 :
		TR_13 = RG_rl_128 ;
	7'h66 :
		TR_13 = RG_rl_128 ;
	7'h67 :
		TR_13 = RG_rl_128 ;
	7'h68 :
		TR_13 = RG_rl_128 ;
	7'h69 :
		TR_13 = RG_rl_128 ;
	7'h6a :
		TR_13 = RG_rl_128 ;
	7'h6b :
		TR_13 = RG_rl_128 ;
	7'h6c :
		TR_13 = RG_rl_128 ;
	7'h6d :
		TR_13 = RG_rl_128 ;
	7'h6e :
		TR_13 = RG_rl_128 ;
	7'h6f :
		TR_13 = RG_rl_128 ;
	7'h70 :
		TR_13 = RG_rl_128 ;
	7'h71 :
		TR_13 = RG_rl_128 ;
	7'h72 :
		TR_13 = RG_rl_128 ;
	7'h73 :
		TR_13 = RG_rl_128 ;
	7'h74 :
		TR_13 = RG_rl_128 ;
	7'h75 :
		TR_13 = RG_rl_128 ;
	7'h76 :
		TR_13 = RG_rl_128 ;
	7'h77 :
		TR_13 = RG_rl_128 ;
	7'h78 :
		TR_13 = RG_rl_128 ;
	7'h79 :
		TR_13 = RG_rl_128 ;
	7'h7a :
		TR_13 = RG_rl_128 ;
	7'h7b :
		TR_13 = RG_rl_128 ;
	7'h7c :
		TR_13 = RG_rl_128 ;
	7'h7d :
		TR_13 = RG_rl_128 ;
	7'h7e :
		TR_13 = RG_rl_128 ;
	7'h7f :
		TR_13 = RG_rl_128 ;
	default :
		TR_13 = 9'hx ;
	endcase
always @ ( RG_rl_129 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_14 = RG_rl_129 ;
	7'h01 :
		TR_14 = RG_rl_129 ;
	7'h02 :
		TR_14 = 9'h000 ;	// line#=../rle.cpp:79
	7'h03 :
		TR_14 = RG_rl_129 ;
	7'h04 :
		TR_14 = RG_rl_129 ;
	7'h05 :
		TR_14 = RG_rl_129 ;
	7'h06 :
		TR_14 = RG_rl_129 ;
	7'h07 :
		TR_14 = RG_rl_129 ;
	7'h08 :
		TR_14 = RG_rl_129 ;
	7'h09 :
		TR_14 = RG_rl_129 ;
	7'h0a :
		TR_14 = RG_rl_129 ;
	7'h0b :
		TR_14 = RG_rl_129 ;
	7'h0c :
		TR_14 = RG_rl_129 ;
	7'h0d :
		TR_14 = RG_rl_129 ;
	7'h0e :
		TR_14 = RG_rl_129 ;
	7'h0f :
		TR_14 = RG_rl_129 ;
	7'h10 :
		TR_14 = RG_rl_129 ;
	7'h11 :
		TR_14 = RG_rl_129 ;
	7'h12 :
		TR_14 = RG_rl_129 ;
	7'h13 :
		TR_14 = RG_rl_129 ;
	7'h14 :
		TR_14 = RG_rl_129 ;
	7'h15 :
		TR_14 = RG_rl_129 ;
	7'h16 :
		TR_14 = RG_rl_129 ;
	7'h17 :
		TR_14 = RG_rl_129 ;
	7'h18 :
		TR_14 = RG_rl_129 ;
	7'h19 :
		TR_14 = RG_rl_129 ;
	7'h1a :
		TR_14 = RG_rl_129 ;
	7'h1b :
		TR_14 = RG_rl_129 ;
	7'h1c :
		TR_14 = RG_rl_129 ;
	7'h1d :
		TR_14 = RG_rl_129 ;
	7'h1e :
		TR_14 = RG_rl_129 ;
	7'h1f :
		TR_14 = RG_rl_129 ;
	7'h20 :
		TR_14 = RG_rl_129 ;
	7'h21 :
		TR_14 = RG_rl_129 ;
	7'h22 :
		TR_14 = RG_rl_129 ;
	7'h23 :
		TR_14 = RG_rl_129 ;
	7'h24 :
		TR_14 = RG_rl_129 ;
	7'h25 :
		TR_14 = RG_rl_129 ;
	7'h26 :
		TR_14 = RG_rl_129 ;
	7'h27 :
		TR_14 = RG_rl_129 ;
	7'h28 :
		TR_14 = RG_rl_129 ;
	7'h29 :
		TR_14 = RG_rl_129 ;
	7'h2a :
		TR_14 = RG_rl_129 ;
	7'h2b :
		TR_14 = RG_rl_129 ;
	7'h2c :
		TR_14 = RG_rl_129 ;
	7'h2d :
		TR_14 = RG_rl_129 ;
	7'h2e :
		TR_14 = RG_rl_129 ;
	7'h2f :
		TR_14 = RG_rl_129 ;
	7'h30 :
		TR_14 = RG_rl_129 ;
	7'h31 :
		TR_14 = RG_rl_129 ;
	7'h32 :
		TR_14 = RG_rl_129 ;
	7'h33 :
		TR_14 = RG_rl_129 ;
	7'h34 :
		TR_14 = RG_rl_129 ;
	7'h35 :
		TR_14 = RG_rl_129 ;
	7'h36 :
		TR_14 = RG_rl_129 ;
	7'h37 :
		TR_14 = RG_rl_129 ;
	7'h38 :
		TR_14 = RG_rl_129 ;
	7'h39 :
		TR_14 = RG_rl_129 ;
	7'h3a :
		TR_14 = RG_rl_129 ;
	7'h3b :
		TR_14 = RG_rl_129 ;
	7'h3c :
		TR_14 = RG_rl_129 ;
	7'h3d :
		TR_14 = RG_rl_129 ;
	7'h3e :
		TR_14 = RG_rl_129 ;
	7'h3f :
		TR_14 = RG_rl_129 ;
	7'h40 :
		TR_14 = RG_rl_129 ;
	7'h41 :
		TR_14 = RG_rl_129 ;
	7'h42 :
		TR_14 = RG_rl_129 ;
	7'h43 :
		TR_14 = RG_rl_129 ;
	7'h44 :
		TR_14 = RG_rl_129 ;
	7'h45 :
		TR_14 = RG_rl_129 ;
	7'h46 :
		TR_14 = RG_rl_129 ;
	7'h47 :
		TR_14 = RG_rl_129 ;
	7'h48 :
		TR_14 = RG_rl_129 ;
	7'h49 :
		TR_14 = RG_rl_129 ;
	7'h4a :
		TR_14 = RG_rl_129 ;
	7'h4b :
		TR_14 = RG_rl_129 ;
	7'h4c :
		TR_14 = RG_rl_129 ;
	7'h4d :
		TR_14 = RG_rl_129 ;
	7'h4e :
		TR_14 = RG_rl_129 ;
	7'h4f :
		TR_14 = RG_rl_129 ;
	7'h50 :
		TR_14 = RG_rl_129 ;
	7'h51 :
		TR_14 = RG_rl_129 ;
	7'h52 :
		TR_14 = RG_rl_129 ;
	7'h53 :
		TR_14 = RG_rl_129 ;
	7'h54 :
		TR_14 = RG_rl_129 ;
	7'h55 :
		TR_14 = RG_rl_129 ;
	7'h56 :
		TR_14 = RG_rl_129 ;
	7'h57 :
		TR_14 = RG_rl_129 ;
	7'h58 :
		TR_14 = RG_rl_129 ;
	7'h59 :
		TR_14 = RG_rl_129 ;
	7'h5a :
		TR_14 = RG_rl_129 ;
	7'h5b :
		TR_14 = RG_rl_129 ;
	7'h5c :
		TR_14 = RG_rl_129 ;
	7'h5d :
		TR_14 = RG_rl_129 ;
	7'h5e :
		TR_14 = RG_rl_129 ;
	7'h5f :
		TR_14 = RG_rl_129 ;
	7'h60 :
		TR_14 = RG_rl_129 ;
	7'h61 :
		TR_14 = RG_rl_129 ;
	7'h62 :
		TR_14 = RG_rl_129 ;
	7'h63 :
		TR_14 = RG_rl_129 ;
	7'h64 :
		TR_14 = RG_rl_129 ;
	7'h65 :
		TR_14 = RG_rl_129 ;
	7'h66 :
		TR_14 = RG_rl_129 ;
	7'h67 :
		TR_14 = RG_rl_129 ;
	7'h68 :
		TR_14 = RG_rl_129 ;
	7'h69 :
		TR_14 = RG_rl_129 ;
	7'h6a :
		TR_14 = RG_rl_129 ;
	7'h6b :
		TR_14 = RG_rl_129 ;
	7'h6c :
		TR_14 = RG_rl_129 ;
	7'h6d :
		TR_14 = RG_rl_129 ;
	7'h6e :
		TR_14 = RG_rl_129 ;
	7'h6f :
		TR_14 = RG_rl_129 ;
	7'h70 :
		TR_14 = RG_rl_129 ;
	7'h71 :
		TR_14 = RG_rl_129 ;
	7'h72 :
		TR_14 = RG_rl_129 ;
	7'h73 :
		TR_14 = RG_rl_129 ;
	7'h74 :
		TR_14 = RG_rl_129 ;
	7'h75 :
		TR_14 = RG_rl_129 ;
	7'h76 :
		TR_14 = RG_rl_129 ;
	7'h77 :
		TR_14 = RG_rl_129 ;
	7'h78 :
		TR_14 = RG_rl_129 ;
	7'h79 :
		TR_14 = RG_rl_129 ;
	7'h7a :
		TR_14 = RG_rl_129 ;
	7'h7b :
		TR_14 = RG_rl_129 ;
	7'h7c :
		TR_14 = RG_rl_129 ;
	7'h7d :
		TR_14 = RG_rl_129 ;
	7'h7e :
		TR_14 = RG_rl_129 ;
	7'h7f :
		TR_14 = RG_rl_129 ;
	default :
		TR_14 = 9'hx ;
	endcase
always @ ( RG_rl_130 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_15 = RG_rl_130 ;
	7'h01 :
		TR_15 = RG_rl_130 ;
	7'h02 :
		TR_15 = RG_rl_130 ;
	7'h03 :
		TR_15 = 9'h000 ;	// line#=../rle.cpp:79
	7'h04 :
		TR_15 = RG_rl_130 ;
	7'h05 :
		TR_15 = RG_rl_130 ;
	7'h06 :
		TR_15 = RG_rl_130 ;
	7'h07 :
		TR_15 = RG_rl_130 ;
	7'h08 :
		TR_15 = RG_rl_130 ;
	7'h09 :
		TR_15 = RG_rl_130 ;
	7'h0a :
		TR_15 = RG_rl_130 ;
	7'h0b :
		TR_15 = RG_rl_130 ;
	7'h0c :
		TR_15 = RG_rl_130 ;
	7'h0d :
		TR_15 = RG_rl_130 ;
	7'h0e :
		TR_15 = RG_rl_130 ;
	7'h0f :
		TR_15 = RG_rl_130 ;
	7'h10 :
		TR_15 = RG_rl_130 ;
	7'h11 :
		TR_15 = RG_rl_130 ;
	7'h12 :
		TR_15 = RG_rl_130 ;
	7'h13 :
		TR_15 = RG_rl_130 ;
	7'h14 :
		TR_15 = RG_rl_130 ;
	7'h15 :
		TR_15 = RG_rl_130 ;
	7'h16 :
		TR_15 = RG_rl_130 ;
	7'h17 :
		TR_15 = RG_rl_130 ;
	7'h18 :
		TR_15 = RG_rl_130 ;
	7'h19 :
		TR_15 = RG_rl_130 ;
	7'h1a :
		TR_15 = RG_rl_130 ;
	7'h1b :
		TR_15 = RG_rl_130 ;
	7'h1c :
		TR_15 = RG_rl_130 ;
	7'h1d :
		TR_15 = RG_rl_130 ;
	7'h1e :
		TR_15 = RG_rl_130 ;
	7'h1f :
		TR_15 = RG_rl_130 ;
	7'h20 :
		TR_15 = RG_rl_130 ;
	7'h21 :
		TR_15 = RG_rl_130 ;
	7'h22 :
		TR_15 = RG_rl_130 ;
	7'h23 :
		TR_15 = RG_rl_130 ;
	7'h24 :
		TR_15 = RG_rl_130 ;
	7'h25 :
		TR_15 = RG_rl_130 ;
	7'h26 :
		TR_15 = RG_rl_130 ;
	7'h27 :
		TR_15 = RG_rl_130 ;
	7'h28 :
		TR_15 = RG_rl_130 ;
	7'h29 :
		TR_15 = RG_rl_130 ;
	7'h2a :
		TR_15 = RG_rl_130 ;
	7'h2b :
		TR_15 = RG_rl_130 ;
	7'h2c :
		TR_15 = RG_rl_130 ;
	7'h2d :
		TR_15 = RG_rl_130 ;
	7'h2e :
		TR_15 = RG_rl_130 ;
	7'h2f :
		TR_15 = RG_rl_130 ;
	7'h30 :
		TR_15 = RG_rl_130 ;
	7'h31 :
		TR_15 = RG_rl_130 ;
	7'h32 :
		TR_15 = RG_rl_130 ;
	7'h33 :
		TR_15 = RG_rl_130 ;
	7'h34 :
		TR_15 = RG_rl_130 ;
	7'h35 :
		TR_15 = RG_rl_130 ;
	7'h36 :
		TR_15 = RG_rl_130 ;
	7'h37 :
		TR_15 = RG_rl_130 ;
	7'h38 :
		TR_15 = RG_rl_130 ;
	7'h39 :
		TR_15 = RG_rl_130 ;
	7'h3a :
		TR_15 = RG_rl_130 ;
	7'h3b :
		TR_15 = RG_rl_130 ;
	7'h3c :
		TR_15 = RG_rl_130 ;
	7'h3d :
		TR_15 = RG_rl_130 ;
	7'h3e :
		TR_15 = RG_rl_130 ;
	7'h3f :
		TR_15 = RG_rl_130 ;
	7'h40 :
		TR_15 = RG_rl_130 ;
	7'h41 :
		TR_15 = RG_rl_130 ;
	7'h42 :
		TR_15 = RG_rl_130 ;
	7'h43 :
		TR_15 = RG_rl_130 ;
	7'h44 :
		TR_15 = RG_rl_130 ;
	7'h45 :
		TR_15 = RG_rl_130 ;
	7'h46 :
		TR_15 = RG_rl_130 ;
	7'h47 :
		TR_15 = RG_rl_130 ;
	7'h48 :
		TR_15 = RG_rl_130 ;
	7'h49 :
		TR_15 = RG_rl_130 ;
	7'h4a :
		TR_15 = RG_rl_130 ;
	7'h4b :
		TR_15 = RG_rl_130 ;
	7'h4c :
		TR_15 = RG_rl_130 ;
	7'h4d :
		TR_15 = RG_rl_130 ;
	7'h4e :
		TR_15 = RG_rl_130 ;
	7'h4f :
		TR_15 = RG_rl_130 ;
	7'h50 :
		TR_15 = RG_rl_130 ;
	7'h51 :
		TR_15 = RG_rl_130 ;
	7'h52 :
		TR_15 = RG_rl_130 ;
	7'h53 :
		TR_15 = RG_rl_130 ;
	7'h54 :
		TR_15 = RG_rl_130 ;
	7'h55 :
		TR_15 = RG_rl_130 ;
	7'h56 :
		TR_15 = RG_rl_130 ;
	7'h57 :
		TR_15 = RG_rl_130 ;
	7'h58 :
		TR_15 = RG_rl_130 ;
	7'h59 :
		TR_15 = RG_rl_130 ;
	7'h5a :
		TR_15 = RG_rl_130 ;
	7'h5b :
		TR_15 = RG_rl_130 ;
	7'h5c :
		TR_15 = RG_rl_130 ;
	7'h5d :
		TR_15 = RG_rl_130 ;
	7'h5e :
		TR_15 = RG_rl_130 ;
	7'h5f :
		TR_15 = RG_rl_130 ;
	7'h60 :
		TR_15 = RG_rl_130 ;
	7'h61 :
		TR_15 = RG_rl_130 ;
	7'h62 :
		TR_15 = RG_rl_130 ;
	7'h63 :
		TR_15 = RG_rl_130 ;
	7'h64 :
		TR_15 = RG_rl_130 ;
	7'h65 :
		TR_15 = RG_rl_130 ;
	7'h66 :
		TR_15 = RG_rl_130 ;
	7'h67 :
		TR_15 = RG_rl_130 ;
	7'h68 :
		TR_15 = RG_rl_130 ;
	7'h69 :
		TR_15 = RG_rl_130 ;
	7'h6a :
		TR_15 = RG_rl_130 ;
	7'h6b :
		TR_15 = RG_rl_130 ;
	7'h6c :
		TR_15 = RG_rl_130 ;
	7'h6d :
		TR_15 = RG_rl_130 ;
	7'h6e :
		TR_15 = RG_rl_130 ;
	7'h6f :
		TR_15 = RG_rl_130 ;
	7'h70 :
		TR_15 = RG_rl_130 ;
	7'h71 :
		TR_15 = RG_rl_130 ;
	7'h72 :
		TR_15 = RG_rl_130 ;
	7'h73 :
		TR_15 = RG_rl_130 ;
	7'h74 :
		TR_15 = RG_rl_130 ;
	7'h75 :
		TR_15 = RG_rl_130 ;
	7'h76 :
		TR_15 = RG_rl_130 ;
	7'h77 :
		TR_15 = RG_rl_130 ;
	7'h78 :
		TR_15 = RG_rl_130 ;
	7'h79 :
		TR_15 = RG_rl_130 ;
	7'h7a :
		TR_15 = RG_rl_130 ;
	7'h7b :
		TR_15 = RG_rl_130 ;
	7'h7c :
		TR_15 = RG_rl_130 ;
	7'h7d :
		TR_15 = RG_rl_130 ;
	7'h7e :
		TR_15 = RG_rl_130 ;
	7'h7f :
		TR_15 = RG_rl_130 ;
	default :
		TR_15 = 9'hx ;
	endcase
always @ ( RG_rl_131 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_16 = RG_rl_131 ;
	7'h01 :
		TR_16 = RG_rl_131 ;
	7'h02 :
		TR_16 = RG_rl_131 ;
	7'h03 :
		TR_16 = RG_rl_131 ;
	7'h04 :
		TR_16 = 9'h000 ;	// line#=../rle.cpp:79
	7'h05 :
		TR_16 = RG_rl_131 ;
	7'h06 :
		TR_16 = RG_rl_131 ;
	7'h07 :
		TR_16 = RG_rl_131 ;
	7'h08 :
		TR_16 = RG_rl_131 ;
	7'h09 :
		TR_16 = RG_rl_131 ;
	7'h0a :
		TR_16 = RG_rl_131 ;
	7'h0b :
		TR_16 = RG_rl_131 ;
	7'h0c :
		TR_16 = RG_rl_131 ;
	7'h0d :
		TR_16 = RG_rl_131 ;
	7'h0e :
		TR_16 = RG_rl_131 ;
	7'h0f :
		TR_16 = RG_rl_131 ;
	7'h10 :
		TR_16 = RG_rl_131 ;
	7'h11 :
		TR_16 = RG_rl_131 ;
	7'h12 :
		TR_16 = RG_rl_131 ;
	7'h13 :
		TR_16 = RG_rl_131 ;
	7'h14 :
		TR_16 = RG_rl_131 ;
	7'h15 :
		TR_16 = RG_rl_131 ;
	7'h16 :
		TR_16 = RG_rl_131 ;
	7'h17 :
		TR_16 = RG_rl_131 ;
	7'h18 :
		TR_16 = RG_rl_131 ;
	7'h19 :
		TR_16 = RG_rl_131 ;
	7'h1a :
		TR_16 = RG_rl_131 ;
	7'h1b :
		TR_16 = RG_rl_131 ;
	7'h1c :
		TR_16 = RG_rl_131 ;
	7'h1d :
		TR_16 = RG_rl_131 ;
	7'h1e :
		TR_16 = RG_rl_131 ;
	7'h1f :
		TR_16 = RG_rl_131 ;
	7'h20 :
		TR_16 = RG_rl_131 ;
	7'h21 :
		TR_16 = RG_rl_131 ;
	7'h22 :
		TR_16 = RG_rl_131 ;
	7'h23 :
		TR_16 = RG_rl_131 ;
	7'h24 :
		TR_16 = RG_rl_131 ;
	7'h25 :
		TR_16 = RG_rl_131 ;
	7'h26 :
		TR_16 = RG_rl_131 ;
	7'h27 :
		TR_16 = RG_rl_131 ;
	7'h28 :
		TR_16 = RG_rl_131 ;
	7'h29 :
		TR_16 = RG_rl_131 ;
	7'h2a :
		TR_16 = RG_rl_131 ;
	7'h2b :
		TR_16 = RG_rl_131 ;
	7'h2c :
		TR_16 = RG_rl_131 ;
	7'h2d :
		TR_16 = RG_rl_131 ;
	7'h2e :
		TR_16 = RG_rl_131 ;
	7'h2f :
		TR_16 = RG_rl_131 ;
	7'h30 :
		TR_16 = RG_rl_131 ;
	7'h31 :
		TR_16 = RG_rl_131 ;
	7'h32 :
		TR_16 = RG_rl_131 ;
	7'h33 :
		TR_16 = RG_rl_131 ;
	7'h34 :
		TR_16 = RG_rl_131 ;
	7'h35 :
		TR_16 = RG_rl_131 ;
	7'h36 :
		TR_16 = RG_rl_131 ;
	7'h37 :
		TR_16 = RG_rl_131 ;
	7'h38 :
		TR_16 = RG_rl_131 ;
	7'h39 :
		TR_16 = RG_rl_131 ;
	7'h3a :
		TR_16 = RG_rl_131 ;
	7'h3b :
		TR_16 = RG_rl_131 ;
	7'h3c :
		TR_16 = RG_rl_131 ;
	7'h3d :
		TR_16 = RG_rl_131 ;
	7'h3e :
		TR_16 = RG_rl_131 ;
	7'h3f :
		TR_16 = RG_rl_131 ;
	7'h40 :
		TR_16 = RG_rl_131 ;
	7'h41 :
		TR_16 = RG_rl_131 ;
	7'h42 :
		TR_16 = RG_rl_131 ;
	7'h43 :
		TR_16 = RG_rl_131 ;
	7'h44 :
		TR_16 = RG_rl_131 ;
	7'h45 :
		TR_16 = RG_rl_131 ;
	7'h46 :
		TR_16 = RG_rl_131 ;
	7'h47 :
		TR_16 = RG_rl_131 ;
	7'h48 :
		TR_16 = RG_rl_131 ;
	7'h49 :
		TR_16 = RG_rl_131 ;
	7'h4a :
		TR_16 = RG_rl_131 ;
	7'h4b :
		TR_16 = RG_rl_131 ;
	7'h4c :
		TR_16 = RG_rl_131 ;
	7'h4d :
		TR_16 = RG_rl_131 ;
	7'h4e :
		TR_16 = RG_rl_131 ;
	7'h4f :
		TR_16 = RG_rl_131 ;
	7'h50 :
		TR_16 = RG_rl_131 ;
	7'h51 :
		TR_16 = RG_rl_131 ;
	7'h52 :
		TR_16 = RG_rl_131 ;
	7'h53 :
		TR_16 = RG_rl_131 ;
	7'h54 :
		TR_16 = RG_rl_131 ;
	7'h55 :
		TR_16 = RG_rl_131 ;
	7'h56 :
		TR_16 = RG_rl_131 ;
	7'h57 :
		TR_16 = RG_rl_131 ;
	7'h58 :
		TR_16 = RG_rl_131 ;
	7'h59 :
		TR_16 = RG_rl_131 ;
	7'h5a :
		TR_16 = RG_rl_131 ;
	7'h5b :
		TR_16 = RG_rl_131 ;
	7'h5c :
		TR_16 = RG_rl_131 ;
	7'h5d :
		TR_16 = RG_rl_131 ;
	7'h5e :
		TR_16 = RG_rl_131 ;
	7'h5f :
		TR_16 = RG_rl_131 ;
	7'h60 :
		TR_16 = RG_rl_131 ;
	7'h61 :
		TR_16 = RG_rl_131 ;
	7'h62 :
		TR_16 = RG_rl_131 ;
	7'h63 :
		TR_16 = RG_rl_131 ;
	7'h64 :
		TR_16 = RG_rl_131 ;
	7'h65 :
		TR_16 = RG_rl_131 ;
	7'h66 :
		TR_16 = RG_rl_131 ;
	7'h67 :
		TR_16 = RG_rl_131 ;
	7'h68 :
		TR_16 = RG_rl_131 ;
	7'h69 :
		TR_16 = RG_rl_131 ;
	7'h6a :
		TR_16 = RG_rl_131 ;
	7'h6b :
		TR_16 = RG_rl_131 ;
	7'h6c :
		TR_16 = RG_rl_131 ;
	7'h6d :
		TR_16 = RG_rl_131 ;
	7'h6e :
		TR_16 = RG_rl_131 ;
	7'h6f :
		TR_16 = RG_rl_131 ;
	7'h70 :
		TR_16 = RG_rl_131 ;
	7'h71 :
		TR_16 = RG_rl_131 ;
	7'h72 :
		TR_16 = RG_rl_131 ;
	7'h73 :
		TR_16 = RG_rl_131 ;
	7'h74 :
		TR_16 = RG_rl_131 ;
	7'h75 :
		TR_16 = RG_rl_131 ;
	7'h76 :
		TR_16 = RG_rl_131 ;
	7'h77 :
		TR_16 = RG_rl_131 ;
	7'h78 :
		TR_16 = RG_rl_131 ;
	7'h79 :
		TR_16 = RG_rl_131 ;
	7'h7a :
		TR_16 = RG_rl_131 ;
	7'h7b :
		TR_16 = RG_rl_131 ;
	7'h7c :
		TR_16 = RG_rl_131 ;
	7'h7d :
		TR_16 = RG_rl_131 ;
	7'h7e :
		TR_16 = RG_rl_131 ;
	7'h7f :
		TR_16 = RG_rl_131 ;
	default :
		TR_16 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_17 = RG_quantized_block_rl ;
	7'h01 :
		TR_17 = RG_quantized_block_rl ;
	7'h02 :
		TR_17 = RG_quantized_block_rl ;
	7'h03 :
		TR_17 = RG_quantized_block_rl ;
	7'h04 :
		TR_17 = RG_quantized_block_rl ;
	7'h05 :
		TR_17 = 9'h000 ;	// line#=../rle.cpp:79
	7'h06 :
		TR_17 = RG_quantized_block_rl ;
	7'h07 :
		TR_17 = RG_quantized_block_rl ;
	7'h08 :
		TR_17 = RG_quantized_block_rl ;
	7'h09 :
		TR_17 = RG_quantized_block_rl ;
	7'h0a :
		TR_17 = RG_quantized_block_rl ;
	7'h0b :
		TR_17 = RG_quantized_block_rl ;
	7'h0c :
		TR_17 = RG_quantized_block_rl ;
	7'h0d :
		TR_17 = RG_quantized_block_rl ;
	7'h0e :
		TR_17 = RG_quantized_block_rl ;
	7'h0f :
		TR_17 = RG_quantized_block_rl ;
	7'h10 :
		TR_17 = RG_quantized_block_rl ;
	7'h11 :
		TR_17 = RG_quantized_block_rl ;
	7'h12 :
		TR_17 = RG_quantized_block_rl ;
	7'h13 :
		TR_17 = RG_quantized_block_rl ;
	7'h14 :
		TR_17 = RG_quantized_block_rl ;
	7'h15 :
		TR_17 = RG_quantized_block_rl ;
	7'h16 :
		TR_17 = RG_quantized_block_rl ;
	7'h17 :
		TR_17 = RG_quantized_block_rl ;
	7'h18 :
		TR_17 = RG_quantized_block_rl ;
	7'h19 :
		TR_17 = RG_quantized_block_rl ;
	7'h1a :
		TR_17 = RG_quantized_block_rl ;
	7'h1b :
		TR_17 = RG_quantized_block_rl ;
	7'h1c :
		TR_17 = RG_quantized_block_rl ;
	7'h1d :
		TR_17 = RG_quantized_block_rl ;
	7'h1e :
		TR_17 = RG_quantized_block_rl ;
	7'h1f :
		TR_17 = RG_quantized_block_rl ;
	7'h20 :
		TR_17 = RG_quantized_block_rl ;
	7'h21 :
		TR_17 = RG_quantized_block_rl ;
	7'h22 :
		TR_17 = RG_quantized_block_rl ;
	7'h23 :
		TR_17 = RG_quantized_block_rl ;
	7'h24 :
		TR_17 = RG_quantized_block_rl ;
	7'h25 :
		TR_17 = RG_quantized_block_rl ;
	7'h26 :
		TR_17 = RG_quantized_block_rl ;
	7'h27 :
		TR_17 = RG_quantized_block_rl ;
	7'h28 :
		TR_17 = RG_quantized_block_rl ;
	7'h29 :
		TR_17 = RG_quantized_block_rl ;
	7'h2a :
		TR_17 = RG_quantized_block_rl ;
	7'h2b :
		TR_17 = RG_quantized_block_rl ;
	7'h2c :
		TR_17 = RG_quantized_block_rl ;
	7'h2d :
		TR_17 = RG_quantized_block_rl ;
	7'h2e :
		TR_17 = RG_quantized_block_rl ;
	7'h2f :
		TR_17 = RG_quantized_block_rl ;
	7'h30 :
		TR_17 = RG_quantized_block_rl ;
	7'h31 :
		TR_17 = RG_quantized_block_rl ;
	7'h32 :
		TR_17 = RG_quantized_block_rl ;
	7'h33 :
		TR_17 = RG_quantized_block_rl ;
	7'h34 :
		TR_17 = RG_quantized_block_rl ;
	7'h35 :
		TR_17 = RG_quantized_block_rl ;
	7'h36 :
		TR_17 = RG_quantized_block_rl ;
	7'h37 :
		TR_17 = RG_quantized_block_rl ;
	7'h38 :
		TR_17 = RG_quantized_block_rl ;
	7'h39 :
		TR_17 = RG_quantized_block_rl ;
	7'h3a :
		TR_17 = RG_quantized_block_rl ;
	7'h3b :
		TR_17 = RG_quantized_block_rl ;
	7'h3c :
		TR_17 = RG_quantized_block_rl ;
	7'h3d :
		TR_17 = RG_quantized_block_rl ;
	7'h3e :
		TR_17 = RG_quantized_block_rl ;
	7'h3f :
		TR_17 = RG_quantized_block_rl ;
	7'h40 :
		TR_17 = RG_quantized_block_rl ;
	7'h41 :
		TR_17 = RG_quantized_block_rl ;
	7'h42 :
		TR_17 = RG_quantized_block_rl ;
	7'h43 :
		TR_17 = RG_quantized_block_rl ;
	7'h44 :
		TR_17 = RG_quantized_block_rl ;
	7'h45 :
		TR_17 = RG_quantized_block_rl ;
	7'h46 :
		TR_17 = RG_quantized_block_rl ;
	7'h47 :
		TR_17 = RG_quantized_block_rl ;
	7'h48 :
		TR_17 = RG_quantized_block_rl ;
	7'h49 :
		TR_17 = RG_quantized_block_rl ;
	7'h4a :
		TR_17 = RG_quantized_block_rl ;
	7'h4b :
		TR_17 = RG_quantized_block_rl ;
	7'h4c :
		TR_17 = RG_quantized_block_rl ;
	7'h4d :
		TR_17 = RG_quantized_block_rl ;
	7'h4e :
		TR_17 = RG_quantized_block_rl ;
	7'h4f :
		TR_17 = RG_quantized_block_rl ;
	7'h50 :
		TR_17 = RG_quantized_block_rl ;
	7'h51 :
		TR_17 = RG_quantized_block_rl ;
	7'h52 :
		TR_17 = RG_quantized_block_rl ;
	7'h53 :
		TR_17 = RG_quantized_block_rl ;
	7'h54 :
		TR_17 = RG_quantized_block_rl ;
	7'h55 :
		TR_17 = RG_quantized_block_rl ;
	7'h56 :
		TR_17 = RG_quantized_block_rl ;
	7'h57 :
		TR_17 = RG_quantized_block_rl ;
	7'h58 :
		TR_17 = RG_quantized_block_rl ;
	7'h59 :
		TR_17 = RG_quantized_block_rl ;
	7'h5a :
		TR_17 = RG_quantized_block_rl ;
	7'h5b :
		TR_17 = RG_quantized_block_rl ;
	7'h5c :
		TR_17 = RG_quantized_block_rl ;
	7'h5d :
		TR_17 = RG_quantized_block_rl ;
	7'h5e :
		TR_17 = RG_quantized_block_rl ;
	7'h5f :
		TR_17 = RG_quantized_block_rl ;
	7'h60 :
		TR_17 = RG_quantized_block_rl ;
	7'h61 :
		TR_17 = RG_quantized_block_rl ;
	7'h62 :
		TR_17 = RG_quantized_block_rl ;
	7'h63 :
		TR_17 = RG_quantized_block_rl ;
	7'h64 :
		TR_17 = RG_quantized_block_rl ;
	7'h65 :
		TR_17 = RG_quantized_block_rl ;
	7'h66 :
		TR_17 = RG_quantized_block_rl ;
	7'h67 :
		TR_17 = RG_quantized_block_rl ;
	7'h68 :
		TR_17 = RG_quantized_block_rl ;
	7'h69 :
		TR_17 = RG_quantized_block_rl ;
	7'h6a :
		TR_17 = RG_quantized_block_rl ;
	7'h6b :
		TR_17 = RG_quantized_block_rl ;
	7'h6c :
		TR_17 = RG_quantized_block_rl ;
	7'h6d :
		TR_17 = RG_quantized_block_rl ;
	7'h6e :
		TR_17 = RG_quantized_block_rl ;
	7'h6f :
		TR_17 = RG_quantized_block_rl ;
	7'h70 :
		TR_17 = RG_quantized_block_rl ;
	7'h71 :
		TR_17 = RG_quantized_block_rl ;
	7'h72 :
		TR_17 = RG_quantized_block_rl ;
	7'h73 :
		TR_17 = RG_quantized_block_rl ;
	7'h74 :
		TR_17 = RG_quantized_block_rl ;
	7'h75 :
		TR_17 = RG_quantized_block_rl ;
	7'h76 :
		TR_17 = RG_quantized_block_rl ;
	7'h77 :
		TR_17 = RG_quantized_block_rl ;
	7'h78 :
		TR_17 = RG_quantized_block_rl ;
	7'h79 :
		TR_17 = RG_quantized_block_rl ;
	7'h7a :
		TR_17 = RG_quantized_block_rl ;
	7'h7b :
		TR_17 = RG_quantized_block_rl ;
	7'h7c :
		TR_17 = RG_quantized_block_rl ;
	7'h7d :
		TR_17 = RG_quantized_block_rl ;
	7'h7e :
		TR_17 = RG_quantized_block_rl ;
	7'h7f :
		TR_17 = RG_quantized_block_rl ;
	default :
		TR_17 = 9'hx ;
	endcase
always @ ( RG_rl_132 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_18 = RG_rl_132 ;
	7'h01 :
		TR_18 = RG_rl_132 ;
	7'h02 :
		TR_18 = RG_rl_132 ;
	7'h03 :
		TR_18 = RG_rl_132 ;
	7'h04 :
		TR_18 = RG_rl_132 ;
	7'h05 :
		TR_18 = RG_rl_132 ;
	7'h06 :
		TR_18 = 9'h000 ;	// line#=../rle.cpp:79
	7'h07 :
		TR_18 = RG_rl_132 ;
	7'h08 :
		TR_18 = RG_rl_132 ;
	7'h09 :
		TR_18 = RG_rl_132 ;
	7'h0a :
		TR_18 = RG_rl_132 ;
	7'h0b :
		TR_18 = RG_rl_132 ;
	7'h0c :
		TR_18 = RG_rl_132 ;
	7'h0d :
		TR_18 = RG_rl_132 ;
	7'h0e :
		TR_18 = RG_rl_132 ;
	7'h0f :
		TR_18 = RG_rl_132 ;
	7'h10 :
		TR_18 = RG_rl_132 ;
	7'h11 :
		TR_18 = RG_rl_132 ;
	7'h12 :
		TR_18 = RG_rl_132 ;
	7'h13 :
		TR_18 = RG_rl_132 ;
	7'h14 :
		TR_18 = RG_rl_132 ;
	7'h15 :
		TR_18 = RG_rl_132 ;
	7'h16 :
		TR_18 = RG_rl_132 ;
	7'h17 :
		TR_18 = RG_rl_132 ;
	7'h18 :
		TR_18 = RG_rl_132 ;
	7'h19 :
		TR_18 = RG_rl_132 ;
	7'h1a :
		TR_18 = RG_rl_132 ;
	7'h1b :
		TR_18 = RG_rl_132 ;
	7'h1c :
		TR_18 = RG_rl_132 ;
	7'h1d :
		TR_18 = RG_rl_132 ;
	7'h1e :
		TR_18 = RG_rl_132 ;
	7'h1f :
		TR_18 = RG_rl_132 ;
	7'h20 :
		TR_18 = RG_rl_132 ;
	7'h21 :
		TR_18 = RG_rl_132 ;
	7'h22 :
		TR_18 = RG_rl_132 ;
	7'h23 :
		TR_18 = RG_rl_132 ;
	7'h24 :
		TR_18 = RG_rl_132 ;
	7'h25 :
		TR_18 = RG_rl_132 ;
	7'h26 :
		TR_18 = RG_rl_132 ;
	7'h27 :
		TR_18 = RG_rl_132 ;
	7'h28 :
		TR_18 = RG_rl_132 ;
	7'h29 :
		TR_18 = RG_rl_132 ;
	7'h2a :
		TR_18 = RG_rl_132 ;
	7'h2b :
		TR_18 = RG_rl_132 ;
	7'h2c :
		TR_18 = RG_rl_132 ;
	7'h2d :
		TR_18 = RG_rl_132 ;
	7'h2e :
		TR_18 = RG_rl_132 ;
	7'h2f :
		TR_18 = RG_rl_132 ;
	7'h30 :
		TR_18 = RG_rl_132 ;
	7'h31 :
		TR_18 = RG_rl_132 ;
	7'h32 :
		TR_18 = RG_rl_132 ;
	7'h33 :
		TR_18 = RG_rl_132 ;
	7'h34 :
		TR_18 = RG_rl_132 ;
	7'h35 :
		TR_18 = RG_rl_132 ;
	7'h36 :
		TR_18 = RG_rl_132 ;
	7'h37 :
		TR_18 = RG_rl_132 ;
	7'h38 :
		TR_18 = RG_rl_132 ;
	7'h39 :
		TR_18 = RG_rl_132 ;
	7'h3a :
		TR_18 = RG_rl_132 ;
	7'h3b :
		TR_18 = RG_rl_132 ;
	7'h3c :
		TR_18 = RG_rl_132 ;
	7'h3d :
		TR_18 = RG_rl_132 ;
	7'h3e :
		TR_18 = RG_rl_132 ;
	7'h3f :
		TR_18 = RG_rl_132 ;
	7'h40 :
		TR_18 = RG_rl_132 ;
	7'h41 :
		TR_18 = RG_rl_132 ;
	7'h42 :
		TR_18 = RG_rl_132 ;
	7'h43 :
		TR_18 = RG_rl_132 ;
	7'h44 :
		TR_18 = RG_rl_132 ;
	7'h45 :
		TR_18 = RG_rl_132 ;
	7'h46 :
		TR_18 = RG_rl_132 ;
	7'h47 :
		TR_18 = RG_rl_132 ;
	7'h48 :
		TR_18 = RG_rl_132 ;
	7'h49 :
		TR_18 = RG_rl_132 ;
	7'h4a :
		TR_18 = RG_rl_132 ;
	7'h4b :
		TR_18 = RG_rl_132 ;
	7'h4c :
		TR_18 = RG_rl_132 ;
	7'h4d :
		TR_18 = RG_rl_132 ;
	7'h4e :
		TR_18 = RG_rl_132 ;
	7'h4f :
		TR_18 = RG_rl_132 ;
	7'h50 :
		TR_18 = RG_rl_132 ;
	7'h51 :
		TR_18 = RG_rl_132 ;
	7'h52 :
		TR_18 = RG_rl_132 ;
	7'h53 :
		TR_18 = RG_rl_132 ;
	7'h54 :
		TR_18 = RG_rl_132 ;
	7'h55 :
		TR_18 = RG_rl_132 ;
	7'h56 :
		TR_18 = RG_rl_132 ;
	7'h57 :
		TR_18 = RG_rl_132 ;
	7'h58 :
		TR_18 = RG_rl_132 ;
	7'h59 :
		TR_18 = RG_rl_132 ;
	7'h5a :
		TR_18 = RG_rl_132 ;
	7'h5b :
		TR_18 = RG_rl_132 ;
	7'h5c :
		TR_18 = RG_rl_132 ;
	7'h5d :
		TR_18 = RG_rl_132 ;
	7'h5e :
		TR_18 = RG_rl_132 ;
	7'h5f :
		TR_18 = RG_rl_132 ;
	7'h60 :
		TR_18 = RG_rl_132 ;
	7'h61 :
		TR_18 = RG_rl_132 ;
	7'h62 :
		TR_18 = RG_rl_132 ;
	7'h63 :
		TR_18 = RG_rl_132 ;
	7'h64 :
		TR_18 = RG_rl_132 ;
	7'h65 :
		TR_18 = RG_rl_132 ;
	7'h66 :
		TR_18 = RG_rl_132 ;
	7'h67 :
		TR_18 = RG_rl_132 ;
	7'h68 :
		TR_18 = RG_rl_132 ;
	7'h69 :
		TR_18 = RG_rl_132 ;
	7'h6a :
		TR_18 = RG_rl_132 ;
	7'h6b :
		TR_18 = RG_rl_132 ;
	7'h6c :
		TR_18 = RG_rl_132 ;
	7'h6d :
		TR_18 = RG_rl_132 ;
	7'h6e :
		TR_18 = RG_rl_132 ;
	7'h6f :
		TR_18 = RG_rl_132 ;
	7'h70 :
		TR_18 = RG_rl_132 ;
	7'h71 :
		TR_18 = RG_rl_132 ;
	7'h72 :
		TR_18 = RG_rl_132 ;
	7'h73 :
		TR_18 = RG_rl_132 ;
	7'h74 :
		TR_18 = RG_rl_132 ;
	7'h75 :
		TR_18 = RG_rl_132 ;
	7'h76 :
		TR_18 = RG_rl_132 ;
	7'h77 :
		TR_18 = RG_rl_132 ;
	7'h78 :
		TR_18 = RG_rl_132 ;
	7'h79 :
		TR_18 = RG_rl_132 ;
	7'h7a :
		TR_18 = RG_rl_132 ;
	7'h7b :
		TR_18 = RG_rl_132 ;
	7'h7c :
		TR_18 = RG_rl_132 ;
	7'h7d :
		TR_18 = RG_rl_132 ;
	7'h7e :
		TR_18 = RG_rl_132 ;
	7'h7f :
		TR_18 = RG_rl_132 ;
	default :
		TR_18 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_1 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h01 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h02 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h03 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h04 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h05 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h06 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h07 :
		TR_19 = 9'h000 ;	// line#=../rle.cpp:79
	7'h08 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h09 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h0a :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h0b :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h0c :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h0d :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h0e :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h0f :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h10 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h11 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h12 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h13 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h14 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h15 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h16 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h17 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h18 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h19 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h1a :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h1b :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h1c :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h1d :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h1e :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h1f :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h20 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h21 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h22 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h23 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h24 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h25 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h26 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h27 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h28 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h29 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h2a :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h2b :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h2c :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h2d :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h2e :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h2f :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h30 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h31 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h32 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h33 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h34 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h35 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h36 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h37 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h38 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h39 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h3a :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h3b :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h3c :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h3d :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h3e :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h3f :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h40 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h41 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h42 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h43 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h44 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h45 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h46 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h47 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h48 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h49 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h4a :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h4b :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h4c :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h4d :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h4e :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h4f :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h50 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h51 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h52 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h53 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h54 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h55 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h56 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h57 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h58 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h59 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h5a :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h5b :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h5c :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h5d :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h5e :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h5f :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h60 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h61 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h62 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h63 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h64 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h65 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h66 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h67 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h68 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h69 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h6a :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h6b :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h6c :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h6d :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h6e :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h6f :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h70 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h71 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h72 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h73 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h74 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h75 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h76 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h77 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h78 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h79 :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h7a :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h7b :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h7c :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h7d :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h7e :
		TR_19 = RG_quantized_block_rl_1 ;
	7'h7f :
		TR_19 = RG_quantized_block_rl_1 ;
	default :
		TR_19 = 9'hx ;
	endcase
always @ ( RG_rl_133 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_20 = RG_rl_133 ;
	7'h01 :
		TR_20 = RG_rl_133 ;
	7'h02 :
		TR_20 = RG_rl_133 ;
	7'h03 :
		TR_20 = RG_rl_133 ;
	7'h04 :
		TR_20 = RG_rl_133 ;
	7'h05 :
		TR_20 = RG_rl_133 ;
	7'h06 :
		TR_20 = RG_rl_133 ;
	7'h07 :
		TR_20 = RG_rl_133 ;
	7'h08 :
		TR_20 = 9'h000 ;	// line#=../rle.cpp:79
	7'h09 :
		TR_20 = RG_rl_133 ;
	7'h0a :
		TR_20 = RG_rl_133 ;
	7'h0b :
		TR_20 = RG_rl_133 ;
	7'h0c :
		TR_20 = RG_rl_133 ;
	7'h0d :
		TR_20 = RG_rl_133 ;
	7'h0e :
		TR_20 = RG_rl_133 ;
	7'h0f :
		TR_20 = RG_rl_133 ;
	7'h10 :
		TR_20 = RG_rl_133 ;
	7'h11 :
		TR_20 = RG_rl_133 ;
	7'h12 :
		TR_20 = RG_rl_133 ;
	7'h13 :
		TR_20 = RG_rl_133 ;
	7'h14 :
		TR_20 = RG_rl_133 ;
	7'h15 :
		TR_20 = RG_rl_133 ;
	7'h16 :
		TR_20 = RG_rl_133 ;
	7'h17 :
		TR_20 = RG_rl_133 ;
	7'h18 :
		TR_20 = RG_rl_133 ;
	7'h19 :
		TR_20 = RG_rl_133 ;
	7'h1a :
		TR_20 = RG_rl_133 ;
	7'h1b :
		TR_20 = RG_rl_133 ;
	7'h1c :
		TR_20 = RG_rl_133 ;
	7'h1d :
		TR_20 = RG_rl_133 ;
	7'h1e :
		TR_20 = RG_rl_133 ;
	7'h1f :
		TR_20 = RG_rl_133 ;
	7'h20 :
		TR_20 = RG_rl_133 ;
	7'h21 :
		TR_20 = RG_rl_133 ;
	7'h22 :
		TR_20 = RG_rl_133 ;
	7'h23 :
		TR_20 = RG_rl_133 ;
	7'h24 :
		TR_20 = RG_rl_133 ;
	7'h25 :
		TR_20 = RG_rl_133 ;
	7'h26 :
		TR_20 = RG_rl_133 ;
	7'h27 :
		TR_20 = RG_rl_133 ;
	7'h28 :
		TR_20 = RG_rl_133 ;
	7'h29 :
		TR_20 = RG_rl_133 ;
	7'h2a :
		TR_20 = RG_rl_133 ;
	7'h2b :
		TR_20 = RG_rl_133 ;
	7'h2c :
		TR_20 = RG_rl_133 ;
	7'h2d :
		TR_20 = RG_rl_133 ;
	7'h2e :
		TR_20 = RG_rl_133 ;
	7'h2f :
		TR_20 = RG_rl_133 ;
	7'h30 :
		TR_20 = RG_rl_133 ;
	7'h31 :
		TR_20 = RG_rl_133 ;
	7'h32 :
		TR_20 = RG_rl_133 ;
	7'h33 :
		TR_20 = RG_rl_133 ;
	7'h34 :
		TR_20 = RG_rl_133 ;
	7'h35 :
		TR_20 = RG_rl_133 ;
	7'h36 :
		TR_20 = RG_rl_133 ;
	7'h37 :
		TR_20 = RG_rl_133 ;
	7'h38 :
		TR_20 = RG_rl_133 ;
	7'h39 :
		TR_20 = RG_rl_133 ;
	7'h3a :
		TR_20 = RG_rl_133 ;
	7'h3b :
		TR_20 = RG_rl_133 ;
	7'h3c :
		TR_20 = RG_rl_133 ;
	7'h3d :
		TR_20 = RG_rl_133 ;
	7'h3e :
		TR_20 = RG_rl_133 ;
	7'h3f :
		TR_20 = RG_rl_133 ;
	7'h40 :
		TR_20 = RG_rl_133 ;
	7'h41 :
		TR_20 = RG_rl_133 ;
	7'h42 :
		TR_20 = RG_rl_133 ;
	7'h43 :
		TR_20 = RG_rl_133 ;
	7'h44 :
		TR_20 = RG_rl_133 ;
	7'h45 :
		TR_20 = RG_rl_133 ;
	7'h46 :
		TR_20 = RG_rl_133 ;
	7'h47 :
		TR_20 = RG_rl_133 ;
	7'h48 :
		TR_20 = RG_rl_133 ;
	7'h49 :
		TR_20 = RG_rl_133 ;
	7'h4a :
		TR_20 = RG_rl_133 ;
	7'h4b :
		TR_20 = RG_rl_133 ;
	7'h4c :
		TR_20 = RG_rl_133 ;
	7'h4d :
		TR_20 = RG_rl_133 ;
	7'h4e :
		TR_20 = RG_rl_133 ;
	7'h4f :
		TR_20 = RG_rl_133 ;
	7'h50 :
		TR_20 = RG_rl_133 ;
	7'h51 :
		TR_20 = RG_rl_133 ;
	7'h52 :
		TR_20 = RG_rl_133 ;
	7'h53 :
		TR_20 = RG_rl_133 ;
	7'h54 :
		TR_20 = RG_rl_133 ;
	7'h55 :
		TR_20 = RG_rl_133 ;
	7'h56 :
		TR_20 = RG_rl_133 ;
	7'h57 :
		TR_20 = RG_rl_133 ;
	7'h58 :
		TR_20 = RG_rl_133 ;
	7'h59 :
		TR_20 = RG_rl_133 ;
	7'h5a :
		TR_20 = RG_rl_133 ;
	7'h5b :
		TR_20 = RG_rl_133 ;
	7'h5c :
		TR_20 = RG_rl_133 ;
	7'h5d :
		TR_20 = RG_rl_133 ;
	7'h5e :
		TR_20 = RG_rl_133 ;
	7'h5f :
		TR_20 = RG_rl_133 ;
	7'h60 :
		TR_20 = RG_rl_133 ;
	7'h61 :
		TR_20 = RG_rl_133 ;
	7'h62 :
		TR_20 = RG_rl_133 ;
	7'h63 :
		TR_20 = RG_rl_133 ;
	7'h64 :
		TR_20 = RG_rl_133 ;
	7'h65 :
		TR_20 = RG_rl_133 ;
	7'h66 :
		TR_20 = RG_rl_133 ;
	7'h67 :
		TR_20 = RG_rl_133 ;
	7'h68 :
		TR_20 = RG_rl_133 ;
	7'h69 :
		TR_20 = RG_rl_133 ;
	7'h6a :
		TR_20 = RG_rl_133 ;
	7'h6b :
		TR_20 = RG_rl_133 ;
	7'h6c :
		TR_20 = RG_rl_133 ;
	7'h6d :
		TR_20 = RG_rl_133 ;
	7'h6e :
		TR_20 = RG_rl_133 ;
	7'h6f :
		TR_20 = RG_rl_133 ;
	7'h70 :
		TR_20 = RG_rl_133 ;
	7'h71 :
		TR_20 = RG_rl_133 ;
	7'h72 :
		TR_20 = RG_rl_133 ;
	7'h73 :
		TR_20 = RG_rl_133 ;
	7'h74 :
		TR_20 = RG_rl_133 ;
	7'h75 :
		TR_20 = RG_rl_133 ;
	7'h76 :
		TR_20 = RG_rl_133 ;
	7'h77 :
		TR_20 = RG_rl_133 ;
	7'h78 :
		TR_20 = RG_rl_133 ;
	7'h79 :
		TR_20 = RG_rl_133 ;
	7'h7a :
		TR_20 = RG_rl_133 ;
	7'h7b :
		TR_20 = RG_rl_133 ;
	7'h7c :
		TR_20 = RG_rl_133 ;
	7'h7d :
		TR_20 = RG_rl_133 ;
	7'h7e :
		TR_20 = RG_rl_133 ;
	7'h7f :
		TR_20 = RG_rl_133 ;
	default :
		TR_20 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_2 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h01 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h02 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h03 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h04 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h05 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h06 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h07 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h08 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h09 :
		TR_21 = 9'h000 ;	// line#=../rle.cpp:79
	7'h0a :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h0b :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h0c :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h0d :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h0e :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h0f :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h10 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h11 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h12 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h13 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h14 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h15 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h16 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h17 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h18 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h19 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h1a :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h1b :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h1c :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h1d :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h1e :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h1f :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h20 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h21 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h22 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h23 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h24 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h25 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h26 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h27 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h28 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h29 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h2a :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h2b :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h2c :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h2d :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h2e :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h2f :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h30 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h31 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h32 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h33 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h34 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h35 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h36 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h37 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h38 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h39 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h3a :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h3b :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h3c :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h3d :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h3e :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h3f :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h40 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h41 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h42 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h43 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h44 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h45 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h46 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h47 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h48 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h49 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h4a :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h4b :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h4c :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h4d :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h4e :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h4f :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h50 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h51 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h52 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h53 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h54 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h55 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h56 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h57 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h58 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h59 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h5a :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h5b :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h5c :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h5d :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h5e :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h5f :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h60 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h61 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h62 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h63 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h64 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h65 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h66 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h67 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h68 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h69 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h6a :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h6b :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h6c :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h6d :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h6e :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h6f :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h70 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h71 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h72 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h73 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h74 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h75 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h76 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h77 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h78 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h79 :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h7a :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h7b :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h7c :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h7d :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h7e :
		TR_21 = RG_quantized_block_rl_2 ;
	7'h7f :
		TR_21 = RG_quantized_block_rl_2 ;
	default :
		TR_21 = 9'hx ;
	endcase
always @ ( RG_rl_134 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_22 = RG_rl_134 ;
	7'h01 :
		TR_22 = RG_rl_134 ;
	7'h02 :
		TR_22 = RG_rl_134 ;
	7'h03 :
		TR_22 = RG_rl_134 ;
	7'h04 :
		TR_22 = RG_rl_134 ;
	7'h05 :
		TR_22 = RG_rl_134 ;
	7'h06 :
		TR_22 = RG_rl_134 ;
	7'h07 :
		TR_22 = RG_rl_134 ;
	7'h08 :
		TR_22 = RG_rl_134 ;
	7'h09 :
		TR_22 = RG_rl_134 ;
	7'h0a :
		TR_22 = 9'h000 ;	// line#=../rle.cpp:79
	7'h0b :
		TR_22 = RG_rl_134 ;
	7'h0c :
		TR_22 = RG_rl_134 ;
	7'h0d :
		TR_22 = RG_rl_134 ;
	7'h0e :
		TR_22 = RG_rl_134 ;
	7'h0f :
		TR_22 = RG_rl_134 ;
	7'h10 :
		TR_22 = RG_rl_134 ;
	7'h11 :
		TR_22 = RG_rl_134 ;
	7'h12 :
		TR_22 = RG_rl_134 ;
	7'h13 :
		TR_22 = RG_rl_134 ;
	7'h14 :
		TR_22 = RG_rl_134 ;
	7'h15 :
		TR_22 = RG_rl_134 ;
	7'h16 :
		TR_22 = RG_rl_134 ;
	7'h17 :
		TR_22 = RG_rl_134 ;
	7'h18 :
		TR_22 = RG_rl_134 ;
	7'h19 :
		TR_22 = RG_rl_134 ;
	7'h1a :
		TR_22 = RG_rl_134 ;
	7'h1b :
		TR_22 = RG_rl_134 ;
	7'h1c :
		TR_22 = RG_rl_134 ;
	7'h1d :
		TR_22 = RG_rl_134 ;
	7'h1e :
		TR_22 = RG_rl_134 ;
	7'h1f :
		TR_22 = RG_rl_134 ;
	7'h20 :
		TR_22 = RG_rl_134 ;
	7'h21 :
		TR_22 = RG_rl_134 ;
	7'h22 :
		TR_22 = RG_rl_134 ;
	7'h23 :
		TR_22 = RG_rl_134 ;
	7'h24 :
		TR_22 = RG_rl_134 ;
	7'h25 :
		TR_22 = RG_rl_134 ;
	7'h26 :
		TR_22 = RG_rl_134 ;
	7'h27 :
		TR_22 = RG_rl_134 ;
	7'h28 :
		TR_22 = RG_rl_134 ;
	7'h29 :
		TR_22 = RG_rl_134 ;
	7'h2a :
		TR_22 = RG_rl_134 ;
	7'h2b :
		TR_22 = RG_rl_134 ;
	7'h2c :
		TR_22 = RG_rl_134 ;
	7'h2d :
		TR_22 = RG_rl_134 ;
	7'h2e :
		TR_22 = RG_rl_134 ;
	7'h2f :
		TR_22 = RG_rl_134 ;
	7'h30 :
		TR_22 = RG_rl_134 ;
	7'h31 :
		TR_22 = RG_rl_134 ;
	7'h32 :
		TR_22 = RG_rl_134 ;
	7'h33 :
		TR_22 = RG_rl_134 ;
	7'h34 :
		TR_22 = RG_rl_134 ;
	7'h35 :
		TR_22 = RG_rl_134 ;
	7'h36 :
		TR_22 = RG_rl_134 ;
	7'h37 :
		TR_22 = RG_rl_134 ;
	7'h38 :
		TR_22 = RG_rl_134 ;
	7'h39 :
		TR_22 = RG_rl_134 ;
	7'h3a :
		TR_22 = RG_rl_134 ;
	7'h3b :
		TR_22 = RG_rl_134 ;
	7'h3c :
		TR_22 = RG_rl_134 ;
	7'h3d :
		TR_22 = RG_rl_134 ;
	7'h3e :
		TR_22 = RG_rl_134 ;
	7'h3f :
		TR_22 = RG_rl_134 ;
	7'h40 :
		TR_22 = RG_rl_134 ;
	7'h41 :
		TR_22 = RG_rl_134 ;
	7'h42 :
		TR_22 = RG_rl_134 ;
	7'h43 :
		TR_22 = RG_rl_134 ;
	7'h44 :
		TR_22 = RG_rl_134 ;
	7'h45 :
		TR_22 = RG_rl_134 ;
	7'h46 :
		TR_22 = RG_rl_134 ;
	7'h47 :
		TR_22 = RG_rl_134 ;
	7'h48 :
		TR_22 = RG_rl_134 ;
	7'h49 :
		TR_22 = RG_rl_134 ;
	7'h4a :
		TR_22 = RG_rl_134 ;
	7'h4b :
		TR_22 = RG_rl_134 ;
	7'h4c :
		TR_22 = RG_rl_134 ;
	7'h4d :
		TR_22 = RG_rl_134 ;
	7'h4e :
		TR_22 = RG_rl_134 ;
	7'h4f :
		TR_22 = RG_rl_134 ;
	7'h50 :
		TR_22 = RG_rl_134 ;
	7'h51 :
		TR_22 = RG_rl_134 ;
	7'h52 :
		TR_22 = RG_rl_134 ;
	7'h53 :
		TR_22 = RG_rl_134 ;
	7'h54 :
		TR_22 = RG_rl_134 ;
	7'h55 :
		TR_22 = RG_rl_134 ;
	7'h56 :
		TR_22 = RG_rl_134 ;
	7'h57 :
		TR_22 = RG_rl_134 ;
	7'h58 :
		TR_22 = RG_rl_134 ;
	7'h59 :
		TR_22 = RG_rl_134 ;
	7'h5a :
		TR_22 = RG_rl_134 ;
	7'h5b :
		TR_22 = RG_rl_134 ;
	7'h5c :
		TR_22 = RG_rl_134 ;
	7'h5d :
		TR_22 = RG_rl_134 ;
	7'h5e :
		TR_22 = RG_rl_134 ;
	7'h5f :
		TR_22 = RG_rl_134 ;
	7'h60 :
		TR_22 = RG_rl_134 ;
	7'h61 :
		TR_22 = RG_rl_134 ;
	7'h62 :
		TR_22 = RG_rl_134 ;
	7'h63 :
		TR_22 = RG_rl_134 ;
	7'h64 :
		TR_22 = RG_rl_134 ;
	7'h65 :
		TR_22 = RG_rl_134 ;
	7'h66 :
		TR_22 = RG_rl_134 ;
	7'h67 :
		TR_22 = RG_rl_134 ;
	7'h68 :
		TR_22 = RG_rl_134 ;
	7'h69 :
		TR_22 = RG_rl_134 ;
	7'h6a :
		TR_22 = RG_rl_134 ;
	7'h6b :
		TR_22 = RG_rl_134 ;
	7'h6c :
		TR_22 = RG_rl_134 ;
	7'h6d :
		TR_22 = RG_rl_134 ;
	7'h6e :
		TR_22 = RG_rl_134 ;
	7'h6f :
		TR_22 = RG_rl_134 ;
	7'h70 :
		TR_22 = RG_rl_134 ;
	7'h71 :
		TR_22 = RG_rl_134 ;
	7'h72 :
		TR_22 = RG_rl_134 ;
	7'h73 :
		TR_22 = RG_rl_134 ;
	7'h74 :
		TR_22 = RG_rl_134 ;
	7'h75 :
		TR_22 = RG_rl_134 ;
	7'h76 :
		TR_22 = RG_rl_134 ;
	7'h77 :
		TR_22 = RG_rl_134 ;
	7'h78 :
		TR_22 = RG_rl_134 ;
	7'h79 :
		TR_22 = RG_rl_134 ;
	7'h7a :
		TR_22 = RG_rl_134 ;
	7'h7b :
		TR_22 = RG_rl_134 ;
	7'h7c :
		TR_22 = RG_rl_134 ;
	7'h7d :
		TR_22 = RG_rl_134 ;
	7'h7e :
		TR_22 = RG_rl_134 ;
	7'h7f :
		TR_22 = RG_rl_134 ;
	default :
		TR_22 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_3 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h01 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h02 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h03 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h04 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h05 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h06 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h07 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h08 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h09 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h0a :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h0b :
		TR_23 = 9'h000 ;	// line#=../rle.cpp:79
	7'h0c :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h0d :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h0e :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h0f :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h10 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h11 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h12 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h13 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h14 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h15 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h16 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h17 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h18 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h19 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h1a :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h1b :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h1c :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h1d :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h1e :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h1f :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h20 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h21 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h22 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h23 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h24 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h25 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h26 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h27 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h28 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h29 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h2a :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h2b :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h2c :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h2d :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h2e :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h2f :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h30 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h31 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h32 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h33 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h34 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h35 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h36 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h37 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h38 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h39 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h3a :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h3b :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h3c :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h3d :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h3e :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h3f :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h40 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h41 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h42 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h43 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h44 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h45 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h46 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h47 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h48 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h49 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h4a :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h4b :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h4c :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h4d :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h4e :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h4f :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h50 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h51 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h52 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h53 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h54 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h55 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h56 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h57 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h58 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h59 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h5a :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h5b :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h5c :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h5d :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h5e :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h5f :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h60 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h61 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h62 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h63 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h64 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h65 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h66 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h67 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h68 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h69 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h6a :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h6b :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h6c :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h6d :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h6e :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h6f :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h70 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h71 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h72 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h73 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h74 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h75 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h76 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h77 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h78 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h79 :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h7a :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h7b :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h7c :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h7d :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h7e :
		TR_23 = RG_quantized_block_rl_3 ;
	7'h7f :
		TR_23 = RG_quantized_block_rl_3 ;
	default :
		TR_23 = 9'hx ;
	endcase
always @ ( RG_rl_135 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_24 = RG_rl_135 ;
	7'h01 :
		TR_24 = RG_rl_135 ;
	7'h02 :
		TR_24 = RG_rl_135 ;
	7'h03 :
		TR_24 = RG_rl_135 ;
	7'h04 :
		TR_24 = RG_rl_135 ;
	7'h05 :
		TR_24 = RG_rl_135 ;
	7'h06 :
		TR_24 = RG_rl_135 ;
	7'h07 :
		TR_24 = RG_rl_135 ;
	7'h08 :
		TR_24 = RG_rl_135 ;
	7'h09 :
		TR_24 = RG_rl_135 ;
	7'h0a :
		TR_24 = RG_rl_135 ;
	7'h0b :
		TR_24 = RG_rl_135 ;
	7'h0c :
		TR_24 = 9'h000 ;	// line#=../rle.cpp:79
	7'h0d :
		TR_24 = RG_rl_135 ;
	7'h0e :
		TR_24 = RG_rl_135 ;
	7'h0f :
		TR_24 = RG_rl_135 ;
	7'h10 :
		TR_24 = RG_rl_135 ;
	7'h11 :
		TR_24 = RG_rl_135 ;
	7'h12 :
		TR_24 = RG_rl_135 ;
	7'h13 :
		TR_24 = RG_rl_135 ;
	7'h14 :
		TR_24 = RG_rl_135 ;
	7'h15 :
		TR_24 = RG_rl_135 ;
	7'h16 :
		TR_24 = RG_rl_135 ;
	7'h17 :
		TR_24 = RG_rl_135 ;
	7'h18 :
		TR_24 = RG_rl_135 ;
	7'h19 :
		TR_24 = RG_rl_135 ;
	7'h1a :
		TR_24 = RG_rl_135 ;
	7'h1b :
		TR_24 = RG_rl_135 ;
	7'h1c :
		TR_24 = RG_rl_135 ;
	7'h1d :
		TR_24 = RG_rl_135 ;
	7'h1e :
		TR_24 = RG_rl_135 ;
	7'h1f :
		TR_24 = RG_rl_135 ;
	7'h20 :
		TR_24 = RG_rl_135 ;
	7'h21 :
		TR_24 = RG_rl_135 ;
	7'h22 :
		TR_24 = RG_rl_135 ;
	7'h23 :
		TR_24 = RG_rl_135 ;
	7'h24 :
		TR_24 = RG_rl_135 ;
	7'h25 :
		TR_24 = RG_rl_135 ;
	7'h26 :
		TR_24 = RG_rl_135 ;
	7'h27 :
		TR_24 = RG_rl_135 ;
	7'h28 :
		TR_24 = RG_rl_135 ;
	7'h29 :
		TR_24 = RG_rl_135 ;
	7'h2a :
		TR_24 = RG_rl_135 ;
	7'h2b :
		TR_24 = RG_rl_135 ;
	7'h2c :
		TR_24 = RG_rl_135 ;
	7'h2d :
		TR_24 = RG_rl_135 ;
	7'h2e :
		TR_24 = RG_rl_135 ;
	7'h2f :
		TR_24 = RG_rl_135 ;
	7'h30 :
		TR_24 = RG_rl_135 ;
	7'h31 :
		TR_24 = RG_rl_135 ;
	7'h32 :
		TR_24 = RG_rl_135 ;
	7'h33 :
		TR_24 = RG_rl_135 ;
	7'h34 :
		TR_24 = RG_rl_135 ;
	7'h35 :
		TR_24 = RG_rl_135 ;
	7'h36 :
		TR_24 = RG_rl_135 ;
	7'h37 :
		TR_24 = RG_rl_135 ;
	7'h38 :
		TR_24 = RG_rl_135 ;
	7'h39 :
		TR_24 = RG_rl_135 ;
	7'h3a :
		TR_24 = RG_rl_135 ;
	7'h3b :
		TR_24 = RG_rl_135 ;
	7'h3c :
		TR_24 = RG_rl_135 ;
	7'h3d :
		TR_24 = RG_rl_135 ;
	7'h3e :
		TR_24 = RG_rl_135 ;
	7'h3f :
		TR_24 = RG_rl_135 ;
	7'h40 :
		TR_24 = RG_rl_135 ;
	7'h41 :
		TR_24 = RG_rl_135 ;
	7'h42 :
		TR_24 = RG_rl_135 ;
	7'h43 :
		TR_24 = RG_rl_135 ;
	7'h44 :
		TR_24 = RG_rl_135 ;
	7'h45 :
		TR_24 = RG_rl_135 ;
	7'h46 :
		TR_24 = RG_rl_135 ;
	7'h47 :
		TR_24 = RG_rl_135 ;
	7'h48 :
		TR_24 = RG_rl_135 ;
	7'h49 :
		TR_24 = RG_rl_135 ;
	7'h4a :
		TR_24 = RG_rl_135 ;
	7'h4b :
		TR_24 = RG_rl_135 ;
	7'h4c :
		TR_24 = RG_rl_135 ;
	7'h4d :
		TR_24 = RG_rl_135 ;
	7'h4e :
		TR_24 = RG_rl_135 ;
	7'h4f :
		TR_24 = RG_rl_135 ;
	7'h50 :
		TR_24 = RG_rl_135 ;
	7'h51 :
		TR_24 = RG_rl_135 ;
	7'h52 :
		TR_24 = RG_rl_135 ;
	7'h53 :
		TR_24 = RG_rl_135 ;
	7'h54 :
		TR_24 = RG_rl_135 ;
	7'h55 :
		TR_24 = RG_rl_135 ;
	7'h56 :
		TR_24 = RG_rl_135 ;
	7'h57 :
		TR_24 = RG_rl_135 ;
	7'h58 :
		TR_24 = RG_rl_135 ;
	7'h59 :
		TR_24 = RG_rl_135 ;
	7'h5a :
		TR_24 = RG_rl_135 ;
	7'h5b :
		TR_24 = RG_rl_135 ;
	7'h5c :
		TR_24 = RG_rl_135 ;
	7'h5d :
		TR_24 = RG_rl_135 ;
	7'h5e :
		TR_24 = RG_rl_135 ;
	7'h5f :
		TR_24 = RG_rl_135 ;
	7'h60 :
		TR_24 = RG_rl_135 ;
	7'h61 :
		TR_24 = RG_rl_135 ;
	7'h62 :
		TR_24 = RG_rl_135 ;
	7'h63 :
		TR_24 = RG_rl_135 ;
	7'h64 :
		TR_24 = RG_rl_135 ;
	7'h65 :
		TR_24 = RG_rl_135 ;
	7'h66 :
		TR_24 = RG_rl_135 ;
	7'h67 :
		TR_24 = RG_rl_135 ;
	7'h68 :
		TR_24 = RG_rl_135 ;
	7'h69 :
		TR_24 = RG_rl_135 ;
	7'h6a :
		TR_24 = RG_rl_135 ;
	7'h6b :
		TR_24 = RG_rl_135 ;
	7'h6c :
		TR_24 = RG_rl_135 ;
	7'h6d :
		TR_24 = RG_rl_135 ;
	7'h6e :
		TR_24 = RG_rl_135 ;
	7'h6f :
		TR_24 = RG_rl_135 ;
	7'h70 :
		TR_24 = RG_rl_135 ;
	7'h71 :
		TR_24 = RG_rl_135 ;
	7'h72 :
		TR_24 = RG_rl_135 ;
	7'h73 :
		TR_24 = RG_rl_135 ;
	7'h74 :
		TR_24 = RG_rl_135 ;
	7'h75 :
		TR_24 = RG_rl_135 ;
	7'h76 :
		TR_24 = RG_rl_135 ;
	7'h77 :
		TR_24 = RG_rl_135 ;
	7'h78 :
		TR_24 = RG_rl_135 ;
	7'h79 :
		TR_24 = RG_rl_135 ;
	7'h7a :
		TR_24 = RG_rl_135 ;
	7'h7b :
		TR_24 = RG_rl_135 ;
	7'h7c :
		TR_24 = RG_rl_135 ;
	7'h7d :
		TR_24 = RG_rl_135 ;
	7'h7e :
		TR_24 = RG_rl_135 ;
	7'h7f :
		TR_24 = RG_rl_135 ;
	default :
		TR_24 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_4 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h01 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h02 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h03 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h04 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h05 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h06 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h07 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h08 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h09 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h0a :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h0b :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h0c :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h0d :
		TR_25 = 9'h000 ;	// line#=../rle.cpp:79
	7'h0e :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h0f :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h10 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h11 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h12 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h13 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h14 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h15 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h16 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h17 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h18 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h19 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h1a :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h1b :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h1c :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h1d :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h1e :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h1f :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h20 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h21 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h22 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h23 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h24 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h25 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h26 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h27 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h28 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h29 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h2a :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h2b :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h2c :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h2d :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h2e :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h2f :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h30 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h31 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h32 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h33 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h34 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h35 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h36 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h37 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h38 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h39 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h3a :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h3b :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h3c :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h3d :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h3e :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h3f :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h40 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h41 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h42 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h43 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h44 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h45 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h46 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h47 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h48 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h49 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h4a :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h4b :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h4c :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h4d :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h4e :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h4f :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h50 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h51 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h52 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h53 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h54 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h55 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h56 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h57 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h58 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h59 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h5a :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h5b :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h5c :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h5d :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h5e :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h5f :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h60 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h61 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h62 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h63 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h64 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h65 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h66 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h67 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h68 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h69 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h6a :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h6b :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h6c :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h6d :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h6e :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h6f :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h70 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h71 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h72 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h73 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h74 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h75 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h76 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h77 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h78 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h79 :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h7a :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h7b :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h7c :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h7d :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h7e :
		TR_25 = RG_quantized_block_rl_4 ;
	7'h7f :
		TR_25 = RG_quantized_block_rl_4 ;
	default :
		TR_25 = 9'hx ;
	endcase
always @ ( RG_rl_136 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_26 = RG_rl_136 ;
	7'h01 :
		TR_26 = RG_rl_136 ;
	7'h02 :
		TR_26 = RG_rl_136 ;
	7'h03 :
		TR_26 = RG_rl_136 ;
	7'h04 :
		TR_26 = RG_rl_136 ;
	7'h05 :
		TR_26 = RG_rl_136 ;
	7'h06 :
		TR_26 = RG_rl_136 ;
	7'h07 :
		TR_26 = RG_rl_136 ;
	7'h08 :
		TR_26 = RG_rl_136 ;
	7'h09 :
		TR_26 = RG_rl_136 ;
	7'h0a :
		TR_26 = RG_rl_136 ;
	7'h0b :
		TR_26 = RG_rl_136 ;
	7'h0c :
		TR_26 = RG_rl_136 ;
	7'h0d :
		TR_26 = RG_rl_136 ;
	7'h0e :
		TR_26 = 9'h000 ;	// line#=../rle.cpp:79
	7'h0f :
		TR_26 = RG_rl_136 ;
	7'h10 :
		TR_26 = RG_rl_136 ;
	7'h11 :
		TR_26 = RG_rl_136 ;
	7'h12 :
		TR_26 = RG_rl_136 ;
	7'h13 :
		TR_26 = RG_rl_136 ;
	7'h14 :
		TR_26 = RG_rl_136 ;
	7'h15 :
		TR_26 = RG_rl_136 ;
	7'h16 :
		TR_26 = RG_rl_136 ;
	7'h17 :
		TR_26 = RG_rl_136 ;
	7'h18 :
		TR_26 = RG_rl_136 ;
	7'h19 :
		TR_26 = RG_rl_136 ;
	7'h1a :
		TR_26 = RG_rl_136 ;
	7'h1b :
		TR_26 = RG_rl_136 ;
	7'h1c :
		TR_26 = RG_rl_136 ;
	7'h1d :
		TR_26 = RG_rl_136 ;
	7'h1e :
		TR_26 = RG_rl_136 ;
	7'h1f :
		TR_26 = RG_rl_136 ;
	7'h20 :
		TR_26 = RG_rl_136 ;
	7'h21 :
		TR_26 = RG_rl_136 ;
	7'h22 :
		TR_26 = RG_rl_136 ;
	7'h23 :
		TR_26 = RG_rl_136 ;
	7'h24 :
		TR_26 = RG_rl_136 ;
	7'h25 :
		TR_26 = RG_rl_136 ;
	7'h26 :
		TR_26 = RG_rl_136 ;
	7'h27 :
		TR_26 = RG_rl_136 ;
	7'h28 :
		TR_26 = RG_rl_136 ;
	7'h29 :
		TR_26 = RG_rl_136 ;
	7'h2a :
		TR_26 = RG_rl_136 ;
	7'h2b :
		TR_26 = RG_rl_136 ;
	7'h2c :
		TR_26 = RG_rl_136 ;
	7'h2d :
		TR_26 = RG_rl_136 ;
	7'h2e :
		TR_26 = RG_rl_136 ;
	7'h2f :
		TR_26 = RG_rl_136 ;
	7'h30 :
		TR_26 = RG_rl_136 ;
	7'h31 :
		TR_26 = RG_rl_136 ;
	7'h32 :
		TR_26 = RG_rl_136 ;
	7'h33 :
		TR_26 = RG_rl_136 ;
	7'h34 :
		TR_26 = RG_rl_136 ;
	7'h35 :
		TR_26 = RG_rl_136 ;
	7'h36 :
		TR_26 = RG_rl_136 ;
	7'h37 :
		TR_26 = RG_rl_136 ;
	7'h38 :
		TR_26 = RG_rl_136 ;
	7'h39 :
		TR_26 = RG_rl_136 ;
	7'h3a :
		TR_26 = RG_rl_136 ;
	7'h3b :
		TR_26 = RG_rl_136 ;
	7'h3c :
		TR_26 = RG_rl_136 ;
	7'h3d :
		TR_26 = RG_rl_136 ;
	7'h3e :
		TR_26 = RG_rl_136 ;
	7'h3f :
		TR_26 = RG_rl_136 ;
	7'h40 :
		TR_26 = RG_rl_136 ;
	7'h41 :
		TR_26 = RG_rl_136 ;
	7'h42 :
		TR_26 = RG_rl_136 ;
	7'h43 :
		TR_26 = RG_rl_136 ;
	7'h44 :
		TR_26 = RG_rl_136 ;
	7'h45 :
		TR_26 = RG_rl_136 ;
	7'h46 :
		TR_26 = RG_rl_136 ;
	7'h47 :
		TR_26 = RG_rl_136 ;
	7'h48 :
		TR_26 = RG_rl_136 ;
	7'h49 :
		TR_26 = RG_rl_136 ;
	7'h4a :
		TR_26 = RG_rl_136 ;
	7'h4b :
		TR_26 = RG_rl_136 ;
	7'h4c :
		TR_26 = RG_rl_136 ;
	7'h4d :
		TR_26 = RG_rl_136 ;
	7'h4e :
		TR_26 = RG_rl_136 ;
	7'h4f :
		TR_26 = RG_rl_136 ;
	7'h50 :
		TR_26 = RG_rl_136 ;
	7'h51 :
		TR_26 = RG_rl_136 ;
	7'h52 :
		TR_26 = RG_rl_136 ;
	7'h53 :
		TR_26 = RG_rl_136 ;
	7'h54 :
		TR_26 = RG_rl_136 ;
	7'h55 :
		TR_26 = RG_rl_136 ;
	7'h56 :
		TR_26 = RG_rl_136 ;
	7'h57 :
		TR_26 = RG_rl_136 ;
	7'h58 :
		TR_26 = RG_rl_136 ;
	7'h59 :
		TR_26 = RG_rl_136 ;
	7'h5a :
		TR_26 = RG_rl_136 ;
	7'h5b :
		TR_26 = RG_rl_136 ;
	7'h5c :
		TR_26 = RG_rl_136 ;
	7'h5d :
		TR_26 = RG_rl_136 ;
	7'h5e :
		TR_26 = RG_rl_136 ;
	7'h5f :
		TR_26 = RG_rl_136 ;
	7'h60 :
		TR_26 = RG_rl_136 ;
	7'h61 :
		TR_26 = RG_rl_136 ;
	7'h62 :
		TR_26 = RG_rl_136 ;
	7'h63 :
		TR_26 = RG_rl_136 ;
	7'h64 :
		TR_26 = RG_rl_136 ;
	7'h65 :
		TR_26 = RG_rl_136 ;
	7'h66 :
		TR_26 = RG_rl_136 ;
	7'h67 :
		TR_26 = RG_rl_136 ;
	7'h68 :
		TR_26 = RG_rl_136 ;
	7'h69 :
		TR_26 = RG_rl_136 ;
	7'h6a :
		TR_26 = RG_rl_136 ;
	7'h6b :
		TR_26 = RG_rl_136 ;
	7'h6c :
		TR_26 = RG_rl_136 ;
	7'h6d :
		TR_26 = RG_rl_136 ;
	7'h6e :
		TR_26 = RG_rl_136 ;
	7'h6f :
		TR_26 = RG_rl_136 ;
	7'h70 :
		TR_26 = RG_rl_136 ;
	7'h71 :
		TR_26 = RG_rl_136 ;
	7'h72 :
		TR_26 = RG_rl_136 ;
	7'h73 :
		TR_26 = RG_rl_136 ;
	7'h74 :
		TR_26 = RG_rl_136 ;
	7'h75 :
		TR_26 = RG_rl_136 ;
	7'h76 :
		TR_26 = RG_rl_136 ;
	7'h77 :
		TR_26 = RG_rl_136 ;
	7'h78 :
		TR_26 = RG_rl_136 ;
	7'h79 :
		TR_26 = RG_rl_136 ;
	7'h7a :
		TR_26 = RG_rl_136 ;
	7'h7b :
		TR_26 = RG_rl_136 ;
	7'h7c :
		TR_26 = RG_rl_136 ;
	7'h7d :
		TR_26 = RG_rl_136 ;
	7'h7e :
		TR_26 = RG_rl_136 ;
	7'h7f :
		TR_26 = RG_rl_136 ;
	default :
		TR_26 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_5 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h01 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h02 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h03 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h04 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h05 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h06 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h07 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h08 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h09 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h0a :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h0b :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h0c :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h0d :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h0e :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h0f :
		TR_27 = 9'h000 ;	// line#=../rle.cpp:79
	7'h10 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h11 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h12 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h13 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h14 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h15 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h16 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h17 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h18 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h19 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h1a :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h1b :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h1c :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h1d :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h1e :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h1f :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h20 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h21 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h22 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h23 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h24 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h25 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h26 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h27 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h28 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h29 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h2a :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h2b :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h2c :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h2d :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h2e :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h2f :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h30 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h31 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h32 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h33 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h34 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h35 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h36 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h37 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h38 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h39 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h3a :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h3b :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h3c :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h3d :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h3e :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h3f :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h40 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h41 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h42 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h43 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h44 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h45 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h46 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h47 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h48 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h49 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h4a :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h4b :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h4c :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h4d :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h4e :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h4f :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h50 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h51 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h52 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h53 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h54 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h55 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h56 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h57 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h58 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h59 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h5a :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h5b :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h5c :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h5d :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h5e :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h5f :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h60 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h61 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h62 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h63 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h64 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h65 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h66 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h67 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h68 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h69 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h6a :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h6b :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h6c :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h6d :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h6e :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h6f :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h70 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h71 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h72 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h73 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h74 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h75 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h76 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h77 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h78 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h79 :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h7a :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h7b :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h7c :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h7d :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h7e :
		TR_27 = RG_quantized_block_rl_5 ;
	7'h7f :
		TR_27 = RG_quantized_block_rl_5 ;
	default :
		TR_27 = 9'hx ;
	endcase
always @ ( RG_rl_137 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_28 = RG_rl_137 ;
	7'h01 :
		TR_28 = RG_rl_137 ;
	7'h02 :
		TR_28 = RG_rl_137 ;
	7'h03 :
		TR_28 = RG_rl_137 ;
	7'h04 :
		TR_28 = RG_rl_137 ;
	7'h05 :
		TR_28 = RG_rl_137 ;
	7'h06 :
		TR_28 = RG_rl_137 ;
	7'h07 :
		TR_28 = RG_rl_137 ;
	7'h08 :
		TR_28 = RG_rl_137 ;
	7'h09 :
		TR_28 = RG_rl_137 ;
	7'h0a :
		TR_28 = RG_rl_137 ;
	7'h0b :
		TR_28 = RG_rl_137 ;
	7'h0c :
		TR_28 = RG_rl_137 ;
	7'h0d :
		TR_28 = RG_rl_137 ;
	7'h0e :
		TR_28 = RG_rl_137 ;
	7'h0f :
		TR_28 = RG_rl_137 ;
	7'h10 :
		TR_28 = 9'h000 ;	// line#=../rle.cpp:79
	7'h11 :
		TR_28 = RG_rl_137 ;
	7'h12 :
		TR_28 = RG_rl_137 ;
	7'h13 :
		TR_28 = RG_rl_137 ;
	7'h14 :
		TR_28 = RG_rl_137 ;
	7'h15 :
		TR_28 = RG_rl_137 ;
	7'h16 :
		TR_28 = RG_rl_137 ;
	7'h17 :
		TR_28 = RG_rl_137 ;
	7'h18 :
		TR_28 = RG_rl_137 ;
	7'h19 :
		TR_28 = RG_rl_137 ;
	7'h1a :
		TR_28 = RG_rl_137 ;
	7'h1b :
		TR_28 = RG_rl_137 ;
	7'h1c :
		TR_28 = RG_rl_137 ;
	7'h1d :
		TR_28 = RG_rl_137 ;
	7'h1e :
		TR_28 = RG_rl_137 ;
	7'h1f :
		TR_28 = RG_rl_137 ;
	7'h20 :
		TR_28 = RG_rl_137 ;
	7'h21 :
		TR_28 = RG_rl_137 ;
	7'h22 :
		TR_28 = RG_rl_137 ;
	7'h23 :
		TR_28 = RG_rl_137 ;
	7'h24 :
		TR_28 = RG_rl_137 ;
	7'h25 :
		TR_28 = RG_rl_137 ;
	7'h26 :
		TR_28 = RG_rl_137 ;
	7'h27 :
		TR_28 = RG_rl_137 ;
	7'h28 :
		TR_28 = RG_rl_137 ;
	7'h29 :
		TR_28 = RG_rl_137 ;
	7'h2a :
		TR_28 = RG_rl_137 ;
	7'h2b :
		TR_28 = RG_rl_137 ;
	7'h2c :
		TR_28 = RG_rl_137 ;
	7'h2d :
		TR_28 = RG_rl_137 ;
	7'h2e :
		TR_28 = RG_rl_137 ;
	7'h2f :
		TR_28 = RG_rl_137 ;
	7'h30 :
		TR_28 = RG_rl_137 ;
	7'h31 :
		TR_28 = RG_rl_137 ;
	7'h32 :
		TR_28 = RG_rl_137 ;
	7'h33 :
		TR_28 = RG_rl_137 ;
	7'h34 :
		TR_28 = RG_rl_137 ;
	7'h35 :
		TR_28 = RG_rl_137 ;
	7'h36 :
		TR_28 = RG_rl_137 ;
	7'h37 :
		TR_28 = RG_rl_137 ;
	7'h38 :
		TR_28 = RG_rl_137 ;
	7'h39 :
		TR_28 = RG_rl_137 ;
	7'h3a :
		TR_28 = RG_rl_137 ;
	7'h3b :
		TR_28 = RG_rl_137 ;
	7'h3c :
		TR_28 = RG_rl_137 ;
	7'h3d :
		TR_28 = RG_rl_137 ;
	7'h3e :
		TR_28 = RG_rl_137 ;
	7'h3f :
		TR_28 = RG_rl_137 ;
	7'h40 :
		TR_28 = RG_rl_137 ;
	7'h41 :
		TR_28 = RG_rl_137 ;
	7'h42 :
		TR_28 = RG_rl_137 ;
	7'h43 :
		TR_28 = RG_rl_137 ;
	7'h44 :
		TR_28 = RG_rl_137 ;
	7'h45 :
		TR_28 = RG_rl_137 ;
	7'h46 :
		TR_28 = RG_rl_137 ;
	7'h47 :
		TR_28 = RG_rl_137 ;
	7'h48 :
		TR_28 = RG_rl_137 ;
	7'h49 :
		TR_28 = RG_rl_137 ;
	7'h4a :
		TR_28 = RG_rl_137 ;
	7'h4b :
		TR_28 = RG_rl_137 ;
	7'h4c :
		TR_28 = RG_rl_137 ;
	7'h4d :
		TR_28 = RG_rl_137 ;
	7'h4e :
		TR_28 = RG_rl_137 ;
	7'h4f :
		TR_28 = RG_rl_137 ;
	7'h50 :
		TR_28 = RG_rl_137 ;
	7'h51 :
		TR_28 = RG_rl_137 ;
	7'h52 :
		TR_28 = RG_rl_137 ;
	7'h53 :
		TR_28 = RG_rl_137 ;
	7'h54 :
		TR_28 = RG_rl_137 ;
	7'h55 :
		TR_28 = RG_rl_137 ;
	7'h56 :
		TR_28 = RG_rl_137 ;
	7'h57 :
		TR_28 = RG_rl_137 ;
	7'h58 :
		TR_28 = RG_rl_137 ;
	7'h59 :
		TR_28 = RG_rl_137 ;
	7'h5a :
		TR_28 = RG_rl_137 ;
	7'h5b :
		TR_28 = RG_rl_137 ;
	7'h5c :
		TR_28 = RG_rl_137 ;
	7'h5d :
		TR_28 = RG_rl_137 ;
	7'h5e :
		TR_28 = RG_rl_137 ;
	7'h5f :
		TR_28 = RG_rl_137 ;
	7'h60 :
		TR_28 = RG_rl_137 ;
	7'h61 :
		TR_28 = RG_rl_137 ;
	7'h62 :
		TR_28 = RG_rl_137 ;
	7'h63 :
		TR_28 = RG_rl_137 ;
	7'h64 :
		TR_28 = RG_rl_137 ;
	7'h65 :
		TR_28 = RG_rl_137 ;
	7'h66 :
		TR_28 = RG_rl_137 ;
	7'h67 :
		TR_28 = RG_rl_137 ;
	7'h68 :
		TR_28 = RG_rl_137 ;
	7'h69 :
		TR_28 = RG_rl_137 ;
	7'h6a :
		TR_28 = RG_rl_137 ;
	7'h6b :
		TR_28 = RG_rl_137 ;
	7'h6c :
		TR_28 = RG_rl_137 ;
	7'h6d :
		TR_28 = RG_rl_137 ;
	7'h6e :
		TR_28 = RG_rl_137 ;
	7'h6f :
		TR_28 = RG_rl_137 ;
	7'h70 :
		TR_28 = RG_rl_137 ;
	7'h71 :
		TR_28 = RG_rl_137 ;
	7'h72 :
		TR_28 = RG_rl_137 ;
	7'h73 :
		TR_28 = RG_rl_137 ;
	7'h74 :
		TR_28 = RG_rl_137 ;
	7'h75 :
		TR_28 = RG_rl_137 ;
	7'h76 :
		TR_28 = RG_rl_137 ;
	7'h77 :
		TR_28 = RG_rl_137 ;
	7'h78 :
		TR_28 = RG_rl_137 ;
	7'h79 :
		TR_28 = RG_rl_137 ;
	7'h7a :
		TR_28 = RG_rl_137 ;
	7'h7b :
		TR_28 = RG_rl_137 ;
	7'h7c :
		TR_28 = RG_rl_137 ;
	7'h7d :
		TR_28 = RG_rl_137 ;
	7'h7e :
		TR_28 = RG_rl_137 ;
	7'h7f :
		TR_28 = RG_rl_137 ;
	default :
		TR_28 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_6 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h01 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h02 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h03 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h04 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h05 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h06 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h07 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h08 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h09 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h0a :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h0b :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h0c :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h0d :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h0e :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h0f :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h10 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h11 :
		TR_29 = 9'h000 ;	// line#=../rle.cpp:79
	7'h12 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h13 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h14 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h15 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h16 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h17 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h18 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h19 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h1a :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h1b :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h1c :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h1d :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h1e :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h1f :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h20 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h21 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h22 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h23 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h24 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h25 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h26 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h27 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h28 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h29 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h2a :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h2b :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h2c :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h2d :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h2e :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h2f :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h30 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h31 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h32 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h33 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h34 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h35 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h36 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h37 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h38 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h39 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h3a :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h3b :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h3c :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h3d :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h3e :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h3f :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h40 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h41 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h42 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h43 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h44 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h45 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h46 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h47 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h48 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h49 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h4a :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h4b :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h4c :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h4d :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h4e :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h4f :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h50 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h51 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h52 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h53 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h54 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h55 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h56 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h57 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h58 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h59 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h5a :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h5b :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h5c :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h5d :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h5e :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h5f :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h60 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h61 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h62 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h63 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h64 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h65 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h66 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h67 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h68 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h69 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h6a :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h6b :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h6c :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h6d :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h6e :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h6f :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h70 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h71 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h72 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h73 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h74 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h75 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h76 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h77 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h78 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h79 :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h7a :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h7b :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h7c :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h7d :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h7e :
		TR_29 = RG_quantized_block_rl_6 ;
	7'h7f :
		TR_29 = RG_quantized_block_rl_6 ;
	default :
		TR_29 = 9'hx ;
	endcase
always @ ( RG_rl_138 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_30 = RG_rl_138 ;
	7'h01 :
		TR_30 = RG_rl_138 ;
	7'h02 :
		TR_30 = RG_rl_138 ;
	7'h03 :
		TR_30 = RG_rl_138 ;
	7'h04 :
		TR_30 = RG_rl_138 ;
	7'h05 :
		TR_30 = RG_rl_138 ;
	7'h06 :
		TR_30 = RG_rl_138 ;
	7'h07 :
		TR_30 = RG_rl_138 ;
	7'h08 :
		TR_30 = RG_rl_138 ;
	7'h09 :
		TR_30 = RG_rl_138 ;
	7'h0a :
		TR_30 = RG_rl_138 ;
	7'h0b :
		TR_30 = RG_rl_138 ;
	7'h0c :
		TR_30 = RG_rl_138 ;
	7'h0d :
		TR_30 = RG_rl_138 ;
	7'h0e :
		TR_30 = RG_rl_138 ;
	7'h0f :
		TR_30 = RG_rl_138 ;
	7'h10 :
		TR_30 = RG_rl_138 ;
	7'h11 :
		TR_30 = RG_rl_138 ;
	7'h12 :
		TR_30 = 9'h000 ;	// line#=../rle.cpp:79
	7'h13 :
		TR_30 = RG_rl_138 ;
	7'h14 :
		TR_30 = RG_rl_138 ;
	7'h15 :
		TR_30 = RG_rl_138 ;
	7'h16 :
		TR_30 = RG_rl_138 ;
	7'h17 :
		TR_30 = RG_rl_138 ;
	7'h18 :
		TR_30 = RG_rl_138 ;
	7'h19 :
		TR_30 = RG_rl_138 ;
	7'h1a :
		TR_30 = RG_rl_138 ;
	7'h1b :
		TR_30 = RG_rl_138 ;
	7'h1c :
		TR_30 = RG_rl_138 ;
	7'h1d :
		TR_30 = RG_rl_138 ;
	7'h1e :
		TR_30 = RG_rl_138 ;
	7'h1f :
		TR_30 = RG_rl_138 ;
	7'h20 :
		TR_30 = RG_rl_138 ;
	7'h21 :
		TR_30 = RG_rl_138 ;
	7'h22 :
		TR_30 = RG_rl_138 ;
	7'h23 :
		TR_30 = RG_rl_138 ;
	7'h24 :
		TR_30 = RG_rl_138 ;
	7'h25 :
		TR_30 = RG_rl_138 ;
	7'h26 :
		TR_30 = RG_rl_138 ;
	7'h27 :
		TR_30 = RG_rl_138 ;
	7'h28 :
		TR_30 = RG_rl_138 ;
	7'h29 :
		TR_30 = RG_rl_138 ;
	7'h2a :
		TR_30 = RG_rl_138 ;
	7'h2b :
		TR_30 = RG_rl_138 ;
	7'h2c :
		TR_30 = RG_rl_138 ;
	7'h2d :
		TR_30 = RG_rl_138 ;
	7'h2e :
		TR_30 = RG_rl_138 ;
	7'h2f :
		TR_30 = RG_rl_138 ;
	7'h30 :
		TR_30 = RG_rl_138 ;
	7'h31 :
		TR_30 = RG_rl_138 ;
	7'h32 :
		TR_30 = RG_rl_138 ;
	7'h33 :
		TR_30 = RG_rl_138 ;
	7'h34 :
		TR_30 = RG_rl_138 ;
	7'h35 :
		TR_30 = RG_rl_138 ;
	7'h36 :
		TR_30 = RG_rl_138 ;
	7'h37 :
		TR_30 = RG_rl_138 ;
	7'h38 :
		TR_30 = RG_rl_138 ;
	7'h39 :
		TR_30 = RG_rl_138 ;
	7'h3a :
		TR_30 = RG_rl_138 ;
	7'h3b :
		TR_30 = RG_rl_138 ;
	7'h3c :
		TR_30 = RG_rl_138 ;
	7'h3d :
		TR_30 = RG_rl_138 ;
	7'h3e :
		TR_30 = RG_rl_138 ;
	7'h3f :
		TR_30 = RG_rl_138 ;
	7'h40 :
		TR_30 = RG_rl_138 ;
	7'h41 :
		TR_30 = RG_rl_138 ;
	7'h42 :
		TR_30 = RG_rl_138 ;
	7'h43 :
		TR_30 = RG_rl_138 ;
	7'h44 :
		TR_30 = RG_rl_138 ;
	7'h45 :
		TR_30 = RG_rl_138 ;
	7'h46 :
		TR_30 = RG_rl_138 ;
	7'h47 :
		TR_30 = RG_rl_138 ;
	7'h48 :
		TR_30 = RG_rl_138 ;
	7'h49 :
		TR_30 = RG_rl_138 ;
	7'h4a :
		TR_30 = RG_rl_138 ;
	7'h4b :
		TR_30 = RG_rl_138 ;
	7'h4c :
		TR_30 = RG_rl_138 ;
	7'h4d :
		TR_30 = RG_rl_138 ;
	7'h4e :
		TR_30 = RG_rl_138 ;
	7'h4f :
		TR_30 = RG_rl_138 ;
	7'h50 :
		TR_30 = RG_rl_138 ;
	7'h51 :
		TR_30 = RG_rl_138 ;
	7'h52 :
		TR_30 = RG_rl_138 ;
	7'h53 :
		TR_30 = RG_rl_138 ;
	7'h54 :
		TR_30 = RG_rl_138 ;
	7'h55 :
		TR_30 = RG_rl_138 ;
	7'h56 :
		TR_30 = RG_rl_138 ;
	7'h57 :
		TR_30 = RG_rl_138 ;
	7'h58 :
		TR_30 = RG_rl_138 ;
	7'h59 :
		TR_30 = RG_rl_138 ;
	7'h5a :
		TR_30 = RG_rl_138 ;
	7'h5b :
		TR_30 = RG_rl_138 ;
	7'h5c :
		TR_30 = RG_rl_138 ;
	7'h5d :
		TR_30 = RG_rl_138 ;
	7'h5e :
		TR_30 = RG_rl_138 ;
	7'h5f :
		TR_30 = RG_rl_138 ;
	7'h60 :
		TR_30 = RG_rl_138 ;
	7'h61 :
		TR_30 = RG_rl_138 ;
	7'h62 :
		TR_30 = RG_rl_138 ;
	7'h63 :
		TR_30 = RG_rl_138 ;
	7'h64 :
		TR_30 = RG_rl_138 ;
	7'h65 :
		TR_30 = RG_rl_138 ;
	7'h66 :
		TR_30 = RG_rl_138 ;
	7'h67 :
		TR_30 = RG_rl_138 ;
	7'h68 :
		TR_30 = RG_rl_138 ;
	7'h69 :
		TR_30 = RG_rl_138 ;
	7'h6a :
		TR_30 = RG_rl_138 ;
	7'h6b :
		TR_30 = RG_rl_138 ;
	7'h6c :
		TR_30 = RG_rl_138 ;
	7'h6d :
		TR_30 = RG_rl_138 ;
	7'h6e :
		TR_30 = RG_rl_138 ;
	7'h6f :
		TR_30 = RG_rl_138 ;
	7'h70 :
		TR_30 = RG_rl_138 ;
	7'h71 :
		TR_30 = RG_rl_138 ;
	7'h72 :
		TR_30 = RG_rl_138 ;
	7'h73 :
		TR_30 = RG_rl_138 ;
	7'h74 :
		TR_30 = RG_rl_138 ;
	7'h75 :
		TR_30 = RG_rl_138 ;
	7'h76 :
		TR_30 = RG_rl_138 ;
	7'h77 :
		TR_30 = RG_rl_138 ;
	7'h78 :
		TR_30 = RG_rl_138 ;
	7'h79 :
		TR_30 = RG_rl_138 ;
	7'h7a :
		TR_30 = RG_rl_138 ;
	7'h7b :
		TR_30 = RG_rl_138 ;
	7'h7c :
		TR_30 = RG_rl_138 ;
	7'h7d :
		TR_30 = RG_rl_138 ;
	7'h7e :
		TR_30 = RG_rl_138 ;
	7'h7f :
		TR_30 = RG_rl_138 ;
	default :
		TR_30 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_7 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h01 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h02 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h03 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h04 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h05 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h06 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h07 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h08 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h09 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h0a :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h0b :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h0c :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h0d :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h0e :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h0f :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h10 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h11 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h12 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h13 :
		TR_31 = 9'h000 ;	// line#=../rle.cpp:79
	7'h14 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h15 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h16 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h17 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h18 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h19 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h1a :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h1b :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h1c :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h1d :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h1e :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h1f :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h20 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h21 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h22 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h23 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h24 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h25 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h26 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h27 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h28 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h29 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h2a :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h2b :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h2c :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h2d :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h2e :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h2f :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h30 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h31 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h32 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h33 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h34 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h35 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h36 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h37 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h38 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h39 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h3a :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h3b :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h3c :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h3d :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h3e :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h3f :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h40 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h41 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h42 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h43 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h44 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h45 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h46 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h47 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h48 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h49 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h4a :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h4b :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h4c :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h4d :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h4e :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h4f :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h50 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h51 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h52 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h53 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h54 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h55 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h56 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h57 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h58 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h59 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h5a :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h5b :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h5c :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h5d :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h5e :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h5f :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h60 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h61 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h62 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h63 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h64 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h65 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h66 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h67 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h68 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h69 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h6a :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h6b :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h6c :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h6d :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h6e :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h6f :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h70 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h71 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h72 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h73 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h74 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h75 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h76 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h77 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h78 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h79 :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h7a :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h7b :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h7c :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h7d :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h7e :
		TR_31 = RG_quantized_block_rl_7 ;
	7'h7f :
		TR_31 = RG_quantized_block_rl_7 ;
	default :
		TR_31 = 9'hx ;
	endcase
always @ ( RG_rl_139 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_32 = RG_rl_139 ;
	7'h01 :
		TR_32 = RG_rl_139 ;
	7'h02 :
		TR_32 = RG_rl_139 ;
	7'h03 :
		TR_32 = RG_rl_139 ;
	7'h04 :
		TR_32 = RG_rl_139 ;
	7'h05 :
		TR_32 = RG_rl_139 ;
	7'h06 :
		TR_32 = RG_rl_139 ;
	7'h07 :
		TR_32 = RG_rl_139 ;
	7'h08 :
		TR_32 = RG_rl_139 ;
	7'h09 :
		TR_32 = RG_rl_139 ;
	7'h0a :
		TR_32 = RG_rl_139 ;
	7'h0b :
		TR_32 = RG_rl_139 ;
	7'h0c :
		TR_32 = RG_rl_139 ;
	7'h0d :
		TR_32 = RG_rl_139 ;
	7'h0e :
		TR_32 = RG_rl_139 ;
	7'h0f :
		TR_32 = RG_rl_139 ;
	7'h10 :
		TR_32 = RG_rl_139 ;
	7'h11 :
		TR_32 = RG_rl_139 ;
	7'h12 :
		TR_32 = RG_rl_139 ;
	7'h13 :
		TR_32 = RG_rl_139 ;
	7'h14 :
		TR_32 = 9'h000 ;	// line#=../rle.cpp:79
	7'h15 :
		TR_32 = RG_rl_139 ;
	7'h16 :
		TR_32 = RG_rl_139 ;
	7'h17 :
		TR_32 = RG_rl_139 ;
	7'h18 :
		TR_32 = RG_rl_139 ;
	7'h19 :
		TR_32 = RG_rl_139 ;
	7'h1a :
		TR_32 = RG_rl_139 ;
	7'h1b :
		TR_32 = RG_rl_139 ;
	7'h1c :
		TR_32 = RG_rl_139 ;
	7'h1d :
		TR_32 = RG_rl_139 ;
	7'h1e :
		TR_32 = RG_rl_139 ;
	7'h1f :
		TR_32 = RG_rl_139 ;
	7'h20 :
		TR_32 = RG_rl_139 ;
	7'h21 :
		TR_32 = RG_rl_139 ;
	7'h22 :
		TR_32 = RG_rl_139 ;
	7'h23 :
		TR_32 = RG_rl_139 ;
	7'h24 :
		TR_32 = RG_rl_139 ;
	7'h25 :
		TR_32 = RG_rl_139 ;
	7'h26 :
		TR_32 = RG_rl_139 ;
	7'h27 :
		TR_32 = RG_rl_139 ;
	7'h28 :
		TR_32 = RG_rl_139 ;
	7'h29 :
		TR_32 = RG_rl_139 ;
	7'h2a :
		TR_32 = RG_rl_139 ;
	7'h2b :
		TR_32 = RG_rl_139 ;
	7'h2c :
		TR_32 = RG_rl_139 ;
	7'h2d :
		TR_32 = RG_rl_139 ;
	7'h2e :
		TR_32 = RG_rl_139 ;
	7'h2f :
		TR_32 = RG_rl_139 ;
	7'h30 :
		TR_32 = RG_rl_139 ;
	7'h31 :
		TR_32 = RG_rl_139 ;
	7'h32 :
		TR_32 = RG_rl_139 ;
	7'h33 :
		TR_32 = RG_rl_139 ;
	7'h34 :
		TR_32 = RG_rl_139 ;
	7'h35 :
		TR_32 = RG_rl_139 ;
	7'h36 :
		TR_32 = RG_rl_139 ;
	7'h37 :
		TR_32 = RG_rl_139 ;
	7'h38 :
		TR_32 = RG_rl_139 ;
	7'h39 :
		TR_32 = RG_rl_139 ;
	7'h3a :
		TR_32 = RG_rl_139 ;
	7'h3b :
		TR_32 = RG_rl_139 ;
	7'h3c :
		TR_32 = RG_rl_139 ;
	7'h3d :
		TR_32 = RG_rl_139 ;
	7'h3e :
		TR_32 = RG_rl_139 ;
	7'h3f :
		TR_32 = RG_rl_139 ;
	7'h40 :
		TR_32 = RG_rl_139 ;
	7'h41 :
		TR_32 = RG_rl_139 ;
	7'h42 :
		TR_32 = RG_rl_139 ;
	7'h43 :
		TR_32 = RG_rl_139 ;
	7'h44 :
		TR_32 = RG_rl_139 ;
	7'h45 :
		TR_32 = RG_rl_139 ;
	7'h46 :
		TR_32 = RG_rl_139 ;
	7'h47 :
		TR_32 = RG_rl_139 ;
	7'h48 :
		TR_32 = RG_rl_139 ;
	7'h49 :
		TR_32 = RG_rl_139 ;
	7'h4a :
		TR_32 = RG_rl_139 ;
	7'h4b :
		TR_32 = RG_rl_139 ;
	7'h4c :
		TR_32 = RG_rl_139 ;
	7'h4d :
		TR_32 = RG_rl_139 ;
	7'h4e :
		TR_32 = RG_rl_139 ;
	7'h4f :
		TR_32 = RG_rl_139 ;
	7'h50 :
		TR_32 = RG_rl_139 ;
	7'h51 :
		TR_32 = RG_rl_139 ;
	7'h52 :
		TR_32 = RG_rl_139 ;
	7'h53 :
		TR_32 = RG_rl_139 ;
	7'h54 :
		TR_32 = RG_rl_139 ;
	7'h55 :
		TR_32 = RG_rl_139 ;
	7'h56 :
		TR_32 = RG_rl_139 ;
	7'h57 :
		TR_32 = RG_rl_139 ;
	7'h58 :
		TR_32 = RG_rl_139 ;
	7'h59 :
		TR_32 = RG_rl_139 ;
	7'h5a :
		TR_32 = RG_rl_139 ;
	7'h5b :
		TR_32 = RG_rl_139 ;
	7'h5c :
		TR_32 = RG_rl_139 ;
	7'h5d :
		TR_32 = RG_rl_139 ;
	7'h5e :
		TR_32 = RG_rl_139 ;
	7'h5f :
		TR_32 = RG_rl_139 ;
	7'h60 :
		TR_32 = RG_rl_139 ;
	7'h61 :
		TR_32 = RG_rl_139 ;
	7'h62 :
		TR_32 = RG_rl_139 ;
	7'h63 :
		TR_32 = RG_rl_139 ;
	7'h64 :
		TR_32 = RG_rl_139 ;
	7'h65 :
		TR_32 = RG_rl_139 ;
	7'h66 :
		TR_32 = RG_rl_139 ;
	7'h67 :
		TR_32 = RG_rl_139 ;
	7'h68 :
		TR_32 = RG_rl_139 ;
	7'h69 :
		TR_32 = RG_rl_139 ;
	7'h6a :
		TR_32 = RG_rl_139 ;
	7'h6b :
		TR_32 = RG_rl_139 ;
	7'h6c :
		TR_32 = RG_rl_139 ;
	7'h6d :
		TR_32 = RG_rl_139 ;
	7'h6e :
		TR_32 = RG_rl_139 ;
	7'h6f :
		TR_32 = RG_rl_139 ;
	7'h70 :
		TR_32 = RG_rl_139 ;
	7'h71 :
		TR_32 = RG_rl_139 ;
	7'h72 :
		TR_32 = RG_rl_139 ;
	7'h73 :
		TR_32 = RG_rl_139 ;
	7'h74 :
		TR_32 = RG_rl_139 ;
	7'h75 :
		TR_32 = RG_rl_139 ;
	7'h76 :
		TR_32 = RG_rl_139 ;
	7'h77 :
		TR_32 = RG_rl_139 ;
	7'h78 :
		TR_32 = RG_rl_139 ;
	7'h79 :
		TR_32 = RG_rl_139 ;
	7'h7a :
		TR_32 = RG_rl_139 ;
	7'h7b :
		TR_32 = RG_rl_139 ;
	7'h7c :
		TR_32 = RG_rl_139 ;
	7'h7d :
		TR_32 = RG_rl_139 ;
	7'h7e :
		TR_32 = RG_rl_139 ;
	7'h7f :
		TR_32 = RG_rl_139 ;
	default :
		TR_32 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_8 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h01 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h02 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h03 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h04 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h05 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h06 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h07 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h08 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h09 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h0a :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h0b :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h0c :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h0d :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h0e :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h0f :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h10 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h11 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h12 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h13 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h14 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h15 :
		TR_33 = 9'h000 ;	// line#=../rle.cpp:79
	7'h16 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h17 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h18 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h19 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h1a :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h1b :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h1c :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h1d :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h1e :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h1f :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h20 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h21 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h22 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h23 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h24 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h25 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h26 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h27 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h28 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h29 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h2a :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h2b :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h2c :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h2d :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h2e :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h2f :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h30 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h31 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h32 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h33 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h34 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h35 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h36 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h37 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h38 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h39 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h3a :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h3b :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h3c :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h3d :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h3e :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h3f :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h40 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h41 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h42 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h43 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h44 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h45 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h46 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h47 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h48 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h49 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h4a :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h4b :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h4c :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h4d :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h4e :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h4f :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h50 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h51 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h52 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h53 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h54 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h55 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h56 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h57 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h58 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h59 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h5a :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h5b :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h5c :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h5d :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h5e :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h5f :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h60 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h61 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h62 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h63 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h64 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h65 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h66 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h67 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h68 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h69 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h6a :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h6b :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h6c :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h6d :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h6e :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h6f :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h70 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h71 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h72 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h73 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h74 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h75 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h76 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h77 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h78 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h79 :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h7a :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h7b :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h7c :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h7d :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h7e :
		TR_33 = RG_quantized_block_rl_8 ;
	7'h7f :
		TR_33 = RG_quantized_block_rl_8 ;
	default :
		TR_33 = 9'hx ;
	endcase
always @ ( RG_rl_140 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_34 = RG_rl_140 ;
	7'h01 :
		TR_34 = RG_rl_140 ;
	7'h02 :
		TR_34 = RG_rl_140 ;
	7'h03 :
		TR_34 = RG_rl_140 ;
	7'h04 :
		TR_34 = RG_rl_140 ;
	7'h05 :
		TR_34 = RG_rl_140 ;
	7'h06 :
		TR_34 = RG_rl_140 ;
	7'h07 :
		TR_34 = RG_rl_140 ;
	7'h08 :
		TR_34 = RG_rl_140 ;
	7'h09 :
		TR_34 = RG_rl_140 ;
	7'h0a :
		TR_34 = RG_rl_140 ;
	7'h0b :
		TR_34 = RG_rl_140 ;
	7'h0c :
		TR_34 = RG_rl_140 ;
	7'h0d :
		TR_34 = RG_rl_140 ;
	7'h0e :
		TR_34 = RG_rl_140 ;
	7'h0f :
		TR_34 = RG_rl_140 ;
	7'h10 :
		TR_34 = RG_rl_140 ;
	7'h11 :
		TR_34 = RG_rl_140 ;
	7'h12 :
		TR_34 = RG_rl_140 ;
	7'h13 :
		TR_34 = RG_rl_140 ;
	7'h14 :
		TR_34 = RG_rl_140 ;
	7'h15 :
		TR_34 = RG_rl_140 ;
	7'h16 :
		TR_34 = 9'h000 ;	// line#=../rle.cpp:79
	7'h17 :
		TR_34 = RG_rl_140 ;
	7'h18 :
		TR_34 = RG_rl_140 ;
	7'h19 :
		TR_34 = RG_rl_140 ;
	7'h1a :
		TR_34 = RG_rl_140 ;
	7'h1b :
		TR_34 = RG_rl_140 ;
	7'h1c :
		TR_34 = RG_rl_140 ;
	7'h1d :
		TR_34 = RG_rl_140 ;
	7'h1e :
		TR_34 = RG_rl_140 ;
	7'h1f :
		TR_34 = RG_rl_140 ;
	7'h20 :
		TR_34 = RG_rl_140 ;
	7'h21 :
		TR_34 = RG_rl_140 ;
	7'h22 :
		TR_34 = RG_rl_140 ;
	7'h23 :
		TR_34 = RG_rl_140 ;
	7'h24 :
		TR_34 = RG_rl_140 ;
	7'h25 :
		TR_34 = RG_rl_140 ;
	7'h26 :
		TR_34 = RG_rl_140 ;
	7'h27 :
		TR_34 = RG_rl_140 ;
	7'h28 :
		TR_34 = RG_rl_140 ;
	7'h29 :
		TR_34 = RG_rl_140 ;
	7'h2a :
		TR_34 = RG_rl_140 ;
	7'h2b :
		TR_34 = RG_rl_140 ;
	7'h2c :
		TR_34 = RG_rl_140 ;
	7'h2d :
		TR_34 = RG_rl_140 ;
	7'h2e :
		TR_34 = RG_rl_140 ;
	7'h2f :
		TR_34 = RG_rl_140 ;
	7'h30 :
		TR_34 = RG_rl_140 ;
	7'h31 :
		TR_34 = RG_rl_140 ;
	7'h32 :
		TR_34 = RG_rl_140 ;
	7'h33 :
		TR_34 = RG_rl_140 ;
	7'h34 :
		TR_34 = RG_rl_140 ;
	7'h35 :
		TR_34 = RG_rl_140 ;
	7'h36 :
		TR_34 = RG_rl_140 ;
	7'h37 :
		TR_34 = RG_rl_140 ;
	7'h38 :
		TR_34 = RG_rl_140 ;
	7'h39 :
		TR_34 = RG_rl_140 ;
	7'h3a :
		TR_34 = RG_rl_140 ;
	7'h3b :
		TR_34 = RG_rl_140 ;
	7'h3c :
		TR_34 = RG_rl_140 ;
	7'h3d :
		TR_34 = RG_rl_140 ;
	7'h3e :
		TR_34 = RG_rl_140 ;
	7'h3f :
		TR_34 = RG_rl_140 ;
	7'h40 :
		TR_34 = RG_rl_140 ;
	7'h41 :
		TR_34 = RG_rl_140 ;
	7'h42 :
		TR_34 = RG_rl_140 ;
	7'h43 :
		TR_34 = RG_rl_140 ;
	7'h44 :
		TR_34 = RG_rl_140 ;
	7'h45 :
		TR_34 = RG_rl_140 ;
	7'h46 :
		TR_34 = RG_rl_140 ;
	7'h47 :
		TR_34 = RG_rl_140 ;
	7'h48 :
		TR_34 = RG_rl_140 ;
	7'h49 :
		TR_34 = RG_rl_140 ;
	7'h4a :
		TR_34 = RG_rl_140 ;
	7'h4b :
		TR_34 = RG_rl_140 ;
	7'h4c :
		TR_34 = RG_rl_140 ;
	7'h4d :
		TR_34 = RG_rl_140 ;
	7'h4e :
		TR_34 = RG_rl_140 ;
	7'h4f :
		TR_34 = RG_rl_140 ;
	7'h50 :
		TR_34 = RG_rl_140 ;
	7'h51 :
		TR_34 = RG_rl_140 ;
	7'h52 :
		TR_34 = RG_rl_140 ;
	7'h53 :
		TR_34 = RG_rl_140 ;
	7'h54 :
		TR_34 = RG_rl_140 ;
	7'h55 :
		TR_34 = RG_rl_140 ;
	7'h56 :
		TR_34 = RG_rl_140 ;
	7'h57 :
		TR_34 = RG_rl_140 ;
	7'h58 :
		TR_34 = RG_rl_140 ;
	7'h59 :
		TR_34 = RG_rl_140 ;
	7'h5a :
		TR_34 = RG_rl_140 ;
	7'h5b :
		TR_34 = RG_rl_140 ;
	7'h5c :
		TR_34 = RG_rl_140 ;
	7'h5d :
		TR_34 = RG_rl_140 ;
	7'h5e :
		TR_34 = RG_rl_140 ;
	7'h5f :
		TR_34 = RG_rl_140 ;
	7'h60 :
		TR_34 = RG_rl_140 ;
	7'h61 :
		TR_34 = RG_rl_140 ;
	7'h62 :
		TR_34 = RG_rl_140 ;
	7'h63 :
		TR_34 = RG_rl_140 ;
	7'h64 :
		TR_34 = RG_rl_140 ;
	7'h65 :
		TR_34 = RG_rl_140 ;
	7'h66 :
		TR_34 = RG_rl_140 ;
	7'h67 :
		TR_34 = RG_rl_140 ;
	7'h68 :
		TR_34 = RG_rl_140 ;
	7'h69 :
		TR_34 = RG_rl_140 ;
	7'h6a :
		TR_34 = RG_rl_140 ;
	7'h6b :
		TR_34 = RG_rl_140 ;
	7'h6c :
		TR_34 = RG_rl_140 ;
	7'h6d :
		TR_34 = RG_rl_140 ;
	7'h6e :
		TR_34 = RG_rl_140 ;
	7'h6f :
		TR_34 = RG_rl_140 ;
	7'h70 :
		TR_34 = RG_rl_140 ;
	7'h71 :
		TR_34 = RG_rl_140 ;
	7'h72 :
		TR_34 = RG_rl_140 ;
	7'h73 :
		TR_34 = RG_rl_140 ;
	7'h74 :
		TR_34 = RG_rl_140 ;
	7'h75 :
		TR_34 = RG_rl_140 ;
	7'h76 :
		TR_34 = RG_rl_140 ;
	7'h77 :
		TR_34 = RG_rl_140 ;
	7'h78 :
		TR_34 = RG_rl_140 ;
	7'h79 :
		TR_34 = RG_rl_140 ;
	7'h7a :
		TR_34 = RG_rl_140 ;
	7'h7b :
		TR_34 = RG_rl_140 ;
	7'h7c :
		TR_34 = RG_rl_140 ;
	7'h7d :
		TR_34 = RG_rl_140 ;
	7'h7e :
		TR_34 = RG_rl_140 ;
	7'h7f :
		TR_34 = RG_rl_140 ;
	default :
		TR_34 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_9 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h01 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h02 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h03 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h04 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h05 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h06 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h07 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h08 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h09 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h0a :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h0b :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h0c :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h0d :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h0e :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h0f :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h10 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h11 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h12 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h13 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h14 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h15 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h16 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h17 :
		TR_35 = 9'h000 ;	// line#=../rle.cpp:79
	7'h18 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h19 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h1a :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h1b :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h1c :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h1d :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h1e :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h1f :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h20 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h21 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h22 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h23 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h24 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h25 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h26 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h27 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h28 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h29 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h2a :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h2b :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h2c :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h2d :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h2e :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h2f :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h30 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h31 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h32 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h33 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h34 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h35 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h36 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h37 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h38 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h39 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h3a :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h3b :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h3c :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h3d :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h3e :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h3f :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h40 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h41 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h42 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h43 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h44 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h45 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h46 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h47 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h48 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h49 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h4a :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h4b :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h4c :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h4d :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h4e :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h4f :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h50 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h51 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h52 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h53 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h54 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h55 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h56 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h57 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h58 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h59 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h5a :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h5b :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h5c :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h5d :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h5e :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h5f :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h60 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h61 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h62 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h63 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h64 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h65 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h66 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h67 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h68 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h69 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h6a :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h6b :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h6c :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h6d :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h6e :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h6f :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h70 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h71 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h72 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h73 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h74 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h75 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h76 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h77 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h78 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h79 :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h7a :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h7b :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h7c :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h7d :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h7e :
		TR_35 = RG_quantized_block_rl_9 ;
	7'h7f :
		TR_35 = RG_quantized_block_rl_9 ;
	default :
		TR_35 = 9'hx ;
	endcase
always @ ( RG_rl_141 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_36 = RG_rl_141 ;
	7'h01 :
		TR_36 = RG_rl_141 ;
	7'h02 :
		TR_36 = RG_rl_141 ;
	7'h03 :
		TR_36 = RG_rl_141 ;
	7'h04 :
		TR_36 = RG_rl_141 ;
	7'h05 :
		TR_36 = RG_rl_141 ;
	7'h06 :
		TR_36 = RG_rl_141 ;
	7'h07 :
		TR_36 = RG_rl_141 ;
	7'h08 :
		TR_36 = RG_rl_141 ;
	7'h09 :
		TR_36 = RG_rl_141 ;
	7'h0a :
		TR_36 = RG_rl_141 ;
	7'h0b :
		TR_36 = RG_rl_141 ;
	7'h0c :
		TR_36 = RG_rl_141 ;
	7'h0d :
		TR_36 = RG_rl_141 ;
	7'h0e :
		TR_36 = RG_rl_141 ;
	7'h0f :
		TR_36 = RG_rl_141 ;
	7'h10 :
		TR_36 = RG_rl_141 ;
	7'h11 :
		TR_36 = RG_rl_141 ;
	7'h12 :
		TR_36 = RG_rl_141 ;
	7'h13 :
		TR_36 = RG_rl_141 ;
	7'h14 :
		TR_36 = RG_rl_141 ;
	7'h15 :
		TR_36 = RG_rl_141 ;
	7'h16 :
		TR_36 = RG_rl_141 ;
	7'h17 :
		TR_36 = RG_rl_141 ;
	7'h18 :
		TR_36 = 9'h000 ;	// line#=../rle.cpp:79
	7'h19 :
		TR_36 = RG_rl_141 ;
	7'h1a :
		TR_36 = RG_rl_141 ;
	7'h1b :
		TR_36 = RG_rl_141 ;
	7'h1c :
		TR_36 = RG_rl_141 ;
	7'h1d :
		TR_36 = RG_rl_141 ;
	7'h1e :
		TR_36 = RG_rl_141 ;
	7'h1f :
		TR_36 = RG_rl_141 ;
	7'h20 :
		TR_36 = RG_rl_141 ;
	7'h21 :
		TR_36 = RG_rl_141 ;
	7'h22 :
		TR_36 = RG_rl_141 ;
	7'h23 :
		TR_36 = RG_rl_141 ;
	7'h24 :
		TR_36 = RG_rl_141 ;
	7'h25 :
		TR_36 = RG_rl_141 ;
	7'h26 :
		TR_36 = RG_rl_141 ;
	7'h27 :
		TR_36 = RG_rl_141 ;
	7'h28 :
		TR_36 = RG_rl_141 ;
	7'h29 :
		TR_36 = RG_rl_141 ;
	7'h2a :
		TR_36 = RG_rl_141 ;
	7'h2b :
		TR_36 = RG_rl_141 ;
	7'h2c :
		TR_36 = RG_rl_141 ;
	7'h2d :
		TR_36 = RG_rl_141 ;
	7'h2e :
		TR_36 = RG_rl_141 ;
	7'h2f :
		TR_36 = RG_rl_141 ;
	7'h30 :
		TR_36 = RG_rl_141 ;
	7'h31 :
		TR_36 = RG_rl_141 ;
	7'h32 :
		TR_36 = RG_rl_141 ;
	7'h33 :
		TR_36 = RG_rl_141 ;
	7'h34 :
		TR_36 = RG_rl_141 ;
	7'h35 :
		TR_36 = RG_rl_141 ;
	7'h36 :
		TR_36 = RG_rl_141 ;
	7'h37 :
		TR_36 = RG_rl_141 ;
	7'h38 :
		TR_36 = RG_rl_141 ;
	7'h39 :
		TR_36 = RG_rl_141 ;
	7'h3a :
		TR_36 = RG_rl_141 ;
	7'h3b :
		TR_36 = RG_rl_141 ;
	7'h3c :
		TR_36 = RG_rl_141 ;
	7'h3d :
		TR_36 = RG_rl_141 ;
	7'h3e :
		TR_36 = RG_rl_141 ;
	7'h3f :
		TR_36 = RG_rl_141 ;
	7'h40 :
		TR_36 = RG_rl_141 ;
	7'h41 :
		TR_36 = RG_rl_141 ;
	7'h42 :
		TR_36 = RG_rl_141 ;
	7'h43 :
		TR_36 = RG_rl_141 ;
	7'h44 :
		TR_36 = RG_rl_141 ;
	7'h45 :
		TR_36 = RG_rl_141 ;
	7'h46 :
		TR_36 = RG_rl_141 ;
	7'h47 :
		TR_36 = RG_rl_141 ;
	7'h48 :
		TR_36 = RG_rl_141 ;
	7'h49 :
		TR_36 = RG_rl_141 ;
	7'h4a :
		TR_36 = RG_rl_141 ;
	7'h4b :
		TR_36 = RG_rl_141 ;
	7'h4c :
		TR_36 = RG_rl_141 ;
	7'h4d :
		TR_36 = RG_rl_141 ;
	7'h4e :
		TR_36 = RG_rl_141 ;
	7'h4f :
		TR_36 = RG_rl_141 ;
	7'h50 :
		TR_36 = RG_rl_141 ;
	7'h51 :
		TR_36 = RG_rl_141 ;
	7'h52 :
		TR_36 = RG_rl_141 ;
	7'h53 :
		TR_36 = RG_rl_141 ;
	7'h54 :
		TR_36 = RG_rl_141 ;
	7'h55 :
		TR_36 = RG_rl_141 ;
	7'h56 :
		TR_36 = RG_rl_141 ;
	7'h57 :
		TR_36 = RG_rl_141 ;
	7'h58 :
		TR_36 = RG_rl_141 ;
	7'h59 :
		TR_36 = RG_rl_141 ;
	7'h5a :
		TR_36 = RG_rl_141 ;
	7'h5b :
		TR_36 = RG_rl_141 ;
	7'h5c :
		TR_36 = RG_rl_141 ;
	7'h5d :
		TR_36 = RG_rl_141 ;
	7'h5e :
		TR_36 = RG_rl_141 ;
	7'h5f :
		TR_36 = RG_rl_141 ;
	7'h60 :
		TR_36 = RG_rl_141 ;
	7'h61 :
		TR_36 = RG_rl_141 ;
	7'h62 :
		TR_36 = RG_rl_141 ;
	7'h63 :
		TR_36 = RG_rl_141 ;
	7'h64 :
		TR_36 = RG_rl_141 ;
	7'h65 :
		TR_36 = RG_rl_141 ;
	7'h66 :
		TR_36 = RG_rl_141 ;
	7'h67 :
		TR_36 = RG_rl_141 ;
	7'h68 :
		TR_36 = RG_rl_141 ;
	7'h69 :
		TR_36 = RG_rl_141 ;
	7'h6a :
		TR_36 = RG_rl_141 ;
	7'h6b :
		TR_36 = RG_rl_141 ;
	7'h6c :
		TR_36 = RG_rl_141 ;
	7'h6d :
		TR_36 = RG_rl_141 ;
	7'h6e :
		TR_36 = RG_rl_141 ;
	7'h6f :
		TR_36 = RG_rl_141 ;
	7'h70 :
		TR_36 = RG_rl_141 ;
	7'h71 :
		TR_36 = RG_rl_141 ;
	7'h72 :
		TR_36 = RG_rl_141 ;
	7'h73 :
		TR_36 = RG_rl_141 ;
	7'h74 :
		TR_36 = RG_rl_141 ;
	7'h75 :
		TR_36 = RG_rl_141 ;
	7'h76 :
		TR_36 = RG_rl_141 ;
	7'h77 :
		TR_36 = RG_rl_141 ;
	7'h78 :
		TR_36 = RG_rl_141 ;
	7'h79 :
		TR_36 = RG_rl_141 ;
	7'h7a :
		TR_36 = RG_rl_141 ;
	7'h7b :
		TR_36 = RG_rl_141 ;
	7'h7c :
		TR_36 = RG_rl_141 ;
	7'h7d :
		TR_36 = RG_rl_141 ;
	7'h7e :
		TR_36 = RG_rl_141 ;
	7'h7f :
		TR_36 = RG_rl_141 ;
	default :
		TR_36 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_10 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h01 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h02 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h03 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h04 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h05 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h06 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h07 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h08 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h09 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h0a :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h0b :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h0c :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h0d :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h0e :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h0f :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h10 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h11 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h12 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h13 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h14 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h15 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h16 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h17 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h18 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h19 :
		TR_37 = 9'h000 ;	// line#=../rle.cpp:79
	7'h1a :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h1b :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h1c :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h1d :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h1e :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h1f :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h20 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h21 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h22 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h23 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h24 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h25 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h26 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h27 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h28 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h29 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h2a :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h2b :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h2c :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h2d :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h2e :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h2f :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h30 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h31 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h32 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h33 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h34 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h35 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h36 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h37 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h38 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h39 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h3a :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h3b :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h3c :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h3d :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h3e :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h3f :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h40 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h41 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h42 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h43 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h44 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h45 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h46 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h47 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h48 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h49 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h4a :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h4b :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h4c :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h4d :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h4e :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h4f :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h50 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h51 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h52 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h53 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h54 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h55 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h56 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h57 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h58 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h59 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h5a :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h5b :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h5c :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h5d :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h5e :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h5f :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h60 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h61 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h62 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h63 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h64 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h65 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h66 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h67 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h68 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h69 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h6a :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h6b :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h6c :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h6d :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h6e :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h6f :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h70 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h71 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h72 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h73 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h74 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h75 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h76 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h77 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h78 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h79 :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h7a :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h7b :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h7c :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h7d :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h7e :
		TR_37 = RG_quantized_block_rl_10 ;
	7'h7f :
		TR_37 = RG_quantized_block_rl_10 ;
	default :
		TR_37 = 9'hx ;
	endcase
always @ ( RG_rl_142 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_38 = RG_rl_142 ;
	7'h01 :
		TR_38 = RG_rl_142 ;
	7'h02 :
		TR_38 = RG_rl_142 ;
	7'h03 :
		TR_38 = RG_rl_142 ;
	7'h04 :
		TR_38 = RG_rl_142 ;
	7'h05 :
		TR_38 = RG_rl_142 ;
	7'h06 :
		TR_38 = RG_rl_142 ;
	7'h07 :
		TR_38 = RG_rl_142 ;
	7'h08 :
		TR_38 = RG_rl_142 ;
	7'h09 :
		TR_38 = RG_rl_142 ;
	7'h0a :
		TR_38 = RG_rl_142 ;
	7'h0b :
		TR_38 = RG_rl_142 ;
	7'h0c :
		TR_38 = RG_rl_142 ;
	7'h0d :
		TR_38 = RG_rl_142 ;
	7'h0e :
		TR_38 = RG_rl_142 ;
	7'h0f :
		TR_38 = RG_rl_142 ;
	7'h10 :
		TR_38 = RG_rl_142 ;
	7'h11 :
		TR_38 = RG_rl_142 ;
	7'h12 :
		TR_38 = RG_rl_142 ;
	7'h13 :
		TR_38 = RG_rl_142 ;
	7'h14 :
		TR_38 = RG_rl_142 ;
	7'h15 :
		TR_38 = RG_rl_142 ;
	7'h16 :
		TR_38 = RG_rl_142 ;
	7'h17 :
		TR_38 = RG_rl_142 ;
	7'h18 :
		TR_38 = RG_rl_142 ;
	7'h19 :
		TR_38 = RG_rl_142 ;
	7'h1a :
		TR_38 = 9'h000 ;	// line#=../rle.cpp:79
	7'h1b :
		TR_38 = RG_rl_142 ;
	7'h1c :
		TR_38 = RG_rl_142 ;
	7'h1d :
		TR_38 = RG_rl_142 ;
	7'h1e :
		TR_38 = RG_rl_142 ;
	7'h1f :
		TR_38 = RG_rl_142 ;
	7'h20 :
		TR_38 = RG_rl_142 ;
	7'h21 :
		TR_38 = RG_rl_142 ;
	7'h22 :
		TR_38 = RG_rl_142 ;
	7'h23 :
		TR_38 = RG_rl_142 ;
	7'h24 :
		TR_38 = RG_rl_142 ;
	7'h25 :
		TR_38 = RG_rl_142 ;
	7'h26 :
		TR_38 = RG_rl_142 ;
	7'h27 :
		TR_38 = RG_rl_142 ;
	7'h28 :
		TR_38 = RG_rl_142 ;
	7'h29 :
		TR_38 = RG_rl_142 ;
	7'h2a :
		TR_38 = RG_rl_142 ;
	7'h2b :
		TR_38 = RG_rl_142 ;
	7'h2c :
		TR_38 = RG_rl_142 ;
	7'h2d :
		TR_38 = RG_rl_142 ;
	7'h2e :
		TR_38 = RG_rl_142 ;
	7'h2f :
		TR_38 = RG_rl_142 ;
	7'h30 :
		TR_38 = RG_rl_142 ;
	7'h31 :
		TR_38 = RG_rl_142 ;
	7'h32 :
		TR_38 = RG_rl_142 ;
	7'h33 :
		TR_38 = RG_rl_142 ;
	7'h34 :
		TR_38 = RG_rl_142 ;
	7'h35 :
		TR_38 = RG_rl_142 ;
	7'h36 :
		TR_38 = RG_rl_142 ;
	7'h37 :
		TR_38 = RG_rl_142 ;
	7'h38 :
		TR_38 = RG_rl_142 ;
	7'h39 :
		TR_38 = RG_rl_142 ;
	7'h3a :
		TR_38 = RG_rl_142 ;
	7'h3b :
		TR_38 = RG_rl_142 ;
	7'h3c :
		TR_38 = RG_rl_142 ;
	7'h3d :
		TR_38 = RG_rl_142 ;
	7'h3e :
		TR_38 = RG_rl_142 ;
	7'h3f :
		TR_38 = RG_rl_142 ;
	7'h40 :
		TR_38 = RG_rl_142 ;
	7'h41 :
		TR_38 = RG_rl_142 ;
	7'h42 :
		TR_38 = RG_rl_142 ;
	7'h43 :
		TR_38 = RG_rl_142 ;
	7'h44 :
		TR_38 = RG_rl_142 ;
	7'h45 :
		TR_38 = RG_rl_142 ;
	7'h46 :
		TR_38 = RG_rl_142 ;
	7'h47 :
		TR_38 = RG_rl_142 ;
	7'h48 :
		TR_38 = RG_rl_142 ;
	7'h49 :
		TR_38 = RG_rl_142 ;
	7'h4a :
		TR_38 = RG_rl_142 ;
	7'h4b :
		TR_38 = RG_rl_142 ;
	7'h4c :
		TR_38 = RG_rl_142 ;
	7'h4d :
		TR_38 = RG_rl_142 ;
	7'h4e :
		TR_38 = RG_rl_142 ;
	7'h4f :
		TR_38 = RG_rl_142 ;
	7'h50 :
		TR_38 = RG_rl_142 ;
	7'h51 :
		TR_38 = RG_rl_142 ;
	7'h52 :
		TR_38 = RG_rl_142 ;
	7'h53 :
		TR_38 = RG_rl_142 ;
	7'h54 :
		TR_38 = RG_rl_142 ;
	7'h55 :
		TR_38 = RG_rl_142 ;
	7'h56 :
		TR_38 = RG_rl_142 ;
	7'h57 :
		TR_38 = RG_rl_142 ;
	7'h58 :
		TR_38 = RG_rl_142 ;
	7'h59 :
		TR_38 = RG_rl_142 ;
	7'h5a :
		TR_38 = RG_rl_142 ;
	7'h5b :
		TR_38 = RG_rl_142 ;
	7'h5c :
		TR_38 = RG_rl_142 ;
	7'h5d :
		TR_38 = RG_rl_142 ;
	7'h5e :
		TR_38 = RG_rl_142 ;
	7'h5f :
		TR_38 = RG_rl_142 ;
	7'h60 :
		TR_38 = RG_rl_142 ;
	7'h61 :
		TR_38 = RG_rl_142 ;
	7'h62 :
		TR_38 = RG_rl_142 ;
	7'h63 :
		TR_38 = RG_rl_142 ;
	7'h64 :
		TR_38 = RG_rl_142 ;
	7'h65 :
		TR_38 = RG_rl_142 ;
	7'h66 :
		TR_38 = RG_rl_142 ;
	7'h67 :
		TR_38 = RG_rl_142 ;
	7'h68 :
		TR_38 = RG_rl_142 ;
	7'h69 :
		TR_38 = RG_rl_142 ;
	7'h6a :
		TR_38 = RG_rl_142 ;
	7'h6b :
		TR_38 = RG_rl_142 ;
	7'h6c :
		TR_38 = RG_rl_142 ;
	7'h6d :
		TR_38 = RG_rl_142 ;
	7'h6e :
		TR_38 = RG_rl_142 ;
	7'h6f :
		TR_38 = RG_rl_142 ;
	7'h70 :
		TR_38 = RG_rl_142 ;
	7'h71 :
		TR_38 = RG_rl_142 ;
	7'h72 :
		TR_38 = RG_rl_142 ;
	7'h73 :
		TR_38 = RG_rl_142 ;
	7'h74 :
		TR_38 = RG_rl_142 ;
	7'h75 :
		TR_38 = RG_rl_142 ;
	7'h76 :
		TR_38 = RG_rl_142 ;
	7'h77 :
		TR_38 = RG_rl_142 ;
	7'h78 :
		TR_38 = RG_rl_142 ;
	7'h79 :
		TR_38 = RG_rl_142 ;
	7'h7a :
		TR_38 = RG_rl_142 ;
	7'h7b :
		TR_38 = RG_rl_142 ;
	7'h7c :
		TR_38 = RG_rl_142 ;
	7'h7d :
		TR_38 = RG_rl_142 ;
	7'h7e :
		TR_38 = RG_rl_142 ;
	7'h7f :
		TR_38 = RG_rl_142 ;
	default :
		TR_38 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_11 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h01 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h02 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h03 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h04 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h05 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h06 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h07 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h08 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h09 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h0a :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h0b :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h0c :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h0d :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h0e :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h0f :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h10 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h11 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h12 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h13 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h14 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h15 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h16 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h17 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h18 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h19 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h1a :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h1b :
		TR_39 = 9'h000 ;	// line#=../rle.cpp:79
	7'h1c :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h1d :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h1e :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h1f :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h20 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h21 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h22 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h23 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h24 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h25 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h26 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h27 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h28 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h29 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h2a :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h2b :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h2c :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h2d :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h2e :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h2f :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h30 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h31 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h32 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h33 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h34 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h35 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h36 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h37 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h38 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h39 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h3a :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h3b :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h3c :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h3d :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h3e :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h3f :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h40 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h41 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h42 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h43 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h44 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h45 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h46 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h47 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h48 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h49 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h4a :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h4b :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h4c :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h4d :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h4e :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h4f :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h50 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h51 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h52 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h53 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h54 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h55 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h56 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h57 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h58 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h59 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h5a :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h5b :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h5c :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h5d :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h5e :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h5f :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h60 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h61 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h62 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h63 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h64 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h65 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h66 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h67 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h68 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h69 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h6a :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h6b :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h6c :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h6d :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h6e :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h6f :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h70 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h71 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h72 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h73 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h74 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h75 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h76 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h77 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h78 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h79 :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h7a :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h7b :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h7c :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h7d :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h7e :
		TR_39 = RG_quantized_block_rl_11 ;
	7'h7f :
		TR_39 = RG_quantized_block_rl_11 ;
	default :
		TR_39 = 9'hx ;
	endcase
always @ ( RG_rl_143 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_40 = RG_rl_143 ;
	7'h01 :
		TR_40 = RG_rl_143 ;
	7'h02 :
		TR_40 = RG_rl_143 ;
	7'h03 :
		TR_40 = RG_rl_143 ;
	7'h04 :
		TR_40 = RG_rl_143 ;
	7'h05 :
		TR_40 = RG_rl_143 ;
	7'h06 :
		TR_40 = RG_rl_143 ;
	7'h07 :
		TR_40 = RG_rl_143 ;
	7'h08 :
		TR_40 = RG_rl_143 ;
	7'h09 :
		TR_40 = RG_rl_143 ;
	7'h0a :
		TR_40 = RG_rl_143 ;
	7'h0b :
		TR_40 = RG_rl_143 ;
	7'h0c :
		TR_40 = RG_rl_143 ;
	7'h0d :
		TR_40 = RG_rl_143 ;
	7'h0e :
		TR_40 = RG_rl_143 ;
	7'h0f :
		TR_40 = RG_rl_143 ;
	7'h10 :
		TR_40 = RG_rl_143 ;
	7'h11 :
		TR_40 = RG_rl_143 ;
	7'h12 :
		TR_40 = RG_rl_143 ;
	7'h13 :
		TR_40 = RG_rl_143 ;
	7'h14 :
		TR_40 = RG_rl_143 ;
	7'h15 :
		TR_40 = RG_rl_143 ;
	7'h16 :
		TR_40 = RG_rl_143 ;
	7'h17 :
		TR_40 = RG_rl_143 ;
	7'h18 :
		TR_40 = RG_rl_143 ;
	7'h19 :
		TR_40 = RG_rl_143 ;
	7'h1a :
		TR_40 = RG_rl_143 ;
	7'h1b :
		TR_40 = RG_rl_143 ;
	7'h1c :
		TR_40 = 9'h000 ;	// line#=../rle.cpp:79
	7'h1d :
		TR_40 = RG_rl_143 ;
	7'h1e :
		TR_40 = RG_rl_143 ;
	7'h1f :
		TR_40 = RG_rl_143 ;
	7'h20 :
		TR_40 = RG_rl_143 ;
	7'h21 :
		TR_40 = RG_rl_143 ;
	7'h22 :
		TR_40 = RG_rl_143 ;
	7'h23 :
		TR_40 = RG_rl_143 ;
	7'h24 :
		TR_40 = RG_rl_143 ;
	7'h25 :
		TR_40 = RG_rl_143 ;
	7'h26 :
		TR_40 = RG_rl_143 ;
	7'h27 :
		TR_40 = RG_rl_143 ;
	7'h28 :
		TR_40 = RG_rl_143 ;
	7'h29 :
		TR_40 = RG_rl_143 ;
	7'h2a :
		TR_40 = RG_rl_143 ;
	7'h2b :
		TR_40 = RG_rl_143 ;
	7'h2c :
		TR_40 = RG_rl_143 ;
	7'h2d :
		TR_40 = RG_rl_143 ;
	7'h2e :
		TR_40 = RG_rl_143 ;
	7'h2f :
		TR_40 = RG_rl_143 ;
	7'h30 :
		TR_40 = RG_rl_143 ;
	7'h31 :
		TR_40 = RG_rl_143 ;
	7'h32 :
		TR_40 = RG_rl_143 ;
	7'h33 :
		TR_40 = RG_rl_143 ;
	7'h34 :
		TR_40 = RG_rl_143 ;
	7'h35 :
		TR_40 = RG_rl_143 ;
	7'h36 :
		TR_40 = RG_rl_143 ;
	7'h37 :
		TR_40 = RG_rl_143 ;
	7'h38 :
		TR_40 = RG_rl_143 ;
	7'h39 :
		TR_40 = RG_rl_143 ;
	7'h3a :
		TR_40 = RG_rl_143 ;
	7'h3b :
		TR_40 = RG_rl_143 ;
	7'h3c :
		TR_40 = RG_rl_143 ;
	7'h3d :
		TR_40 = RG_rl_143 ;
	7'h3e :
		TR_40 = RG_rl_143 ;
	7'h3f :
		TR_40 = RG_rl_143 ;
	7'h40 :
		TR_40 = RG_rl_143 ;
	7'h41 :
		TR_40 = RG_rl_143 ;
	7'h42 :
		TR_40 = RG_rl_143 ;
	7'h43 :
		TR_40 = RG_rl_143 ;
	7'h44 :
		TR_40 = RG_rl_143 ;
	7'h45 :
		TR_40 = RG_rl_143 ;
	7'h46 :
		TR_40 = RG_rl_143 ;
	7'h47 :
		TR_40 = RG_rl_143 ;
	7'h48 :
		TR_40 = RG_rl_143 ;
	7'h49 :
		TR_40 = RG_rl_143 ;
	7'h4a :
		TR_40 = RG_rl_143 ;
	7'h4b :
		TR_40 = RG_rl_143 ;
	7'h4c :
		TR_40 = RG_rl_143 ;
	7'h4d :
		TR_40 = RG_rl_143 ;
	7'h4e :
		TR_40 = RG_rl_143 ;
	7'h4f :
		TR_40 = RG_rl_143 ;
	7'h50 :
		TR_40 = RG_rl_143 ;
	7'h51 :
		TR_40 = RG_rl_143 ;
	7'h52 :
		TR_40 = RG_rl_143 ;
	7'h53 :
		TR_40 = RG_rl_143 ;
	7'h54 :
		TR_40 = RG_rl_143 ;
	7'h55 :
		TR_40 = RG_rl_143 ;
	7'h56 :
		TR_40 = RG_rl_143 ;
	7'h57 :
		TR_40 = RG_rl_143 ;
	7'h58 :
		TR_40 = RG_rl_143 ;
	7'h59 :
		TR_40 = RG_rl_143 ;
	7'h5a :
		TR_40 = RG_rl_143 ;
	7'h5b :
		TR_40 = RG_rl_143 ;
	7'h5c :
		TR_40 = RG_rl_143 ;
	7'h5d :
		TR_40 = RG_rl_143 ;
	7'h5e :
		TR_40 = RG_rl_143 ;
	7'h5f :
		TR_40 = RG_rl_143 ;
	7'h60 :
		TR_40 = RG_rl_143 ;
	7'h61 :
		TR_40 = RG_rl_143 ;
	7'h62 :
		TR_40 = RG_rl_143 ;
	7'h63 :
		TR_40 = RG_rl_143 ;
	7'h64 :
		TR_40 = RG_rl_143 ;
	7'h65 :
		TR_40 = RG_rl_143 ;
	7'h66 :
		TR_40 = RG_rl_143 ;
	7'h67 :
		TR_40 = RG_rl_143 ;
	7'h68 :
		TR_40 = RG_rl_143 ;
	7'h69 :
		TR_40 = RG_rl_143 ;
	7'h6a :
		TR_40 = RG_rl_143 ;
	7'h6b :
		TR_40 = RG_rl_143 ;
	7'h6c :
		TR_40 = RG_rl_143 ;
	7'h6d :
		TR_40 = RG_rl_143 ;
	7'h6e :
		TR_40 = RG_rl_143 ;
	7'h6f :
		TR_40 = RG_rl_143 ;
	7'h70 :
		TR_40 = RG_rl_143 ;
	7'h71 :
		TR_40 = RG_rl_143 ;
	7'h72 :
		TR_40 = RG_rl_143 ;
	7'h73 :
		TR_40 = RG_rl_143 ;
	7'h74 :
		TR_40 = RG_rl_143 ;
	7'h75 :
		TR_40 = RG_rl_143 ;
	7'h76 :
		TR_40 = RG_rl_143 ;
	7'h77 :
		TR_40 = RG_rl_143 ;
	7'h78 :
		TR_40 = RG_rl_143 ;
	7'h79 :
		TR_40 = RG_rl_143 ;
	7'h7a :
		TR_40 = RG_rl_143 ;
	7'h7b :
		TR_40 = RG_rl_143 ;
	7'h7c :
		TR_40 = RG_rl_143 ;
	7'h7d :
		TR_40 = RG_rl_143 ;
	7'h7e :
		TR_40 = RG_rl_143 ;
	7'h7f :
		TR_40 = RG_rl_143 ;
	default :
		TR_40 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_12 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h01 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h02 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h03 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h04 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h05 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h06 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h07 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h08 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h09 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h0a :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h0b :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h0c :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h0d :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h0e :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h0f :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h10 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h11 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h12 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h13 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h14 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h15 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h16 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h17 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h18 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h19 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h1a :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h1b :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h1c :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h1d :
		TR_41 = 9'h000 ;	// line#=../rle.cpp:79
	7'h1e :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h1f :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h20 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h21 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h22 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h23 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h24 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h25 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h26 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h27 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h28 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h29 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h2a :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h2b :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h2c :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h2d :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h2e :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h2f :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h30 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h31 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h32 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h33 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h34 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h35 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h36 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h37 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h38 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h39 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h3a :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h3b :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h3c :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h3d :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h3e :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h3f :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h40 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h41 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h42 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h43 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h44 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h45 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h46 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h47 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h48 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h49 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h4a :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h4b :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h4c :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h4d :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h4e :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h4f :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h50 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h51 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h52 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h53 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h54 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h55 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h56 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h57 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h58 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h59 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h5a :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h5b :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h5c :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h5d :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h5e :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h5f :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h60 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h61 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h62 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h63 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h64 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h65 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h66 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h67 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h68 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h69 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h6a :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h6b :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h6c :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h6d :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h6e :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h6f :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h70 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h71 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h72 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h73 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h74 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h75 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h76 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h77 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h78 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h79 :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h7a :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h7b :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h7c :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h7d :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h7e :
		TR_41 = RG_quantized_block_rl_12 ;
	7'h7f :
		TR_41 = RG_quantized_block_rl_12 ;
	default :
		TR_41 = 9'hx ;
	endcase
always @ ( RG_rl_144 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_42 = RG_rl_144 ;
	7'h01 :
		TR_42 = RG_rl_144 ;
	7'h02 :
		TR_42 = RG_rl_144 ;
	7'h03 :
		TR_42 = RG_rl_144 ;
	7'h04 :
		TR_42 = RG_rl_144 ;
	7'h05 :
		TR_42 = RG_rl_144 ;
	7'h06 :
		TR_42 = RG_rl_144 ;
	7'h07 :
		TR_42 = RG_rl_144 ;
	7'h08 :
		TR_42 = RG_rl_144 ;
	7'h09 :
		TR_42 = RG_rl_144 ;
	7'h0a :
		TR_42 = RG_rl_144 ;
	7'h0b :
		TR_42 = RG_rl_144 ;
	7'h0c :
		TR_42 = RG_rl_144 ;
	7'h0d :
		TR_42 = RG_rl_144 ;
	7'h0e :
		TR_42 = RG_rl_144 ;
	7'h0f :
		TR_42 = RG_rl_144 ;
	7'h10 :
		TR_42 = RG_rl_144 ;
	7'h11 :
		TR_42 = RG_rl_144 ;
	7'h12 :
		TR_42 = RG_rl_144 ;
	7'h13 :
		TR_42 = RG_rl_144 ;
	7'h14 :
		TR_42 = RG_rl_144 ;
	7'h15 :
		TR_42 = RG_rl_144 ;
	7'h16 :
		TR_42 = RG_rl_144 ;
	7'h17 :
		TR_42 = RG_rl_144 ;
	7'h18 :
		TR_42 = RG_rl_144 ;
	7'h19 :
		TR_42 = RG_rl_144 ;
	7'h1a :
		TR_42 = RG_rl_144 ;
	7'h1b :
		TR_42 = RG_rl_144 ;
	7'h1c :
		TR_42 = RG_rl_144 ;
	7'h1d :
		TR_42 = RG_rl_144 ;
	7'h1e :
		TR_42 = 9'h000 ;	// line#=../rle.cpp:79
	7'h1f :
		TR_42 = RG_rl_144 ;
	7'h20 :
		TR_42 = RG_rl_144 ;
	7'h21 :
		TR_42 = RG_rl_144 ;
	7'h22 :
		TR_42 = RG_rl_144 ;
	7'h23 :
		TR_42 = RG_rl_144 ;
	7'h24 :
		TR_42 = RG_rl_144 ;
	7'h25 :
		TR_42 = RG_rl_144 ;
	7'h26 :
		TR_42 = RG_rl_144 ;
	7'h27 :
		TR_42 = RG_rl_144 ;
	7'h28 :
		TR_42 = RG_rl_144 ;
	7'h29 :
		TR_42 = RG_rl_144 ;
	7'h2a :
		TR_42 = RG_rl_144 ;
	7'h2b :
		TR_42 = RG_rl_144 ;
	7'h2c :
		TR_42 = RG_rl_144 ;
	7'h2d :
		TR_42 = RG_rl_144 ;
	7'h2e :
		TR_42 = RG_rl_144 ;
	7'h2f :
		TR_42 = RG_rl_144 ;
	7'h30 :
		TR_42 = RG_rl_144 ;
	7'h31 :
		TR_42 = RG_rl_144 ;
	7'h32 :
		TR_42 = RG_rl_144 ;
	7'h33 :
		TR_42 = RG_rl_144 ;
	7'h34 :
		TR_42 = RG_rl_144 ;
	7'h35 :
		TR_42 = RG_rl_144 ;
	7'h36 :
		TR_42 = RG_rl_144 ;
	7'h37 :
		TR_42 = RG_rl_144 ;
	7'h38 :
		TR_42 = RG_rl_144 ;
	7'h39 :
		TR_42 = RG_rl_144 ;
	7'h3a :
		TR_42 = RG_rl_144 ;
	7'h3b :
		TR_42 = RG_rl_144 ;
	7'h3c :
		TR_42 = RG_rl_144 ;
	7'h3d :
		TR_42 = RG_rl_144 ;
	7'h3e :
		TR_42 = RG_rl_144 ;
	7'h3f :
		TR_42 = RG_rl_144 ;
	7'h40 :
		TR_42 = RG_rl_144 ;
	7'h41 :
		TR_42 = RG_rl_144 ;
	7'h42 :
		TR_42 = RG_rl_144 ;
	7'h43 :
		TR_42 = RG_rl_144 ;
	7'h44 :
		TR_42 = RG_rl_144 ;
	7'h45 :
		TR_42 = RG_rl_144 ;
	7'h46 :
		TR_42 = RG_rl_144 ;
	7'h47 :
		TR_42 = RG_rl_144 ;
	7'h48 :
		TR_42 = RG_rl_144 ;
	7'h49 :
		TR_42 = RG_rl_144 ;
	7'h4a :
		TR_42 = RG_rl_144 ;
	7'h4b :
		TR_42 = RG_rl_144 ;
	7'h4c :
		TR_42 = RG_rl_144 ;
	7'h4d :
		TR_42 = RG_rl_144 ;
	7'h4e :
		TR_42 = RG_rl_144 ;
	7'h4f :
		TR_42 = RG_rl_144 ;
	7'h50 :
		TR_42 = RG_rl_144 ;
	7'h51 :
		TR_42 = RG_rl_144 ;
	7'h52 :
		TR_42 = RG_rl_144 ;
	7'h53 :
		TR_42 = RG_rl_144 ;
	7'h54 :
		TR_42 = RG_rl_144 ;
	7'h55 :
		TR_42 = RG_rl_144 ;
	7'h56 :
		TR_42 = RG_rl_144 ;
	7'h57 :
		TR_42 = RG_rl_144 ;
	7'h58 :
		TR_42 = RG_rl_144 ;
	7'h59 :
		TR_42 = RG_rl_144 ;
	7'h5a :
		TR_42 = RG_rl_144 ;
	7'h5b :
		TR_42 = RG_rl_144 ;
	7'h5c :
		TR_42 = RG_rl_144 ;
	7'h5d :
		TR_42 = RG_rl_144 ;
	7'h5e :
		TR_42 = RG_rl_144 ;
	7'h5f :
		TR_42 = RG_rl_144 ;
	7'h60 :
		TR_42 = RG_rl_144 ;
	7'h61 :
		TR_42 = RG_rl_144 ;
	7'h62 :
		TR_42 = RG_rl_144 ;
	7'h63 :
		TR_42 = RG_rl_144 ;
	7'h64 :
		TR_42 = RG_rl_144 ;
	7'h65 :
		TR_42 = RG_rl_144 ;
	7'h66 :
		TR_42 = RG_rl_144 ;
	7'h67 :
		TR_42 = RG_rl_144 ;
	7'h68 :
		TR_42 = RG_rl_144 ;
	7'h69 :
		TR_42 = RG_rl_144 ;
	7'h6a :
		TR_42 = RG_rl_144 ;
	7'h6b :
		TR_42 = RG_rl_144 ;
	7'h6c :
		TR_42 = RG_rl_144 ;
	7'h6d :
		TR_42 = RG_rl_144 ;
	7'h6e :
		TR_42 = RG_rl_144 ;
	7'h6f :
		TR_42 = RG_rl_144 ;
	7'h70 :
		TR_42 = RG_rl_144 ;
	7'h71 :
		TR_42 = RG_rl_144 ;
	7'h72 :
		TR_42 = RG_rl_144 ;
	7'h73 :
		TR_42 = RG_rl_144 ;
	7'h74 :
		TR_42 = RG_rl_144 ;
	7'h75 :
		TR_42 = RG_rl_144 ;
	7'h76 :
		TR_42 = RG_rl_144 ;
	7'h77 :
		TR_42 = RG_rl_144 ;
	7'h78 :
		TR_42 = RG_rl_144 ;
	7'h79 :
		TR_42 = RG_rl_144 ;
	7'h7a :
		TR_42 = RG_rl_144 ;
	7'h7b :
		TR_42 = RG_rl_144 ;
	7'h7c :
		TR_42 = RG_rl_144 ;
	7'h7d :
		TR_42 = RG_rl_144 ;
	7'h7e :
		TR_42 = RG_rl_144 ;
	7'h7f :
		TR_42 = RG_rl_144 ;
	default :
		TR_42 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_13 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h01 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h02 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h03 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h04 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h05 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h06 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h07 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h08 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h09 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h0a :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h0b :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h0c :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h0d :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h0e :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h0f :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h10 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h11 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h12 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h13 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h14 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h15 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h16 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h17 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h18 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h19 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h1a :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h1b :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h1c :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h1d :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h1e :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h1f :
		TR_43 = 9'h000 ;	// line#=../rle.cpp:79
	7'h20 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h21 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h22 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h23 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h24 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h25 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h26 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h27 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h28 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h29 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h2a :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h2b :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h2c :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h2d :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h2e :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h2f :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h30 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h31 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h32 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h33 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h34 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h35 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h36 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h37 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h38 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h39 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h3a :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h3b :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h3c :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h3d :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h3e :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h3f :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h40 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h41 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h42 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h43 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h44 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h45 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h46 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h47 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h48 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h49 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h4a :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h4b :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h4c :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h4d :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h4e :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h4f :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h50 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h51 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h52 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h53 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h54 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h55 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h56 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h57 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h58 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h59 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h5a :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h5b :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h5c :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h5d :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h5e :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h5f :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h60 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h61 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h62 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h63 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h64 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h65 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h66 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h67 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h68 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h69 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h6a :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h6b :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h6c :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h6d :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h6e :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h6f :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h70 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h71 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h72 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h73 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h74 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h75 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h76 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h77 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h78 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h79 :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h7a :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h7b :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h7c :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h7d :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h7e :
		TR_43 = RG_quantized_block_rl_13 ;
	7'h7f :
		TR_43 = RG_quantized_block_rl_13 ;
	default :
		TR_43 = 9'hx ;
	endcase
always @ ( RG_rl_145 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_44 = RG_rl_145 ;
	7'h01 :
		TR_44 = RG_rl_145 ;
	7'h02 :
		TR_44 = RG_rl_145 ;
	7'h03 :
		TR_44 = RG_rl_145 ;
	7'h04 :
		TR_44 = RG_rl_145 ;
	7'h05 :
		TR_44 = RG_rl_145 ;
	7'h06 :
		TR_44 = RG_rl_145 ;
	7'h07 :
		TR_44 = RG_rl_145 ;
	7'h08 :
		TR_44 = RG_rl_145 ;
	7'h09 :
		TR_44 = RG_rl_145 ;
	7'h0a :
		TR_44 = RG_rl_145 ;
	7'h0b :
		TR_44 = RG_rl_145 ;
	7'h0c :
		TR_44 = RG_rl_145 ;
	7'h0d :
		TR_44 = RG_rl_145 ;
	7'h0e :
		TR_44 = RG_rl_145 ;
	7'h0f :
		TR_44 = RG_rl_145 ;
	7'h10 :
		TR_44 = RG_rl_145 ;
	7'h11 :
		TR_44 = RG_rl_145 ;
	7'h12 :
		TR_44 = RG_rl_145 ;
	7'h13 :
		TR_44 = RG_rl_145 ;
	7'h14 :
		TR_44 = RG_rl_145 ;
	7'h15 :
		TR_44 = RG_rl_145 ;
	7'h16 :
		TR_44 = RG_rl_145 ;
	7'h17 :
		TR_44 = RG_rl_145 ;
	7'h18 :
		TR_44 = RG_rl_145 ;
	7'h19 :
		TR_44 = RG_rl_145 ;
	7'h1a :
		TR_44 = RG_rl_145 ;
	7'h1b :
		TR_44 = RG_rl_145 ;
	7'h1c :
		TR_44 = RG_rl_145 ;
	7'h1d :
		TR_44 = RG_rl_145 ;
	7'h1e :
		TR_44 = RG_rl_145 ;
	7'h1f :
		TR_44 = RG_rl_145 ;
	7'h20 :
		TR_44 = 9'h000 ;	// line#=../rle.cpp:79
	7'h21 :
		TR_44 = RG_rl_145 ;
	7'h22 :
		TR_44 = RG_rl_145 ;
	7'h23 :
		TR_44 = RG_rl_145 ;
	7'h24 :
		TR_44 = RG_rl_145 ;
	7'h25 :
		TR_44 = RG_rl_145 ;
	7'h26 :
		TR_44 = RG_rl_145 ;
	7'h27 :
		TR_44 = RG_rl_145 ;
	7'h28 :
		TR_44 = RG_rl_145 ;
	7'h29 :
		TR_44 = RG_rl_145 ;
	7'h2a :
		TR_44 = RG_rl_145 ;
	7'h2b :
		TR_44 = RG_rl_145 ;
	7'h2c :
		TR_44 = RG_rl_145 ;
	7'h2d :
		TR_44 = RG_rl_145 ;
	7'h2e :
		TR_44 = RG_rl_145 ;
	7'h2f :
		TR_44 = RG_rl_145 ;
	7'h30 :
		TR_44 = RG_rl_145 ;
	7'h31 :
		TR_44 = RG_rl_145 ;
	7'h32 :
		TR_44 = RG_rl_145 ;
	7'h33 :
		TR_44 = RG_rl_145 ;
	7'h34 :
		TR_44 = RG_rl_145 ;
	7'h35 :
		TR_44 = RG_rl_145 ;
	7'h36 :
		TR_44 = RG_rl_145 ;
	7'h37 :
		TR_44 = RG_rl_145 ;
	7'h38 :
		TR_44 = RG_rl_145 ;
	7'h39 :
		TR_44 = RG_rl_145 ;
	7'h3a :
		TR_44 = RG_rl_145 ;
	7'h3b :
		TR_44 = RG_rl_145 ;
	7'h3c :
		TR_44 = RG_rl_145 ;
	7'h3d :
		TR_44 = RG_rl_145 ;
	7'h3e :
		TR_44 = RG_rl_145 ;
	7'h3f :
		TR_44 = RG_rl_145 ;
	7'h40 :
		TR_44 = RG_rl_145 ;
	7'h41 :
		TR_44 = RG_rl_145 ;
	7'h42 :
		TR_44 = RG_rl_145 ;
	7'h43 :
		TR_44 = RG_rl_145 ;
	7'h44 :
		TR_44 = RG_rl_145 ;
	7'h45 :
		TR_44 = RG_rl_145 ;
	7'h46 :
		TR_44 = RG_rl_145 ;
	7'h47 :
		TR_44 = RG_rl_145 ;
	7'h48 :
		TR_44 = RG_rl_145 ;
	7'h49 :
		TR_44 = RG_rl_145 ;
	7'h4a :
		TR_44 = RG_rl_145 ;
	7'h4b :
		TR_44 = RG_rl_145 ;
	7'h4c :
		TR_44 = RG_rl_145 ;
	7'h4d :
		TR_44 = RG_rl_145 ;
	7'h4e :
		TR_44 = RG_rl_145 ;
	7'h4f :
		TR_44 = RG_rl_145 ;
	7'h50 :
		TR_44 = RG_rl_145 ;
	7'h51 :
		TR_44 = RG_rl_145 ;
	7'h52 :
		TR_44 = RG_rl_145 ;
	7'h53 :
		TR_44 = RG_rl_145 ;
	7'h54 :
		TR_44 = RG_rl_145 ;
	7'h55 :
		TR_44 = RG_rl_145 ;
	7'h56 :
		TR_44 = RG_rl_145 ;
	7'h57 :
		TR_44 = RG_rl_145 ;
	7'h58 :
		TR_44 = RG_rl_145 ;
	7'h59 :
		TR_44 = RG_rl_145 ;
	7'h5a :
		TR_44 = RG_rl_145 ;
	7'h5b :
		TR_44 = RG_rl_145 ;
	7'h5c :
		TR_44 = RG_rl_145 ;
	7'h5d :
		TR_44 = RG_rl_145 ;
	7'h5e :
		TR_44 = RG_rl_145 ;
	7'h5f :
		TR_44 = RG_rl_145 ;
	7'h60 :
		TR_44 = RG_rl_145 ;
	7'h61 :
		TR_44 = RG_rl_145 ;
	7'h62 :
		TR_44 = RG_rl_145 ;
	7'h63 :
		TR_44 = RG_rl_145 ;
	7'h64 :
		TR_44 = RG_rl_145 ;
	7'h65 :
		TR_44 = RG_rl_145 ;
	7'h66 :
		TR_44 = RG_rl_145 ;
	7'h67 :
		TR_44 = RG_rl_145 ;
	7'h68 :
		TR_44 = RG_rl_145 ;
	7'h69 :
		TR_44 = RG_rl_145 ;
	7'h6a :
		TR_44 = RG_rl_145 ;
	7'h6b :
		TR_44 = RG_rl_145 ;
	7'h6c :
		TR_44 = RG_rl_145 ;
	7'h6d :
		TR_44 = RG_rl_145 ;
	7'h6e :
		TR_44 = RG_rl_145 ;
	7'h6f :
		TR_44 = RG_rl_145 ;
	7'h70 :
		TR_44 = RG_rl_145 ;
	7'h71 :
		TR_44 = RG_rl_145 ;
	7'h72 :
		TR_44 = RG_rl_145 ;
	7'h73 :
		TR_44 = RG_rl_145 ;
	7'h74 :
		TR_44 = RG_rl_145 ;
	7'h75 :
		TR_44 = RG_rl_145 ;
	7'h76 :
		TR_44 = RG_rl_145 ;
	7'h77 :
		TR_44 = RG_rl_145 ;
	7'h78 :
		TR_44 = RG_rl_145 ;
	7'h79 :
		TR_44 = RG_rl_145 ;
	7'h7a :
		TR_44 = RG_rl_145 ;
	7'h7b :
		TR_44 = RG_rl_145 ;
	7'h7c :
		TR_44 = RG_rl_145 ;
	7'h7d :
		TR_44 = RG_rl_145 ;
	7'h7e :
		TR_44 = RG_rl_145 ;
	7'h7f :
		TR_44 = RG_rl_145 ;
	default :
		TR_44 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_14 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h01 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h02 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h03 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h04 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h05 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h06 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h07 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h08 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h09 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h0a :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h0b :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h0c :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h0d :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h0e :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h0f :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h10 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h11 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h12 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h13 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h14 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h15 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h16 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h17 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h18 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h19 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h1a :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h1b :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h1c :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h1d :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h1e :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h1f :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h20 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h21 :
		TR_45 = 9'h000 ;	// line#=../rle.cpp:79
	7'h22 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h23 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h24 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h25 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h26 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h27 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h28 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h29 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h2a :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h2b :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h2c :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h2d :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h2e :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h2f :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h30 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h31 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h32 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h33 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h34 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h35 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h36 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h37 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h38 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h39 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h3a :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h3b :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h3c :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h3d :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h3e :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h3f :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h40 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h41 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h42 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h43 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h44 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h45 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h46 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h47 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h48 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h49 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h4a :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h4b :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h4c :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h4d :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h4e :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h4f :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h50 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h51 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h52 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h53 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h54 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h55 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h56 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h57 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h58 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h59 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h5a :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h5b :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h5c :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h5d :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h5e :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h5f :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h60 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h61 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h62 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h63 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h64 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h65 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h66 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h67 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h68 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h69 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h6a :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h6b :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h6c :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h6d :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h6e :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h6f :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h70 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h71 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h72 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h73 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h74 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h75 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h76 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h77 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h78 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h79 :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h7a :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h7b :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h7c :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h7d :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h7e :
		TR_45 = RG_quantized_block_rl_14 ;
	7'h7f :
		TR_45 = RG_quantized_block_rl_14 ;
	default :
		TR_45 = 9'hx ;
	endcase
always @ ( RG_rl_146 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_46 = RG_rl_146 ;
	7'h01 :
		TR_46 = RG_rl_146 ;
	7'h02 :
		TR_46 = RG_rl_146 ;
	7'h03 :
		TR_46 = RG_rl_146 ;
	7'h04 :
		TR_46 = RG_rl_146 ;
	7'h05 :
		TR_46 = RG_rl_146 ;
	7'h06 :
		TR_46 = RG_rl_146 ;
	7'h07 :
		TR_46 = RG_rl_146 ;
	7'h08 :
		TR_46 = RG_rl_146 ;
	7'h09 :
		TR_46 = RG_rl_146 ;
	7'h0a :
		TR_46 = RG_rl_146 ;
	7'h0b :
		TR_46 = RG_rl_146 ;
	7'h0c :
		TR_46 = RG_rl_146 ;
	7'h0d :
		TR_46 = RG_rl_146 ;
	7'h0e :
		TR_46 = RG_rl_146 ;
	7'h0f :
		TR_46 = RG_rl_146 ;
	7'h10 :
		TR_46 = RG_rl_146 ;
	7'h11 :
		TR_46 = RG_rl_146 ;
	7'h12 :
		TR_46 = RG_rl_146 ;
	7'h13 :
		TR_46 = RG_rl_146 ;
	7'h14 :
		TR_46 = RG_rl_146 ;
	7'h15 :
		TR_46 = RG_rl_146 ;
	7'h16 :
		TR_46 = RG_rl_146 ;
	7'h17 :
		TR_46 = RG_rl_146 ;
	7'h18 :
		TR_46 = RG_rl_146 ;
	7'h19 :
		TR_46 = RG_rl_146 ;
	7'h1a :
		TR_46 = RG_rl_146 ;
	7'h1b :
		TR_46 = RG_rl_146 ;
	7'h1c :
		TR_46 = RG_rl_146 ;
	7'h1d :
		TR_46 = RG_rl_146 ;
	7'h1e :
		TR_46 = RG_rl_146 ;
	7'h1f :
		TR_46 = RG_rl_146 ;
	7'h20 :
		TR_46 = RG_rl_146 ;
	7'h21 :
		TR_46 = RG_rl_146 ;
	7'h22 :
		TR_46 = 9'h000 ;	// line#=../rle.cpp:79
	7'h23 :
		TR_46 = RG_rl_146 ;
	7'h24 :
		TR_46 = RG_rl_146 ;
	7'h25 :
		TR_46 = RG_rl_146 ;
	7'h26 :
		TR_46 = RG_rl_146 ;
	7'h27 :
		TR_46 = RG_rl_146 ;
	7'h28 :
		TR_46 = RG_rl_146 ;
	7'h29 :
		TR_46 = RG_rl_146 ;
	7'h2a :
		TR_46 = RG_rl_146 ;
	7'h2b :
		TR_46 = RG_rl_146 ;
	7'h2c :
		TR_46 = RG_rl_146 ;
	7'h2d :
		TR_46 = RG_rl_146 ;
	7'h2e :
		TR_46 = RG_rl_146 ;
	7'h2f :
		TR_46 = RG_rl_146 ;
	7'h30 :
		TR_46 = RG_rl_146 ;
	7'h31 :
		TR_46 = RG_rl_146 ;
	7'h32 :
		TR_46 = RG_rl_146 ;
	7'h33 :
		TR_46 = RG_rl_146 ;
	7'h34 :
		TR_46 = RG_rl_146 ;
	7'h35 :
		TR_46 = RG_rl_146 ;
	7'h36 :
		TR_46 = RG_rl_146 ;
	7'h37 :
		TR_46 = RG_rl_146 ;
	7'h38 :
		TR_46 = RG_rl_146 ;
	7'h39 :
		TR_46 = RG_rl_146 ;
	7'h3a :
		TR_46 = RG_rl_146 ;
	7'h3b :
		TR_46 = RG_rl_146 ;
	7'h3c :
		TR_46 = RG_rl_146 ;
	7'h3d :
		TR_46 = RG_rl_146 ;
	7'h3e :
		TR_46 = RG_rl_146 ;
	7'h3f :
		TR_46 = RG_rl_146 ;
	7'h40 :
		TR_46 = RG_rl_146 ;
	7'h41 :
		TR_46 = RG_rl_146 ;
	7'h42 :
		TR_46 = RG_rl_146 ;
	7'h43 :
		TR_46 = RG_rl_146 ;
	7'h44 :
		TR_46 = RG_rl_146 ;
	7'h45 :
		TR_46 = RG_rl_146 ;
	7'h46 :
		TR_46 = RG_rl_146 ;
	7'h47 :
		TR_46 = RG_rl_146 ;
	7'h48 :
		TR_46 = RG_rl_146 ;
	7'h49 :
		TR_46 = RG_rl_146 ;
	7'h4a :
		TR_46 = RG_rl_146 ;
	7'h4b :
		TR_46 = RG_rl_146 ;
	7'h4c :
		TR_46 = RG_rl_146 ;
	7'h4d :
		TR_46 = RG_rl_146 ;
	7'h4e :
		TR_46 = RG_rl_146 ;
	7'h4f :
		TR_46 = RG_rl_146 ;
	7'h50 :
		TR_46 = RG_rl_146 ;
	7'h51 :
		TR_46 = RG_rl_146 ;
	7'h52 :
		TR_46 = RG_rl_146 ;
	7'h53 :
		TR_46 = RG_rl_146 ;
	7'h54 :
		TR_46 = RG_rl_146 ;
	7'h55 :
		TR_46 = RG_rl_146 ;
	7'h56 :
		TR_46 = RG_rl_146 ;
	7'h57 :
		TR_46 = RG_rl_146 ;
	7'h58 :
		TR_46 = RG_rl_146 ;
	7'h59 :
		TR_46 = RG_rl_146 ;
	7'h5a :
		TR_46 = RG_rl_146 ;
	7'h5b :
		TR_46 = RG_rl_146 ;
	7'h5c :
		TR_46 = RG_rl_146 ;
	7'h5d :
		TR_46 = RG_rl_146 ;
	7'h5e :
		TR_46 = RG_rl_146 ;
	7'h5f :
		TR_46 = RG_rl_146 ;
	7'h60 :
		TR_46 = RG_rl_146 ;
	7'h61 :
		TR_46 = RG_rl_146 ;
	7'h62 :
		TR_46 = RG_rl_146 ;
	7'h63 :
		TR_46 = RG_rl_146 ;
	7'h64 :
		TR_46 = RG_rl_146 ;
	7'h65 :
		TR_46 = RG_rl_146 ;
	7'h66 :
		TR_46 = RG_rl_146 ;
	7'h67 :
		TR_46 = RG_rl_146 ;
	7'h68 :
		TR_46 = RG_rl_146 ;
	7'h69 :
		TR_46 = RG_rl_146 ;
	7'h6a :
		TR_46 = RG_rl_146 ;
	7'h6b :
		TR_46 = RG_rl_146 ;
	7'h6c :
		TR_46 = RG_rl_146 ;
	7'h6d :
		TR_46 = RG_rl_146 ;
	7'h6e :
		TR_46 = RG_rl_146 ;
	7'h6f :
		TR_46 = RG_rl_146 ;
	7'h70 :
		TR_46 = RG_rl_146 ;
	7'h71 :
		TR_46 = RG_rl_146 ;
	7'h72 :
		TR_46 = RG_rl_146 ;
	7'h73 :
		TR_46 = RG_rl_146 ;
	7'h74 :
		TR_46 = RG_rl_146 ;
	7'h75 :
		TR_46 = RG_rl_146 ;
	7'h76 :
		TR_46 = RG_rl_146 ;
	7'h77 :
		TR_46 = RG_rl_146 ;
	7'h78 :
		TR_46 = RG_rl_146 ;
	7'h79 :
		TR_46 = RG_rl_146 ;
	7'h7a :
		TR_46 = RG_rl_146 ;
	7'h7b :
		TR_46 = RG_rl_146 ;
	7'h7c :
		TR_46 = RG_rl_146 ;
	7'h7d :
		TR_46 = RG_rl_146 ;
	7'h7e :
		TR_46 = RG_rl_146 ;
	7'h7f :
		TR_46 = RG_rl_146 ;
	default :
		TR_46 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_15 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h01 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h02 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h03 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h04 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h05 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h06 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h07 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h08 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h09 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h0a :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h0b :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h0c :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h0d :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h0e :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h0f :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h10 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h11 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h12 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h13 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h14 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h15 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h16 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h17 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h18 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h19 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h1a :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h1b :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h1c :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h1d :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h1e :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h1f :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h20 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h21 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h22 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h23 :
		TR_47 = 9'h000 ;	// line#=../rle.cpp:79
	7'h24 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h25 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h26 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h27 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h28 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h29 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h2a :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h2b :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h2c :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h2d :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h2e :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h2f :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h30 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h31 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h32 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h33 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h34 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h35 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h36 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h37 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h38 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h39 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h3a :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h3b :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h3c :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h3d :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h3e :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h3f :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h40 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h41 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h42 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h43 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h44 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h45 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h46 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h47 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h48 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h49 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h4a :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h4b :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h4c :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h4d :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h4e :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h4f :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h50 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h51 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h52 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h53 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h54 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h55 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h56 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h57 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h58 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h59 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h5a :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h5b :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h5c :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h5d :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h5e :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h5f :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h60 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h61 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h62 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h63 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h64 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h65 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h66 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h67 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h68 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h69 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h6a :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h6b :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h6c :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h6d :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h6e :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h6f :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h70 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h71 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h72 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h73 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h74 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h75 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h76 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h77 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h78 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h79 :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h7a :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h7b :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h7c :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h7d :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h7e :
		TR_47 = RG_quantized_block_rl_15 ;
	7'h7f :
		TR_47 = RG_quantized_block_rl_15 ;
	default :
		TR_47 = 9'hx ;
	endcase
always @ ( RG_rl_147 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_48 = RG_rl_147 ;
	7'h01 :
		TR_48 = RG_rl_147 ;
	7'h02 :
		TR_48 = RG_rl_147 ;
	7'h03 :
		TR_48 = RG_rl_147 ;
	7'h04 :
		TR_48 = RG_rl_147 ;
	7'h05 :
		TR_48 = RG_rl_147 ;
	7'h06 :
		TR_48 = RG_rl_147 ;
	7'h07 :
		TR_48 = RG_rl_147 ;
	7'h08 :
		TR_48 = RG_rl_147 ;
	7'h09 :
		TR_48 = RG_rl_147 ;
	7'h0a :
		TR_48 = RG_rl_147 ;
	7'h0b :
		TR_48 = RG_rl_147 ;
	7'h0c :
		TR_48 = RG_rl_147 ;
	7'h0d :
		TR_48 = RG_rl_147 ;
	7'h0e :
		TR_48 = RG_rl_147 ;
	7'h0f :
		TR_48 = RG_rl_147 ;
	7'h10 :
		TR_48 = RG_rl_147 ;
	7'h11 :
		TR_48 = RG_rl_147 ;
	7'h12 :
		TR_48 = RG_rl_147 ;
	7'h13 :
		TR_48 = RG_rl_147 ;
	7'h14 :
		TR_48 = RG_rl_147 ;
	7'h15 :
		TR_48 = RG_rl_147 ;
	7'h16 :
		TR_48 = RG_rl_147 ;
	7'h17 :
		TR_48 = RG_rl_147 ;
	7'h18 :
		TR_48 = RG_rl_147 ;
	7'h19 :
		TR_48 = RG_rl_147 ;
	7'h1a :
		TR_48 = RG_rl_147 ;
	7'h1b :
		TR_48 = RG_rl_147 ;
	7'h1c :
		TR_48 = RG_rl_147 ;
	7'h1d :
		TR_48 = RG_rl_147 ;
	7'h1e :
		TR_48 = RG_rl_147 ;
	7'h1f :
		TR_48 = RG_rl_147 ;
	7'h20 :
		TR_48 = RG_rl_147 ;
	7'h21 :
		TR_48 = RG_rl_147 ;
	7'h22 :
		TR_48 = RG_rl_147 ;
	7'h23 :
		TR_48 = RG_rl_147 ;
	7'h24 :
		TR_48 = 9'h000 ;	// line#=../rle.cpp:79
	7'h25 :
		TR_48 = RG_rl_147 ;
	7'h26 :
		TR_48 = RG_rl_147 ;
	7'h27 :
		TR_48 = RG_rl_147 ;
	7'h28 :
		TR_48 = RG_rl_147 ;
	7'h29 :
		TR_48 = RG_rl_147 ;
	7'h2a :
		TR_48 = RG_rl_147 ;
	7'h2b :
		TR_48 = RG_rl_147 ;
	7'h2c :
		TR_48 = RG_rl_147 ;
	7'h2d :
		TR_48 = RG_rl_147 ;
	7'h2e :
		TR_48 = RG_rl_147 ;
	7'h2f :
		TR_48 = RG_rl_147 ;
	7'h30 :
		TR_48 = RG_rl_147 ;
	7'h31 :
		TR_48 = RG_rl_147 ;
	7'h32 :
		TR_48 = RG_rl_147 ;
	7'h33 :
		TR_48 = RG_rl_147 ;
	7'h34 :
		TR_48 = RG_rl_147 ;
	7'h35 :
		TR_48 = RG_rl_147 ;
	7'h36 :
		TR_48 = RG_rl_147 ;
	7'h37 :
		TR_48 = RG_rl_147 ;
	7'h38 :
		TR_48 = RG_rl_147 ;
	7'h39 :
		TR_48 = RG_rl_147 ;
	7'h3a :
		TR_48 = RG_rl_147 ;
	7'h3b :
		TR_48 = RG_rl_147 ;
	7'h3c :
		TR_48 = RG_rl_147 ;
	7'h3d :
		TR_48 = RG_rl_147 ;
	7'h3e :
		TR_48 = RG_rl_147 ;
	7'h3f :
		TR_48 = RG_rl_147 ;
	7'h40 :
		TR_48 = RG_rl_147 ;
	7'h41 :
		TR_48 = RG_rl_147 ;
	7'h42 :
		TR_48 = RG_rl_147 ;
	7'h43 :
		TR_48 = RG_rl_147 ;
	7'h44 :
		TR_48 = RG_rl_147 ;
	7'h45 :
		TR_48 = RG_rl_147 ;
	7'h46 :
		TR_48 = RG_rl_147 ;
	7'h47 :
		TR_48 = RG_rl_147 ;
	7'h48 :
		TR_48 = RG_rl_147 ;
	7'h49 :
		TR_48 = RG_rl_147 ;
	7'h4a :
		TR_48 = RG_rl_147 ;
	7'h4b :
		TR_48 = RG_rl_147 ;
	7'h4c :
		TR_48 = RG_rl_147 ;
	7'h4d :
		TR_48 = RG_rl_147 ;
	7'h4e :
		TR_48 = RG_rl_147 ;
	7'h4f :
		TR_48 = RG_rl_147 ;
	7'h50 :
		TR_48 = RG_rl_147 ;
	7'h51 :
		TR_48 = RG_rl_147 ;
	7'h52 :
		TR_48 = RG_rl_147 ;
	7'h53 :
		TR_48 = RG_rl_147 ;
	7'h54 :
		TR_48 = RG_rl_147 ;
	7'h55 :
		TR_48 = RG_rl_147 ;
	7'h56 :
		TR_48 = RG_rl_147 ;
	7'h57 :
		TR_48 = RG_rl_147 ;
	7'h58 :
		TR_48 = RG_rl_147 ;
	7'h59 :
		TR_48 = RG_rl_147 ;
	7'h5a :
		TR_48 = RG_rl_147 ;
	7'h5b :
		TR_48 = RG_rl_147 ;
	7'h5c :
		TR_48 = RG_rl_147 ;
	7'h5d :
		TR_48 = RG_rl_147 ;
	7'h5e :
		TR_48 = RG_rl_147 ;
	7'h5f :
		TR_48 = RG_rl_147 ;
	7'h60 :
		TR_48 = RG_rl_147 ;
	7'h61 :
		TR_48 = RG_rl_147 ;
	7'h62 :
		TR_48 = RG_rl_147 ;
	7'h63 :
		TR_48 = RG_rl_147 ;
	7'h64 :
		TR_48 = RG_rl_147 ;
	7'h65 :
		TR_48 = RG_rl_147 ;
	7'h66 :
		TR_48 = RG_rl_147 ;
	7'h67 :
		TR_48 = RG_rl_147 ;
	7'h68 :
		TR_48 = RG_rl_147 ;
	7'h69 :
		TR_48 = RG_rl_147 ;
	7'h6a :
		TR_48 = RG_rl_147 ;
	7'h6b :
		TR_48 = RG_rl_147 ;
	7'h6c :
		TR_48 = RG_rl_147 ;
	7'h6d :
		TR_48 = RG_rl_147 ;
	7'h6e :
		TR_48 = RG_rl_147 ;
	7'h6f :
		TR_48 = RG_rl_147 ;
	7'h70 :
		TR_48 = RG_rl_147 ;
	7'h71 :
		TR_48 = RG_rl_147 ;
	7'h72 :
		TR_48 = RG_rl_147 ;
	7'h73 :
		TR_48 = RG_rl_147 ;
	7'h74 :
		TR_48 = RG_rl_147 ;
	7'h75 :
		TR_48 = RG_rl_147 ;
	7'h76 :
		TR_48 = RG_rl_147 ;
	7'h77 :
		TR_48 = RG_rl_147 ;
	7'h78 :
		TR_48 = RG_rl_147 ;
	7'h79 :
		TR_48 = RG_rl_147 ;
	7'h7a :
		TR_48 = RG_rl_147 ;
	7'h7b :
		TR_48 = RG_rl_147 ;
	7'h7c :
		TR_48 = RG_rl_147 ;
	7'h7d :
		TR_48 = RG_rl_147 ;
	7'h7e :
		TR_48 = RG_rl_147 ;
	7'h7f :
		TR_48 = RG_rl_147 ;
	default :
		TR_48 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_16 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h01 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h02 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h03 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h04 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h05 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h06 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h07 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h08 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h09 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h0a :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h0b :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h0c :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h0d :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h0e :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h0f :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h10 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h11 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h12 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h13 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h14 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h15 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h16 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h17 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h18 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h19 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h1a :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h1b :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h1c :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h1d :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h1e :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h1f :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h20 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h21 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h22 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h23 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h24 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h25 :
		TR_49 = 9'h000 ;	// line#=../rle.cpp:79
	7'h26 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h27 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h28 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h29 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h2a :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h2b :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h2c :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h2d :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h2e :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h2f :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h30 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h31 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h32 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h33 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h34 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h35 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h36 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h37 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h38 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h39 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h3a :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h3b :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h3c :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h3d :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h3e :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h3f :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h40 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h41 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h42 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h43 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h44 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h45 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h46 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h47 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h48 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h49 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h4a :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h4b :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h4c :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h4d :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h4e :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h4f :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h50 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h51 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h52 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h53 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h54 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h55 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h56 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h57 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h58 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h59 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h5a :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h5b :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h5c :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h5d :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h5e :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h5f :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h60 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h61 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h62 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h63 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h64 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h65 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h66 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h67 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h68 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h69 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h6a :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h6b :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h6c :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h6d :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h6e :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h6f :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h70 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h71 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h72 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h73 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h74 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h75 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h76 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h77 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h78 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h79 :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h7a :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h7b :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h7c :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h7d :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h7e :
		TR_49 = RG_quantized_block_rl_16 ;
	7'h7f :
		TR_49 = RG_quantized_block_rl_16 ;
	default :
		TR_49 = 9'hx ;
	endcase
always @ ( RG_rl_148 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_50 = RG_rl_148 ;
	7'h01 :
		TR_50 = RG_rl_148 ;
	7'h02 :
		TR_50 = RG_rl_148 ;
	7'h03 :
		TR_50 = RG_rl_148 ;
	7'h04 :
		TR_50 = RG_rl_148 ;
	7'h05 :
		TR_50 = RG_rl_148 ;
	7'h06 :
		TR_50 = RG_rl_148 ;
	7'h07 :
		TR_50 = RG_rl_148 ;
	7'h08 :
		TR_50 = RG_rl_148 ;
	7'h09 :
		TR_50 = RG_rl_148 ;
	7'h0a :
		TR_50 = RG_rl_148 ;
	7'h0b :
		TR_50 = RG_rl_148 ;
	7'h0c :
		TR_50 = RG_rl_148 ;
	7'h0d :
		TR_50 = RG_rl_148 ;
	7'h0e :
		TR_50 = RG_rl_148 ;
	7'h0f :
		TR_50 = RG_rl_148 ;
	7'h10 :
		TR_50 = RG_rl_148 ;
	7'h11 :
		TR_50 = RG_rl_148 ;
	7'h12 :
		TR_50 = RG_rl_148 ;
	7'h13 :
		TR_50 = RG_rl_148 ;
	7'h14 :
		TR_50 = RG_rl_148 ;
	7'h15 :
		TR_50 = RG_rl_148 ;
	7'h16 :
		TR_50 = RG_rl_148 ;
	7'h17 :
		TR_50 = RG_rl_148 ;
	7'h18 :
		TR_50 = RG_rl_148 ;
	7'h19 :
		TR_50 = RG_rl_148 ;
	7'h1a :
		TR_50 = RG_rl_148 ;
	7'h1b :
		TR_50 = RG_rl_148 ;
	7'h1c :
		TR_50 = RG_rl_148 ;
	7'h1d :
		TR_50 = RG_rl_148 ;
	7'h1e :
		TR_50 = RG_rl_148 ;
	7'h1f :
		TR_50 = RG_rl_148 ;
	7'h20 :
		TR_50 = RG_rl_148 ;
	7'h21 :
		TR_50 = RG_rl_148 ;
	7'h22 :
		TR_50 = RG_rl_148 ;
	7'h23 :
		TR_50 = RG_rl_148 ;
	7'h24 :
		TR_50 = RG_rl_148 ;
	7'h25 :
		TR_50 = RG_rl_148 ;
	7'h26 :
		TR_50 = 9'h000 ;	// line#=../rle.cpp:79
	7'h27 :
		TR_50 = RG_rl_148 ;
	7'h28 :
		TR_50 = RG_rl_148 ;
	7'h29 :
		TR_50 = RG_rl_148 ;
	7'h2a :
		TR_50 = RG_rl_148 ;
	7'h2b :
		TR_50 = RG_rl_148 ;
	7'h2c :
		TR_50 = RG_rl_148 ;
	7'h2d :
		TR_50 = RG_rl_148 ;
	7'h2e :
		TR_50 = RG_rl_148 ;
	7'h2f :
		TR_50 = RG_rl_148 ;
	7'h30 :
		TR_50 = RG_rl_148 ;
	7'h31 :
		TR_50 = RG_rl_148 ;
	7'h32 :
		TR_50 = RG_rl_148 ;
	7'h33 :
		TR_50 = RG_rl_148 ;
	7'h34 :
		TR_50 = RG_rl_148 ;
	7'h35 :
		TR_50 = RG_rl_148 ;
	7'h36 :
		TR_50 = RG_rl_148 ;
	7'h37 :
		TR_50 = RG_rl_148 ;
	7'h38 :
		TR_50 = RG_rl_148 ;
	7'h39 :
		TR_50 = RG_rl_148 ;
	7'h3a :
		TR_50 = RG_rl_148 ;
	7'h3b :
		TR_50 = RG_rl_148 ;
	7'h3c :
		TR_50 = RG_rl_148 ;
	7'h3d :
		TR_50 = RG_rl_148 ;
	7'h3e :
		TR_50 = RG_rl_148 ;
	7'h3f :
		TR_50 = RG_rl_148 ;
	7'h40 :
		TR_50 = RG_rl_148 ;
	7'h41 :
		TR_50 = RG_rl_148 ;
	7'h42 :
		TR_50 = RG_rl_148 ;
	7'h43 :
		TR_50 = RG_rl_148 ;
	7'h44 :
		TR_50 = RG_rl_148 ;
	7'h45 :
		TR_50 = RG_rl_148 ;
	7'h46 :
		TR_50 = RG_rl_148 ;
	7'h47 :
		TR_50 = RG_rl_148 ;
	7'h48 :
		TR_50 = RG_rl_148 ;
	7'h49 :
		TR_50 = RG_rl_148 ;
	7'h4a :
		TR_50 = RG_rl_148 ;
	7'h4b :
		TR_50 = RG_rl_148 ;
	7'h4c :
		TR_50 = RG_rl_148 ;
	7'h4d :
		TR_50 = RG_rl_148 ;
	7'h4e :
		TR_50 = RG_rl_148 ;
	7'h4f :
		TR_50 = RG_rl_148 ;
	7'h50 :
		TR_50 = RG_rl_148 ;
	7'h51 :
		TR_50 = RG_rl_148 ;
	7'h52 :
		TR_50 = RG_rl_148 ;
	7'h53 :
		TR_50 = RG_rl_148 ;
	7'h54 :
		TR_50 = RG_rl_148 ;
	7'h55 :
		TR_50 = RG_rl_148 ;
	7'h56 :
		TR_50 = RG_rl_148 ;
	7'h57 :
		TR_50 = RG_rl_148 ;
	7'h58 :
		TR_50 = RG_rl_148 ;
	7'h59 :
		TR_50 = RG_rl_148 ;
	7'h5a :
		TR_50 = RG_rl_148 ;
	7'h5b :
		TR_50 = RG_rl_148 ;
	7'h5c :
		TR_50 = RG_rl_148 ;
	7'h5d :
		TR_50 = RG_rl_148 ;
	7'h5e :
		TR_50 = RG_rl_148 ;
	7'h5f :
		TR_50 = RG_rl_148 ;
	7'h60 :
		TR_50 = RG_rl_148 ;
	7'h61 :
		TR_50 = RG_rl_148 ;
	7'h62 :
		TR_50 = RG_rl_148 ;
	7'h63 :
		TR_50 = RG_rl_148 ;
	7'h64 :
		TR_50 = RG_rl_148 ;
	7'h65 :
		TR_50 = RG_rl_148 ;
	7'h66 :
		TR_50 = RG_rl_148 ;
	7'h67 :
		TR_50 = RG_rl_148 ;
	7'h68 :
		TR_50 = RG_rl_148 ;
	7'h69 :
		TR_50 = RG_rl_148 ;
	7'h6a :
		TR_50 = RG_rl_148 ;
	7'h6b :
		TR_50 = RG_rl_148 ;
	7'h6c :
		TR_50 = RG_rl_148 ;
	7'h6d :
		TR_50 = RG_rl_148 ;
	7'h6e :
		TR_50 = RG_rl_148 ;
	7'h6f :
		TR_50 = RG_rl_148 ;
	7'h70 :
		TR_50 = RG_rl_148 ;
	7'h71 :
		TR_50 = RG_rl_148 ;
	7'h72 :
		TR_50 = RG_rl_148 ;
	7'h73 :
		TR_50 = RG_rl_148 ;
	7'h74 :
		TR_50 = RG_rl_148 ;
	7'h75 :
		TR_50 = RG_rl_148 ;
	7'h76 :
		TR_50 = RG_rl_148 ;
	7'h77 :
		TR_50 = RG_rl_148 ;
	7'h78 :
		TR_50 = RG_rl_148 ;
	7'h79 :
		TR_50 = RG_rl_148 ;
	7'h7a :
		TR_50 = RG_rl_148 ;
	7'h7b :
		TR_50 = RG_rl_148 ;
	7'h7c :
		TR_50 = RG_rl_148 ;
	7'h7d :
		TR_50 = RG_rl_148 ;
	7'h7e :
		TR_50 = RG_rl_148 ;
	7'h7f :
		TR_50 = RG_rl_148 ;
	default :
		TR_50 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_17 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h01 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h02 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h03 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h04 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h05 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h06 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h07 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h08 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h09 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h0a :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h0b :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h0c :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h0d :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h0e :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h0f :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h10 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h11 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h12 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h13 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h14 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h15 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h16 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h17 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h18 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h19 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h1a :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h1b :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h1c :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h1d :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h1e :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h1f :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h20 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h21 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h22 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h23 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h24 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h25 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h26 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h27 :
		TR_51 = 9'h000 ;	// line#=../rle.cpp:79
	7'h28 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h29 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h2a :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h2b :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h2c :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h2d :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h2e :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h2f :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h30 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h31 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h32 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h33 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h34 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h35 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h36 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h37 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h38 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h39 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h3a :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h3b :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h3c :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h3d :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h3e :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h3f :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h40 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h41 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h42 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h43 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h44 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h45 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h46 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h47 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h48 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h49 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h4a :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h4b :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h4c :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h4d :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h4e :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h4f :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h50 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h51 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h52 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h53 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h54 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h55 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h56 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h57 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h58 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h59 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h5a :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h5b :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h5c :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h5d :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h5e :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h5f :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h60 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h61 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h62 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h63 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h64 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h65 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h66 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h67 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h68 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h69 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h6a :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h6b :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h6c :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h6d :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h6e :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h6f :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h70 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h71 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h72 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h73 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h74 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h75 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h76 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h77 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h78 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h79 :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h7a :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h7b :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h7c :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h7d :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h7e :
		TR_51 = RG_quantized_block_rl_17 ;
	7'h7f :
		TR_51 = RG_quantized_block_rl_17 ;
	default :
		TR_51 = 9'hx ;
	endcase
always @ ( RG_rl_149 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_52 = RG_rl_149 ;
	7'h01 :
		TR_52 = RG_rl_149 ;
	7'h02 :
		TR_52 = RG_rl_149 ;
	7'h03 :
		TR_52 = RG_rl_149 ;
	7'h04 :
		TR_52 = RG_rl_149 ;
	7'h05 :
		TR_52 = RG_rl_149 ;
	7'h06 :
		TR_52 = RG_rl_149 ;
	7'h07 :
		TR_52 = RG_rl_149 ;
	7'h08 :
		TR_52 = RG_rl_149 ;
	7'h09 :
		TR_52 = RG_rl_149 ;
	7'h0a :
		TR_52 = RG_rl_149 ;
	7'h0b :
		TR_52 = RG_rl_149 ;
	7'h0c :
		TR_52 = RG_rl_149 ;
	7'h0d :
		TR_52 = RG_rl_149 ;
	7'h0e :
		TR_52 = RG_rl_149 ;
	7'h0f :
		TR_52 = RG_rl_149 ;
	7'h10 :
		TR_52 = RG_rl_149 ;
	7'h11 :
		TR_52 = RG_rl_149 ;
	7'h12 :
		TR_52 = RG_rl_149 ;
	7'h13 :
		TR_52 = RG_rl_149 ;
	7'h14 :
		TR_52 = RG_rl_149 ;
	7'h15 :
		TR_52 = RG_rl_149 ;
	7'h16 :
		TR_52 = RG_rl_149 ;
	7'h17 :
		TR_52 = RG_rl_149 ;
	7'h18 :
		TR_52 = RG_rl_149 ;
	7'h19 :
		TR_52 = RG_rl_149 ;
	7'h1a :
		TR_52 = RG_rl_149 ;
	7'h1b :
		TR_52 = RG_rl_149 ;
	7'h1c :
		TR_52 = RG_rl_149 ;
	7'h1d :
		TR_52 = RG_rl_149 ;
	7'h1e :
		TR_52 = RG_rl_149 ;
	7'h1f :
		TR_52 = RG_rl_149 ;
	7'h20 :
		TR_52 = RG_rl_149 ;
	7'h21 :
		TR_52 = RG_rl_149 ;
	7'h22 :
		TR_52 = RG_rl_149 ;
	7'h23 :
		TR_52 = RG_rl_149 ;
	7'h24 :
		TR_52 = RG_rl_149 ;
	7'h25 :
		TR_52 = RG_rl_149 ;
	7'h26 :
		TR_52 = RG_rl_149 ;
	7'h27 :
		TR_52 = RG_rl_149 ;
	7'h28 :
		TR_52 = 9'h000 ;	// line#=../rle.cpp:79
	7'h29 :
		TR_52 = RG_rl_149 ;
	7'h2a :
		TR_52 = RG_rl_149 ;
	7'h2b :
		TR_52 = RG_rl_149 ;
	7'h2c :
		TR_52 = RG_rl_149 ;
	7'h2d :
		TR_52 = RG_rl_149 ;
	7'h2e :
		TR_52 = RG_rl_149 ;
	7'h2f :
		TR_52 = RG_rl_149 ;
	7'h30 :
		TR_52 = RG_rl_149 ;
	7'h31 :
		TR_52 = RG_rl_149 ;
	7'h32 :
		TR_52 = RG_rl_149 ;
	7'h33 :
		TR_52 = RG_rl_149 ;
	7'h34 :
		TR_52 = RG_rl_149 ;
	7'h35 :
		TR_52 = RG_rl_149 ;
	7'h36 :
		TR_52 = RG_rl_149 ;
	7'h37 :
		TR_52 = RG_rl_149 ;
	7'h38 :
		TR_52 = RG_rl_149 ;
	7'h39 :
		TR_52 = RG_rl_149 ;
	7'h3a :
		TR_52 = RG_rl_149 ;
	7'h3b :
		TR_52 = RG_rl_149 ;
	7'h3c :
		TR_52 = RG_rl_149 ;
	7'h3d :
		TR_52 = RG_rl_149 ;
	7'h3e :
		TR_52 = RG_rl_149 ;
	7'h3f :
		TR_52 = RG_rl_149 ;
	7'h40 :
		TR_52 = RG_rl_149 ;
	7'h41 :
		TR_52 = RG_rl_149 ;
	7'h42 :
		TR_52 = RG_rl_149 ;
	7'h43 :
		TR_52 = RG_rl_149 ;
	7'h44 :
		TR_52 = RG_rl_149 ;
	7'h45 :
		TR_52 = RG_rl_149 ;
	7'h46 :
		TR_52 = RG_rl_149 ;
	7'h47 :
		TR_52 = RG_rl_149 ;
	7'h48 :
		TR_52 = RG_rl_149 ;
	7'h49 :
		TR_52 = RG_rl_149 ;
	7'h4a :
		TR_52 = RG_rl_149 ;
	7'h4b :
		TR_52 = RG_rl_149 ;
	7'h4c :
		TR_52 = RG_rl_149 ;
	7'h4d :
		TR_52 = RG_rl_149 ;
	7'h4e :
		TR_52 = RG_rl_149 ;
	7'h4f :
		TR_52 = RG_rl_149 ;
	7'h50 :
		TR_52 = RG_rl_149 ;
	7'h51 :
		TR_52 = RG_rl_149 ;
	7'h52 :
		TR_52 = RG_rl_149 ;
	7'h53 :
		TR_52 = RG_rl_149 ;
	7'h54 :
		TR_52 = RG_rl_149 ;
	7'h55 :
		TR_52 = RG_rl_149 ;
	7'h56 :
		TR_52 = RG_rl_149 ;
	7'h57 :
		TR_52 = RG_rl_149 ;
	7'h58 :
		TR_52 = RG_rl_149 ;
	7'h59 :
		TR_52 = RG_rl_149 ;
	7'h5a :
		TR_52 = RG_rl_149 ;
	7'h5b :
		TR_52 = RG_rl_149 ;
	7'h5c :
		TR_52 = RG_rl_149 ;
	7'h5d :
		TR_52 = RG_rl_149 ;
	7'h5e :
		TR_52 = RG_rl_149 ;
	7'h5f :
		TR_52 = RG_rl_149 ;
	7'h60 :
		TR_52 = RG_rl_149 ;
	7'h61 :
		TR_52 = RG_rl_149 ;
	7'h62 :
		TR_52 = RG_rl_149 ;
	7'h63 :
		TR_52 = RG_rl_149 ;
	7'h64 :
		TR_52 = RG_rl_149 ;
	7'h65 :
		TR_52 = RG_rl_149 ;
	7'h66 :
		TR_52 = RG_rl_149 ;
	7'h67 :
		TR_52 = RG_rl_149 ;
	7'h68 :
		TR_52 = RG_rl_149 ;
	7'h69 :
		TR_52 = RG_rl_149 ;
	7'h6a :
		TR_52 = RG_rl_149 ;
	7'h6b :
		TR_52 = RG_rl_149 ;
	7'h6c :
		TR_52 = RG_rl_149 ;
	7'h6d :
		TR_52 = RG_rl_149 ;
	7'h6e :
		TR_52 = RG_rl_149 ;
	7'h6f :
		TR_52 = RG_rl_149 ;
	7'h70 :
		TR_52 = RG_rl_149 ;
	7'h71 :
		TR_52 = RG_rl_149 ;
	7'h72 :
		TR_52 = RG_rl_149 ;
	7'h73 :
		TR_52 = RG_rl_149 ;
	7'h74 :
		TR_52 = RG_rl_149 ;
	7'h75 :
		TR_52 = RG_rl_149 ;
	7'h76 :
		TR_52 = RG_rl_149 ;
	7'h77 :
		TR_52 = RG_rl_149 ;
	7'h78 :
		TR_52 = RG_rl_149 ;
	7'h79 :
		TR_52 = RG_rl_149 ;
	7'h7a :
		TR_52 = RG_rl_149 ;
	7'h7b :
		TR_52 = RG_rl_149 ;
	7'h7c :
		TR_52 = RG_rl_149 ;
	7'h7d :
		TR_52 = RG_rl_149 ;
	7'h7e :
		TR_52 = RG_rl_149 ;
	7'h7f :
		TR_52 = RG_rl_149 ;
	default :
		TR_52 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_18 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h01 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h02 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h03 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h04 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h05 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h06 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h07 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h08 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h09 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h0a :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h0b :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h0c :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h0d :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h0e :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h0f :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h10 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h11 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h12 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h13 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h14 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h15 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h16 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h17 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h18 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h19 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h1a :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h1b :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h1c :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h1d :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h1e :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h1f :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h20 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h21 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h22 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h23 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h24 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h25 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h26 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h27 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h28 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h29 :
		TR_53 = 9'h000 ;	// line#=../rle.cpp:79
	7'h2a :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h2b :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h2c :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h2d :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h2e :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h2f :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h30 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h31 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h32 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h33 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h34 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h35 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h36 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h37 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h38 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h39 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h3a :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h3b :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h3c :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h3d :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h3e :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h3f :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h40 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h41 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h42 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h43 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h44 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h45 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h46 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h47 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h48 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h49 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h4a :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h4b :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h4c :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h4d :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h4e :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h4f :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h50 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h51 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h52 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h53 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h54 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h55 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h56 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h57 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h58 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h59 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h5a :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h5b :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h5c :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h5d :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h5e :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h5f :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h60 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h61 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h62 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h63 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h64 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h65 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h66 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h67 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h68 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h69 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h6a :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h6b :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h6c :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h6d :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h6e :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h6f :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h70 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h71 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h72 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h73 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h74 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h75 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h76 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h77 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h78 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h79 :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h7a :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h7b :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h7c :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h7d :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h7e :
		TR_53 = RG_quantized_block_rl_18 ;
	7'h7f :
		TR_53 = RG_quantized_block_rl_18 ;
	default :
		TR_53 = 9'hx ;
	endcase
always @ ( RG_rl_150 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_54 = RG_rl_150 ;
	7'h01 :
		TR_54 = RG_rl_150 ;
	7'h02 :
		TR_54 = RG_rl_150 ;
	7'h03 :
		TR_54 = RG_rl_150 ;
	7'h04 :
		TR_54 = RG_rl_150 ;
	7'h05 :
		TR_54 = RG_rl_150 ;
	7'h06 :
		TR_54 = RG_rl_150 ;
	7'h07 :
		TR_54 = RG_rl_150 ;
	7'h08 :
		TR_54 = RG_rl_150 ;
	7'h09 :
		TR_54 = RG_rl_150 ;
	7'h0a :
		TR_54 = RG_rl_150 ;
	7'h0b :
		TR_54 = RG_rl_150 ;
	7'h0c :
		TR_54 = RG_rl_150 ;
	7'h0d :
		TR_54 = RG_rl_150 ;
	7'h0e :
		TR_54 = RG_rl_150 ;
	7'h0f :
		TR_54 = RG_rl_150 ;
	7'h10 :
		TR_54 = RG_rl_150 ;
	7'h11 :
		TR_54 = RG_rl_150 ;
	7'h12 :
		TR_54 = RG_rl_150 ;
	7'h13 :
		TR_54 = RG_rl_150 ;
	7'h14 :
		TR_54 = RG_rl_150 ;
	7'h15 :
		TR_54 = RG_rl_150 ;
	7'h16 :
		TR_54 = RG_rl_150 ;
	7'h17 :
		TR_54 = RG_rl_150 ;
	7'h18 :
		TR_54 = RG_rl_150 ;
	7'h19 :
		TR_54 = RG_rl_150 ;
	7'h1a :
		TR_54 = RG_rl_150 ;
	7'h1b :
		TR_54 = RG_rl_150 ;
	7'h1c :
		TR_54 = RG_rl_150 ;
	7'h1d :
		TR_54 = RG_rl_150 ;
	7'h1e :
		TR_54 = RG_rl_150 ;
	7'h1f :
		TR_54 = RG_rl_150 ;
	7'h20 :
		TR_54 = RG_rl_150 ;
	7'h21 :
		TR_54 = RG_rl_150 ;
	7'h22 :
		TR_54 = RG_rl_150 ;
	7'h23 :
		TR_54 = RG_rl_150 ;
	7'h24 :
		TR_54 = RG_rl_150 ;
	7'h25 :
		TR_54 = RG_rl_150 ;
	7'h26 :
		TR_54 = RG_rl_150 ;
	7'h27 :
		TR_54 = RG_rl_150 ;
	7'h28 :
		TR_54 = RG_rl_150 ;
	7'h29 :
		TR_54 = RG_rl_150 ;
	7'h2a :
		TR_54 = 9'h000 ;	// line#=../rle.cpp:79
	7'h2b :
		TR_54 = RG_rl_150 ;
	7'h2c :
		TR_54 = RG_rl_150 ;
	7'h2d :
		TR_54 = RG_rl_150 ;
	7'h2e :
		TR_54 = RG_rl_150 ;
	7'h2f :
		TR_54 = RG_rl_150 ;
	7'h30 :
		TR_54 = RG_rl_150 ;
	7'h31 :
		TR_54 = RG_rl_150 ;
	7'h32 :
		TR_54 = RG_rl_150 ;
	7'h33 :
		TR_54 = RG_rl_150 ;
	7'h34 :
		TR_54 = RG_rl_150 ;
	7'h35 :
		TR_54 = RG_rl_150 ;
	7'h36 :
		TR_54 = RG_rl_150 ;
	7'h37 :
		TR_54 = RG_rl_150 ;
	7'h38 :
		TR_54 = RG_rl_150 ;
	7'h39 :
		TR_54 = RG_rl_150 ;
	7'h3a :
		TR_54 = RG_rl_150 ;
	7'h3b :
		TR_54 = RG_rl_150 ;
	7'h3c :
		TR_54 = RG_rl_150 ;
	7'h3d :
		TR_54 = RG_rl_150 ;
	7'h3e :
		TR_54 = RG_rl_150 ;
	7'h3f :
		TR_54 = RG_rl_150 ;
	7'h40 :
		TR_54 = RG_rl_150 ;
	7'h41 :
		TR_54 = RG_rl_150 ;
	7'h42 :
		TR_54 = RG_rl_150 ;
	7'h43 :
		TR_54 = RG_rl_150 ;
	7'h44 :
		TR_54 = RG_rl_150 ;
	7'h45 :
		TR_54 = RG_rl_150 ;
	7'h46 :
		TR_54 = RG_rl_150 ;
	7'h47 :
		TR_54 = RG_rl_150 ;
	7'h48 :
		TR_54 = RG_rl_150 ;
	7'h49 :
		TR_54 = RG_rl_150 ;
	7'h4a :
		TR_54 = RG_rl_150 ;
	7'h4b :
		TR_54 = RG_rl_150 ;
	7'h4c :
		TR_54 = RG_rl_150 ;
	7'h4d :
		TR_54 = RG_rl_150 ;
	7'h4e :
		TR_54 = RG_rl_150 ;
	7'h4f :
		TR_54 = RG_rl_150 ;
	7'h50 :
		TR_54 = RG_rl_150 ;
	7'h51 :
		TR_54 = RG_rl_150 ;
	7'h52 :
		TR_54 = RG_rl_150 ;
	7'h53 :
		TR_54 = RG_rl_150 ;
	7'h54 :
		TR_54 = RG_rl_150 ;
	7'h55 :
		TR_54 = RG_rl_150 ;
	7'h56 :
		TR_54 = RG_rl_150 ;
	7'h57 :
		TR_54 = RG_rl_150 ;
	7'h58 :
		TR_54 = RG_rl_150 ;
	7'h59 :
		TR_54 = RG_rl_150 ;
	7'h5a :
		TR_54 = RG_rl_150 ;
	7'h5b :
		TR_54 = RG_rl_150 ;
	7'h5c :
		TR_54 = RG_rl_150 ;
	7'h5d :
		TR_54 = RG_rl_150 ;
	7'h5e :
		TR_54 = RG_rl_150 ;
	7'h5f :
		TR_54 = RG_rl_150 ;
	7'h60 :
		TR_54 = RG_rl_150 ;
	7'h61 :
		TR_54 = RG_rl_150 ;
	7'h62 :
		TR_54 = RG_rl_150 ;
	7'h63 :
		TR_54 = RG_rl_150 ;
	7'h64 :
		TR_54 = RG_rl_150 ;
	7'h65 :
		TR_54 = RG_rl_150 ;
	7'h66 :
		TR_54 = RG_rl_150 ;
	7'h67 :
		TR_54 = RG_rl_150 ;
	7'h68 :
		TR_54 = RG_rl_150 ;
	7'h69 :
		TR_54 = RG_rl_150 ;
	7'h6a :
		TR_54 = RG_rl_150 ;
	7'h6b :
		TR_54 = RG_rl_150 ;
	7'h6c :
		TR_54 = RG_rl_150 ;
	7'h6d :
		TR_54 = RG_rl_150 ;
	7'h6e :
		TR_54 = RG_rl_150 ;
	7'h6f :
		TR_54 = RG_rl_150 ;
	7'h70 :
		TR_54 = RG_rl_150 ;
	7'h71 :
		TR_54 = RG_rl_150 ;
	7'h72 :
		TR_54 = RG_rl_150 ;
	7'h73 :
		TR_54 = RG_rl_150 ;
	7'h74 :
		TR_54 = RG_rl_150 ;
	7'h75 :
		TR_54 = RG_rl_150 ;
	7'h76 :
		TR_54 = RG_rl_150 ;
	7'h77 :
		TR_54 = RG_rl_150 ;
	7'h78 :
		TR_54 = RG_rl_150 ;
	7'h79 :
		TR_54 = RG_rl_150 ;
	7'h7a :
		TR_54 = RG_rl_150 ;
	7'h7b :
		TR_54 = RG_rl_150 ;
	7'h7c :
		TR_54 = RG_rl_150 ;
	7'h7d :
		TR_54 = RG_rl_150 ;
	7'h7e :
		TR_54 = RG_rl_150 ;
	7'h7f :
		TR_54 = RG_rl_150 ;
	default :
		TR_54 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_19 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h01 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h02 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h03 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h04 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h05 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h06 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h07 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h08 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h09 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h0a :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h0b :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h0c :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h0d :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h0e :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h0f :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h10 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h11 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h12 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h13 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h14 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h15 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h16 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h17 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h18 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h19 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h1a :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h1b :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h1c :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h1d :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h1e :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h1f :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h20 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h21 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h22 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h23 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h24 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h25 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h26 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h27 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h28 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h29 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h2a :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h2b :
		TR_55 = 9'h000 ;	// line#=../rle.cpp:79
	7'h2c :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h2d :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h2e :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h2f :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h30 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h31 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h32 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h33 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h34 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h35 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h36 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h37 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h38 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h39 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h3a :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h3b :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h3c :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h3d :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h3e :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h3f :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h40 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h41 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h42 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h43 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h44 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h45 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h46 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h47 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h48 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h49 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h4a :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h4b :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h4c :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h4d :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h4e :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h4f :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h50 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h51 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h52 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h53 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h54 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h55 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h56 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h57 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h58 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h59 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h5a :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h5b :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h5c :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h5d :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h5e :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h5f :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h60 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h61 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h62 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h63 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h64 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h65 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h66 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h67 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h68 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h69 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h6a :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h6b :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h6c :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h6d :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h6e :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h6f :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h70 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h71 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h72 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h73 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h74 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h75 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h76 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h77 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h78 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h79 :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h7a :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h7b :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h7c :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h7d :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h7e :
		TR_55 = RG_quantized_block_rl_19 ;
	7'h7f :
		TR_55 = RG_quantized_block_rl_19 ;
	default :
		TR_55 = 9'hx ;
	endcase
always @ ( RG_rl_151 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_56 = RG_rl_151 ;
	7'h01 :
		TR_56 = RG_rl_151 ;
	7'h02 :
		TR_56 = RG_rl_151 ;
	7'h03 :
		TR_56 = RG_rl_151 ;
	7'h04 :
		TR_56 = RG_rl_151 ;
	7'h05 :
		TR_56 = RG_rl_151 ;
	7'h06 :
		TR_56 = RG_rl_151 ;
	7'h07 :
		TR_56 = RG_rl_151 ;
	7'h08 :
		TR_56 = RG_rl_151 ;
	7'h09 :
		TR_56 = RG_rl_151 ;
	7'h0a :
		TR_56 = RG_rl_151 ;
	7'h0b :
		TR_56 = RG_rl_151 ;
	7'h0c :
		TR_56 = RG_rl_151 ;
	7'h0d :
		TR_56 = RG_rl_151 ;
	7'h0e :
		TR_56 = RG_rl_151 ;
	7'h0f :
		TR_56 = RG_rl_151 ;
	7'h10 :
		TR_56 = RG_rl_151 ;
	7'h11 :
		TR_56 = RG_rl_151 ;
	7'h12 :
		TR_56 = RG_rl_151 ;
	7'h13 :
		TR_56 = RG_rl_151 ;
	7'h14 :
		TR_56 = RG_rl_151 ;
	7'h15 :
		TR_56 = RG_rl_151 ;
	7'h16 :
		TR_56 = RG_rl_151 ;
	7'h17 :
		TR_56 = RG_rl_151 ;
	7'h18 :
		TR_56 = RG_rl_151 ;
	7'h19 :
		TR_56 = RG_rl_151 ;
	7'h1a :
		TR_56 = RG_rl_151 ;
	7'h1b :
		TR_56 = RG_rl_151 ;
	7'h1c :
		TR_56 = RG_rl_151 ;
	7'h1d :
		TR_56 = RG_rl_151 ;
	7'h1e :
		TR_56 = RG_rl_151 ;
	7'h1f :
		TR_56 = RG_rl_151 ;
	7'h20 :
		TR_56 = RG_rl_151 ;
	7'h21 :
		TR_56 = RG_rl_151 ;
	7'h22 :
		TR_56 = RG_rl_151 ;
	7'h23 :
		TR_56 = RG_rl_151 ;
	7'h24 :
		TR_56 = RG_rl_151 ;
	7'h25 :
		TR_56 = RG_rl_151 ;
	7'h26 :
		TR_56 = RG_rl_151 ;
	7'h27 :
		TR_56 = RG_rl_151 ;
	7'h28 :
		TR_56 = RG_rl_151 ;
	7'h29 :
		TR_56 = RG_rl_151 ;
	7'h2a :
		TR_56 = RG_rl_151 ;
	7'h2b :
		TR_56 = RG_rl_151 ;
	7'h2c :
		TR_56 = 9'h000 ;	// line#=../rle.cpp:79
	7'h2d :
		TR_56 = RG_rl_151 ;
	7'h2e :
		TR_56 = RG_rl_151 ;
	7'h2f :
		TR_56 = RG_rl_151 ;
	7'h30 :
		TR_56 = RG_rl_151 ;
	7'h31 :
		TR_56 = RG_rl_151 ;
	7'h32 :
		TR_56 = RG_rl_151 ;
	7'h33 :
		TR_56 = RG_rl_151 ;
	7'h34 :
		TR_56 = RG_rl_151 ;
	7'h35 :
		TR_56 = RG_rl_151 ;
	7'h36 :
		TR_56 = RG_rl_151 ;
	7'h37 :
		TR_56 = RG_rl_151 ;
	7'h38 :
		TR_56 = RG_rl_151 ;
	7'h39 :
		TR_56 = RG_rl_151 ;
	7'h3a :
		TR_56 = RG_rl_151 ;
	7'h3b :
		TR_56 = RG_rl_151 ;
	7'h3c :
		TR_56 = RG_rl_151 ;
	7'h3d :
		TR_56 = RG_rl_151 ;
	7'h3e :
		TR_56 = RG_rl_151 ;
	7'h3f :
		TR_56 = RG_rl_151 ;
	7'h40 :
		TR_56 = RG_rl_151 ;
	7'h41 :
		TR_56 = RG_rl_151 ;
	7'h42 :
		TR_56 = RG_rl_151 ;
	7'h43 :
		TR_56 = RG_rl_151 ;
	7'h44 :
		TR_56 = RG_rl_151 ;
	7'h45 :
		TR_56 = RG_rl_151 ;
	7'h46 :
		TR_56 = RG_rl_151 ;
	7'h47 :
		TR_56 = RG_rl_151 ;
	7'h48 :
		TR_56 = RG_rl_151 ;
	7'h49 :
		TR_56 = RG_rl_151 ;
	7'h4a :
		TR_56 = RG_rl_151 ;
	7'h4b :
		TR_56 = RG_rl_151 ;
	7'h4c :
		TR_56 = RG_rl_151 ;
	7'h4d :
		TR_56 = RG_rl_151 ;
	7'h4e :
		TR_56 = RG_rl_151 ;
	7'h4f :
		TR_56 = RG_rl_151 ;
	7'h50 :
		TR_56 = RG_rl_151 ;
	7'h51 :
		TR_56 = RG_rl_151 ;
	7'h52 :
		TR_56 = RG_rl_151 ;
	7'h53 :
		TR_56 = RG_rl_151 ;
	7'h54 :
		TR_56 = RG_rl_151 ;
	7'h55 :
		TR_56 = RG_rl_151 ;
	7'h56 :
		TR_56 = RG_rl_151 ;
	7'h57 :
		TR_56 = RG_rl_151 ;
	7'h58 :
		TR_56 = RG_rl_151 ;
	7'h59 :
		TR_56 = RG_rl_151 ;
	7'h5a :
		TR_56 = RG_rl_151 ;
	7'h5b :
		TR_56 = RG_rl_151 ;
	7'h5c :
		TR_56 = RG_rl_151 ;
	7'h5d :
		TR_56 = RG_rl_151 ;
	7'h5e :
		TR_56 = RG_rl_151 ;
	7'h5f :
		TR_56 = RG_rl_151 ;
	7'h60 :
		TR_56 = RG_rl_151 ;
	7'h61 :
		TR_56 = RG_rl_151 ;
	7'h62 :
		TR_56 = RG_rl_151 ;
	7'h63 :
		TR_56 = RG_rl_151 ;
	7'h64 :
		TR_56 = RG_rl_151 ;
	7'h65 :
		TR_56 = RG_rl_151 ;
	7'h66 :
		TR_56 = RG_rl_151 ;
	7'h67 :
		TR_56 = RG_rl_151 ;
	7'h68 :
		TR_56 = RG_rl_151 ;
	7'h69 :
		TR_56 = RG_rl_151 ;
	7'h6a :
		TR_56 = RG_rl_151 ;
	7'h6b :
		TR_56 = RG_rl_151 ;
	7'h6c :
		TR_56 = RG_rl_151 ;
	7'h6d :
		TR_56 = RG_rl_151 ;
	7'h6e :
		TR_56 = RG_rl_151 ;
	7'h6f :
		TR_56 = RG_rl_151 ;
	7'h70 :
		TR_56 = RG_rl_151 ;
	7'h71 :
		TR_56 = RG_rl_151 ;
	7'h72 :
		TR_56 = RG_rl_151 ;
	7'h73 :
		TR_56 = RG_rl_151 ;
	7'h74 :
		TR_56 = RG_rl_151 ;
	7'h75 :
		TR_56 = RG_rl_151 ;
	7'h76 :
		TR_56 = RG_rl_151 ;
	7'h77 :
		TR_56 = RG_rl_151 ;
	7'h78 :
		TR_56 = RG_rl_151 ;
	7'h79 :
		TR_56 = RG_rl_151 ;
	7'h7a :
		TR_56 = RG_rl_151 ;
	7'h7b :
		TR_56 = RG_rl_151 ;
	7'h7c :
		TR_56 = RG_rl_151 ;
	7'h7d :
		TR_56 = RG_rl_151 ;
	7'h7e :
		TR_56 = RG_rl_151 ;
	7'h7f :
		TR_56 = RG_rl_151 ;
	default :
		TR_56 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_20 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h01 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h02 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h03 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h04 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h05 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h06 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h07 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h08 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h09 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h0a :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h0b :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h0c :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h0d :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h0e :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h0f :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h10 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h11 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h12 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h13 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h14 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h15 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h16 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h17 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h18 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h19 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h1a :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h1b :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h1c :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h1d :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h1e :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h1f :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h20 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h21 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h22 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h23 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h24 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h25 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h26 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h27 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h28 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h29 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h2a :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h2b :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h2c :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h2d :
		TR_57 = 9'h000 ;	// line#=../rle.cpp:79
	7'h2e :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h2f :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h30 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h31 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h32 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h33 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h34 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h35 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h36 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h37 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h38 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h39 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h3a :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h3b :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h3c :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h3d :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h3e :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h3f :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h40 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h41 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h42 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h43 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h44 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h45 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h46 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h47 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h48 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h49 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h4a :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h4b :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h4c :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h4d :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h4e :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h4f :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h50 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h51 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h52 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h53 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h54 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h55 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h56 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h57 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h58 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h59 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h5a :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h5b :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h5c :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h5d :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h5e :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h5f :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h60 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h61 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h62 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h63 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h64 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h65 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h66 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h67 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h68 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h69 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h6a :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h6b :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h6c :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h6d :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h6e :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h6f :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h70 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h71 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h72 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h73 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h74 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h75 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h76 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h77 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h78 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h79 :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h7a :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h7b :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h7c :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h7d :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h7e :
		TR_57 = RG_quantized_block_rl_20 ;
	7'h7f :
		TR_57 = RG_quantized_block_rl_20 ;
	default :
		TR_57 = 9'hx ;
	endcase
always @ ( RG_rl_152 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_58 = RG_rl_152 ;
	7'h01 :
		TR_58 = RG_rl_152 ;
	7'h02 :
		TR_58 = RG_rl_152 ;
	7'h03 :
		TR_58 = RG_rl_152 ;
	7'h04 :
		TR_58 = RG_rl_152 ;
	7'h05 :
		TR_58 = RG_rl_152 ;
	7'h06 :
		TR_58 = RG_rl_152 ;
	7'h07 :
		TR_58 = RG_rl_152 ;
	7'h08 :
		TR_58 = RG_rl_152 ;
	7'h09 :
		TR_58 = RG_rl_152 ;
	7'h0a :
		TR_58 = RG_rl_152 ;
	7'h0b :
		TR_58 = RG_rl_152 ;
	7'h0c :
		TR_58 = RG_rl_152 ;
	7'h0d :
		TR_58 = RG_rl_152 ;
	7'h0e :
		TR_58 = RG_rl_152 ;
	7'h0f :
		TR_58 = RG_rl_152 ;
	7'h10 :
		TR_58 = RG_rl_152 ;
	7'h11 :
		TR_58 = RG_rl_152 ;
	7'h12 :
		TR_58 = RG_rl_152 ;
	7'h13 :
		TR_58 = RG_rl_152 ;
	7'h14 :
		TR_58 = RG_rl_152 ;
	7'h15 :
		TR_58 = RG_rl_152 ;
	7'h16 :
		TR_58 = RG_rl_152 ;
	7'h17 :
		TR_58 = RG_rl_152 ;
	7'h18 :
		TR_58 = RG_rl_152 ;
	7'h19 :
		TR_58 = RG_rl_152 ;
	7'h1a :
		TR_58 = RG_rl_152 ;
	7'h1b :
		TR_58 = RG_rl_152 ;
	7'h1c :
		TR_58 = RG_rl_152 ;
	7'h1d :
		TR_58 = RG_rl_152 ;
	7'h1e :
		TR_58 = RG_rl_152 ;
	7'h1f :
		TR_58 = RG_rl_152 ;
	7'h20 :
		TR_58 = RG_rl_152 ;
	7'h21 :
		TR_58 = RG_rl_152 ;
	7'h22 :
		TR_58 = RG_rl_152 ;
	7'h23 :
		TR_58 = RG_rl_152 ;
	7'h24 :
		TR_58 = RG_rl_152 ;
	7'h25 :
		TR_58 = RG_rl_152 ;
	7'h26 :
		TR_58 = RG_rl_152 ;
	7'h27 :
		TR_58 = RG_rl_152 ;
	7'h28 :
		TR_58 = RG_rl_152 ;
	7'h29 :
		TR_58 = RG_rl_152 ;
	7'h2a :
		TR_58 = RG_rl_152 ;
	7'h2b :
		TR_58 = RG_rl_152 ;
	7'h2c :
		TR_58 = RG_rl_152 ;
	7'h2d :
		TR_58 = RG_rl_152 ;
	7'h2e :
		TR_58 = 9'h000 ;	// line#=../rle.cpp:79
	7'h2f :
		TR_58 = RG_rl_152 ;
	7'h30 :
		TR_58 = RG_rl_152 ;
	7'h31 :
		TR_58 = RG_rl_152 ;
	7'h32 :
		TR_58 = RG_rl_152 ;
	7'h33 :
		TR_58 = RG_rl_152 ;
	7'h34 :
		TR_58 = RG_rl_152 ;
	7'h35 :
		TR_58 = RG_rl_152 ;
	7'h36 :
		TR_58 = RG_rl_152 ;
	7'h37 :
		TR_58 = RG_rl_152 ;
	7'h38 :
		TR_58 = RG_rl_152 ;
	7'h39 :
		TR_58 = RG_rl_152 ;
	7'h3a :
		TR_58 = RG_rl_152 ;
	7'h3b :
		TR_58 = RG_rl_152 ;
	7'h3c :
		TR_58 = RG_rl_152 ;
	7'h3d :
		TR_58 = RG_rl_152 ;
	7'h3e :
		TR_58 = RG_rl_152 ;
	7'h3f :
		TR_58 = RG_rl_152 ;
	7'h40 :
		TR_58 = RG_rl_152 ;
	7'h41 :
		TR_58 = RG_rl_152 ;
	7'h42 :
		TR_58 = RG_rl_152 ;
	7'h43 :
		TR_58 = RG_rl_152 ;
	7'h44 :
		TR_58 = RG_rl_152 ;
	7'h45 :
		TR_58 = RG_rl_152 ;
	7'h46 :
		TR_58 = RG_rl_152 ;
	7'h47 :
		TR_58 = RG_rl_152 ;
	7'h48 :
		TR_58 = RG_rl_152 ;
	7'h49 :
		TR_58 = RG_rl_152 ;
	7'h4a :
		TR_58 = RG_rl_152 ;
	7'h4b :
		TR_58 = RG_rl_152 ;
	7'h4c :
		TR_58 = RG_rl_152 ;
	7'h4d :
		TR_58 = RG_rl_152 ;
	7'h4e :
		TR_58 = RG_rl_152 ;
	7'h4f :
		TR_58 = RG_rl_152 ;
	7'h50 :
		TR_58 = RG_rl_152 ;
	7'h51 :
		TR_58 = RG_rl_152 ;
	7'h52 :
		TR_58 = RG_rl_152 ;
	7'h53 :
		TR_58 = RG_rl_152 ;
	7'h54 :
		TR_58 = RG_rl_152 ;
	7'h55 :
		TR_58 = RG_rl_152 ;
	7'h56 :
		TR_58 = RG_rl_152 ;
	7'h57 :
		TR_58 = RG_rl_152 ;
	7'h58 :
		TR_58 = RG_rl_152 ;
	7'h59 :
		TR_58 = RG_rl_152 ;
	7'h5a :
		TR_58 = RG_rl_152 ;
	7'h5b :
		TR_58 = RG_rl_152 ;
	7'h5c :
		TR_58 = RG_rl_152 ;
	7'h5d :
		TR_58 = RG_rl_152 ;
	7'h5e :
		TR_58 = RG_rl_152 ;
	7'h5f :
		TR_58 = RG_rl_152 ;
	7'h60 :
		TR_58 = RG_rl_152 ;
	7'h61 :
		TR_58 = RG_rl_152 ;
	7'h62 :
		TR_58 = RG_rl_152 ;
	7'h63 :
		TR_58 = RG_rl_152 ;
	7'h64 :
		TR_58 = RG_rl_152 ;
	7'h65 :
		TR_58 = RG_rl_152 ;
	7'h66 :
		TR_58 = RG_rl_152 ;
	7'h67 :
		TR_58 = RG_rl_152 ;
	7'h68 :
		TR_58 = RG_rl_152 ;
	7'h69 :
		TR_58 = RG_rl_152 ;
	7'h6a :
		TR_58 = RG_rl_152 ;
	7'h6b :
		TR_58 = RG_rl_152 ;
	7'h6c :
		TR_58 = RG_rl_152 ;
	7'h6d :
		TR_58 = RG_rl_152 ;
	7'h6e :
		TR_58 = RG_rl_152 ;
	7'h6f :
		TR_58 = RG_rl_152 ;
	7'h70 :
		TR_58 = RG_rl_152 ;
	7'h71 :
		TR_58 = RG_rl_152 ;
	7'h72 :
		TR_58 = RG_rl_152 ;
	7'h73 :
		TR_58 = RG_rl_152 ;
	7'h74 :
		TR_58 = RG_rl_152 ;
	7'h75 :
		TR_58 = RG_rl_152 ;
	7'h76 :
		TR_58 = RG_rl_152 ;
	7'h77 :
		TR_58 = RG_rl_152 ;
	7'h78 :
		TR_58 = RG_rl_152 ;
	7'h79 :
		TR_58 = RG_rl_152 ;
	7'h7a :
		TR_58 = RG_rl_152 ;
	7'h7b :
		TR_58 = RG_rl_152 ;
	7'h7c :
		TR_58 = RG_rl_152 ;
	7'h7d :
		TR_58 = RG_rl_152 ;
	7'h7e :
		TR_58 = RG_rl_152 ;
	7'h7f :
		TR_58 = RG_rl_152 ;
	default :
		TR_58 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_21 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h01 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h02 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h03 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h04 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h05 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h06 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h07 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h08 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h09 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h0a :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h0b :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h0c :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h0d :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h0e :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h0f :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h10 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h11 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h12 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h13 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h14 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h15 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h16 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h17 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h18 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h19 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h1a :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h1b :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h1c :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h1d :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h1e :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h1f :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h20 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h21 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h22 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h23 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h24 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h25 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h26 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h27 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h28 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h29 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h2a :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h2b :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h2c :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h2d :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h2e :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h2f :
		TR_59 = 9'h000 ;	// line#=../rle.cpp:79
	7'h30 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h31 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h32 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h33 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h34 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h35 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h36 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h37 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h38 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h39 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h3a :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h3b :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h3c :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h3d :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h3e :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h3f :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h40 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h41 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h42 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h43 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h44 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h45 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h46 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h47 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h48 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h49 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h4a :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h4b :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h4c :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h4d :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h4e :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h4f :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h50 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h51 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h52 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h53 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h54 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h55 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h56 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h57 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h58 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h59 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h5a :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h5b :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h5c :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h5d :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h5e :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h5f :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h60 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h61 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h62 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h63 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h64 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h65 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h66 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h67 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h68 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h69 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h6a :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h6b :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h6c :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h6d :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h6e :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h6f :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h70 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h71 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h72 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h73 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h74 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h75 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h76 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h77 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h78 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h79 :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h7a :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h7b :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h7c :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h7d :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h7e :
		TR_59 = RG_quantized_block_rl_21 ;
	7'h7f :
		TR_59 = RG_quantized_block_rl_21 ;
	default :
		TR_59 = 9'hx ;
	endcase
always @ ( RG_rl_153 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_60 = RG_rl_153 ;
	7'h01 :
		TR_60 = RG_rl_153 ;
	7'h02 :
		TR_60 = RG_rl_153 ;
	7'h03 :
		TR_60 = RG_rl_153 ;
	7'h04 :
		TR_60 = RG_rl_153 ;
	7'h05 :
		TR_60 = RG_rl_153 ;
	7'h06 :
		TR_60 = RG_rl_153 ;
	7'h07 :
		TR_60 = RG_rl_153 ;
	7'h08 :
		TR_60 = RG_rl_153 ;
	7'h09 :
		TR_60 = RG_rl_153 ;
	7'h0a :
		TR_60 = RG_rl_153 ;
	7'h0b :
		TR_60 = RG_rl_153 ;
	7'h0c :
		TR_60 = RG_rl_153 ;
	7'h0d :
		TR_60 = RG_rl_153 ;
	7'h0e :
		TR_60 = RG_rl_153 ;
	7'h0f :
		TR_60 = RG_rl_153 ;
	7'h10 :
		TR_60 = RG_rl_153 ;
	7'h11 :
		TR_60 = RG_rl_153 ;
	7'h12 :
		TR_60 = RG_rl_153 ;
	7'h13 :
		TR_60 = RG_rl_153 ;
	7'h14 :
		TR_60 = RG_rl_153 ;
	7'h15 :
		TR_60 = RG_rl_153 ;
	7'h16 :
		TR_60 = RG_rl_153 ;
	7'h17 :
		TR_60 = RG_rl_153 ;
	7'h18 :
		TR_60 = RG_rl_153 ;
	7'h19 :
		TR_60 = RG_rl_153 ;
	7'h1a :
		TR_60 = RG_rl_153 ;
	7'h1b :
		TR_60 = RG_rl_153 ;
	7'h1c :
		TR_60 = RG_rl_153 ;
	7'h1d :
		TR_60 = RG_rl_153 ;
	7'h1e :
		TR_60 = RG_rl_153 ;
	7'h1f :
		TR_60 = RG_rl_153 ;
	7'h20 :
		TR_60 = RG_rl_153 ;
	7'h21 :
		TR_60 = RG_rl_153 ;
	7'h22 :
		TR_60 = RG_rl_153 ;
	7'h23 :
		TR_60 = RG_rl_153 ;
	7'h24 :
		TR_60 = RG_rl_153 ;
	7'h25 :
		TR_60 = RG_rl_153 ;
	7'h26 :
		TR_60 = RG_rl_153 ;
	7'h27 :
		TR_60 = RG_rl_153 ;
	7'h28 :
		TR_60 = RG_rl_153 ;
	7'h29 :
		TR_60 = RG_rl_153 ;
	7'h2a :
		TR_60 = RG_rl_153 ;
	7'h2b :
		TR_60 = RG_rl_153 ;
	7'h2c :
		TR_60 = RG_rl_153 ;
	7'h2d :
		TR_60 = RG_rl_153 ;
	7'h2e :
		TR_60 = RG_rl_153 ;
	7'h2f :
		TR_60 = RG_rl_153 ;
	7'h30 :
		TR_60 = 9'h000 ;	// line#=../rle.cpp:79
	7'h31 :
		TR_60 = RG_rl_153 ;
	7'h32 :
		TR_60 = RG_rl_153 ;
	7'h33 :
		TR_60 = RG_rl_153 ;
	7'h34 :
		TR_60 = RG_rl_153 ;
	7'h35 :
		TR_60 = RG_rl_153 ;
	7'h36 :
		TR_60 = RG_rl_153 ;
	7'h37 :
		TR_60 = RG_rl_153 ;
	7'h38 :
		TR_60 = RG_rl_153 ;
	7'h39 :
		TR_60 = RG_rl_153 ;
	7'h3a :
		TR_60 = RG_rl_153 ;
	7'h3b :
		TR_60 = RG_rl_153 ;
	7'h3c :
		TR_60 = RG_rl_153 ;
	7'h3d :
		TR_60 = RG_rl_153 ;
	7'h3e :
		TR_60 = RG_rl_153 ;
	7'h3f :
		TR_60 = RG_rl_153 ;
	7'h40 :
		TR_60 = RG_rl_153 ;
	7'h41 :
		TR_60 = RG_rl_153 ;
	7'h42 :
		TR_60 = RG_rl_153 ;
	7'h43 :
		TR_60 = RG_rl_153 ;
	7'h44 :
		TR_60 = RG_rl_153 ;
	7'h45 :
		TR_60 = RG_rl_153 ;
	7'h46 :
		TR_60 = RG_rl_153 ;
	7'h47 :
		TR_60 = RG_rl_153 ;
	7'h48 :
		TR_60 = RG_rl_153 ;
	7'h49 :
		TR_60 = RG_rl_153 ;
	7'h4a :
		TR_60 = RG_rl_153 ;
	7'h4b :
		TR_60 = RG_rl_153 ;
	7'h4c :
		TR_60 = RG_rl_153 ;
	7'h4d :
		TR_60 = RG_rl_153 ;
	7'h4e :
		TR_60 = RG_rl_153 ;
	7'h4f :
		TR_60 = RG_rl_153 ;
	7'h50 :
		TR_60 = RG_rl_153 ;
	7'h51 :
		TR_60 = RG_rl_153 ;
	7'h52 :
		TR_60 = RG_rl_153 ;
	7'h53 :
		TR_60 = RG_rl_153 ;
	7'h54 :
		TR_60 = RG_rl_153 ;
	7'h55 :
		TR_60 = RG_rl_153 ;
	7'h56 :
		TR_60 = RG_rl_153 ;
	7'h57 :
		TR_60 = RG_rl_153 ;
	7'h58 :
		TR_60 = RG_rl_153 ;
	7'h59 :
		TR_60 = RG_rl_153 ;
	7'h5a :
		TR_60 = RG_rl_153 ;
	7'h5b :
		TR_60 = RG_rl_153 ;
	7'h5c :
		TR_60 = RG_rl_153 ;
	7'h5d :
		TR_60 = RG_rl_153 ;
	7'h5e :
		TR_60 = RG_rl_153 ;
	7'h5f :
		TR_60 = RG_rl_153 ;
	7'h60 :
		TR_60 = RG_rl_153 ;
	7'h61 :
		TR_60 = RG_rl_153 ;
	7'h62 :
		TR_60 = RG_rl_153 ;
	7'h63 :
		TR_60 = RG_rl_153 ;
	7'h64 :
		TR_60 = RG_rl_153 ;
	7'h65 :
		TR_60 = RG_rl_153 ;
	7'h66 :
		TR_60 = RG_rl_153 ;
	7'h67 :
		TR_60 = RG_rl_153 ;
	7'h68 :
		TR_60 = RG_rl_153 ;
	7'h69 :
		TR_60 = RG_rl_153 ;
	7'h6a :
		TR_60 = RG_rl_153 ;
	7'h6b :
		TR_60 = RG_rl_153 ;
	7'h6c :
		TR_60 = RG_rl_153 ;
	7'h6d :
		TR_60 = RG_rl_153 ;
	7'h6e :
		TR_60 = RG_rl_153 ;
	7'h6f :
		TR_60 = RG_rl_153 ;
	7'h70 :
		TR_60 = RG_rl_153 ;
	7'h71 :
		TR_60 = RG_rl_153 ;
	7'h72 :
		TR_60 = RG_rl_153 ;
	7'h73 :
		TR_60 = RG_rl_153 ;
	7'h74 :
		TR_60 = RG_rl_153 ;
	7'h75 :
		TR_60 = RG_rl_153 ;
	7'h76 :
		TR_60 = RG_rl_153 ;
	7'h77 :
		TR_60 = RG_rl_153 ;
	7'h78 :
		TR_60 = RG_rl_153 ;
	7'h79 :
		TR_60 = RG_rl_153 ;
	7'h7a :
		TR_60 = RG_rl_153 ;
	7'h7b :
		TR_60 = RG_rl_153 ;
	7'h7c :
		TR_60 = RG_rl_153 ;
	7'h7d :
		TR_60 = RG_rl_153 ;
	7'h7e :
		TR_60 = RG_rl_153 ;
	7'h7f :
		TR_60 = RG_rl_153 ;
	default :
		TR_60 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_22 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h01 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h02 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h03 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h04 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h05 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h06 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h07 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h08 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h09 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h0a :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h0b :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h0c :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h0d :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h0e :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h0f :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h10 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h11 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h12 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h13 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h14 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h15 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h16 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h17 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h18 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h19 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h1a :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h1b :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h1c :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h1d :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h1e :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h1f :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h20 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h21 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h22 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h23 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h24 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h25 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h26 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h27 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h28 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h29 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h2a :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h2b :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h2c :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h2d :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h2e :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h2f :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h30 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h31 :
		TR_61 = 9'h000 ;	// line#=../rle.cpp:79
	7'h32 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h33 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h34 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h35 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h36 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h37 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h38 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h39 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h3a :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h3b :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h3c :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h3d :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h3e :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h3f :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h40 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h41 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h42 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h43 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h44 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h45 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h46 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h47 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h48 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h49 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h4a :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h4b :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h4c :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h4d :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h4e :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h4f :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h50 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h51 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h52 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h53 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h54 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h55 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h56 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h57 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h58 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h59 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h5a :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h5b :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h5c :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h5d :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h5e :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h5f :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h60 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h61 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h62 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h63 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h64 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h65 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h66 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h67 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h68 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h69 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h6a :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h6b :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h6c :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h6d :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h6e :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h6f :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h70 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h71 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h72 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h73 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h74 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h75 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h76 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h77 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h78 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h79 :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h7a :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h7b :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h7c :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h7d :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h7e :
		TR_61 = RG_quantized_block_rl_22 ;
	7'h7f :
		TR_61 = RG_quantized_block_rl_22 ;
	default :
		TR_61 = 9'hx ;
	endcase
always @ ( RG_rl_154 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_62 = RG_rl_154 ;
	7'h01 :
		TR_62 = RG_rl_154 ;
	7'h02 :
		TR_62 = RG_rl_154 ;
	7'h03 :
		TR_62 = RG_rl_154 ;
	7'h04 :
		TR_62 = RG_rl_154 ;
	7'h05 :
		TR_62 = RG_rl_154 ;
	7'h06 :
		TR_62 = RG_rl_154 ;
	7'h07 :
		TR_62 = RG_rl_154 ;
	7'h08 :
		TR_62 = RG_rl_154 ;
	7'h09 :
		TR_62 = RG_rl_154 ;
	7'h0a :
		TR_62 = RG_rl_154 ;
	7'h0b :
		TR_62 = RG_rl_154 ;
	7'h0c :
		TR_62 = RG_rl_154 ;
	7'h0d :
		TR_62 = RG_rl_154 ;
	7'h0e :
		TR_62 = RG_rl_154 ;
	7'h0f :
		TR_62 = RG_rl_154 ;
	7'h10 :
		TR_62 = RG_rl_154 ;
	7'h11 :
		TR_62 = RG_rl_154 ;
	7'h12 :
		TR_62 = RG_rl_154 ;
	7'h13 :
		TR_62 = RG_rl_154 ;
	7'h14 :
		TR_62 = RG_rl_154 ;
	7'h15 :
		TR_62 = RG_rl_154 ;
	7'h16 :
		TR_62 = RG_rl_154 ;
	7'h17 :
		TR_62 = RG_rl_154 ;
	7'h18 :
		TR_62 = RG_rl_154 ;
	7'h19 :
		TR_62 = RG_rl_154 ;
	7'h1a :
		TR_62 = RG_rl_154 ;
	7'h1b :
		TR_62 = RG_rl_154 ;
	7'h1c :
		TR_62 = RG_rl_154 ;
	7'h1d :
		TR_62 = RG_rl_154 ;
	7'h1e :
		TR_62 = RG_rl_154 ;
	7'h1f :
		TR_62 = RG_rl_154 ;
	7'h20 :
		TR_62 = RG_rl_154 ;
	7'h21 :
		TR_62 = RG_rl_154 ;
	7'h22 :
		TR_62 = RG_rl_154 ;
	7'h23 :
		TR_62 = RG_rl_154 ;
	7'h24 :
		TR_62 = RG_rl_154 ;
	7'h25 :
		TR_62 = RG_rl_154 ;
	7'h26 :
		TR_62 = RG_rl_154 ;
	7'h27 :
		TR_62 = RG_rl_154 ;
	7'h28 :
		TR_62 = RG_rl_154 ;
	7'h29 :
		TR_62 = RG_rl_154 ;
	7'h2a :
		TR_62 = RG_rl_154 ;
	7'h2b :
		TR_62 = RG_rl_154 ;
	7'h2c :
		TR_62 = RG_rl_154 ;
	7'h2d :
		TR_62 = RG_rl_154 ;
	7'h2e :
		TR_62 = RG_rl_154 ;
	7'h2f :
		TR_62 = RG_rl_154 ;
	7'h30 :
		TR_62 = RG_rl_154 ;
	7'h31 :
		TR_62 = RG_rl_154 ;
	7'h32 :
		TR_62 = 9'h000 ;	// line#=../rle.cpp:79
	7'h33 :
		TR_62 = RG_rl_154 ;
	7'h34 :
		TR_62 = RG_rl_154 ;
	7'h35 :
		TR_62 = RG_rl_154 ;
	7'h36 :
		TR_62 = RG_rl_154 ;
	7'h37 :
		TR_62 = RG_rl_154 ;
	7'h38 :
		TR_62 = RG_rl_154 ;
	7'h39 :
		TR_62 = RG_rl_154 ;
	7'h3a :
		TR_62 = RG_rl_154 ;
	7'h3b :
		TR_62 = RG_rl_154 ;
	7'h3c :
		TR_62 = RG_rl_154 ;
	7'h3d :
		TR_62 = RG_rl_154 ;
	7'h3e :
		TR_62 = RG_rl_154 ;
	7'h3f :
		TR_62 = RG_rl_154 ;
	7'h40 :
		TR_62 = RG_rl_154 ;
	7'h41 :
		TR_62 = RG_rl_154 ;
	7'h42 :
		TR_62 = RG_rl_154 ;
	7'h43 :
		TR_62 = RG_rl_154 ;
	7'h44 :
		TR_62 = RG_rl_154 ;
	7'h45 :
		TR_62 = RG_rl_154 ;
	7'h46 :
		TR_62 = RG_rl_154 ;
	7'h47 :
		TR_62 = RG_rl_154 ;
	7'h48 :
		TR_62 = RG_rl_154 ;
	7'h49 :
		TR_62 = RG_rl_154 ;
	7'h4a :
		TR_62 = RG_rl_154 ;
	7'h4b :
		TR_62 = RG_rl_154 ;
	7'h4c :
		TR_62 = RG_rl_154 ;
	7'h4d :
		TR_62 = RG_rl_154 ;
	7'h4e :
		TR_62 = RG_rl_154 ;
	7'h4f :
		TR_62 = RG_rl_154 ;
	7'h50 :
		TR_62 = RG_rl_154 ;
	7'h51 :
		TR_62 = RG_rl_154 ;
	7'h52 :
		TR_62 = RG_rl_154 ;
	7'h53 :
		TR_62 = RG_rl_154 ;
	7'h54 :
		TR_62 = RG_rl_154 ;
	7'h55 :
		TR_62 = RG_rl_154 ;
	7'h56 :
		TR_62 = RG_rl_154 ;
	7'h57 :
		TR_62 = RG_rl_154 ;
	7'h58 :
		TR_62 = RG_rl_154 ;
	7'h59 :
		TR_62 = RG_rl_154 ;
	7'h5a :
		TR_62 = RG_rl_154 ;
	7'h5b :
		TR_62 = RG_rl_154 ;
	7'h5c :
		TR_62 = RG_rl_154 ;
	7'h5d :
		TR_62 = RG_rl_154 ;
	7'h5e :
		TR_62 = RG_rl_154 ;
	7'h5f :
		TR_62 = RG_rl_154 ;
	7'h60 :
		TR_62 = RG_rl_154 ;
	7'h61 :
		TR_62 = RG_rl_154 ;
	7'h62 :
		TR_62 = RG_rl_154 ;
	7'h63 :
		TR_62 = RG_rl_154 ;
	7'h64 :
		TR_62 = RG_rl_154 ;
	7'h65 :
		TR_62 = RG_rl_154 ;
	7'h66 :
		TR_62 = RG_rl_154 ;
	7'h67 :
		TR_62 = RG_rl_154 ;
	7'h68 :
		TR_62 = RG_rl_154 ;
	7'h69 :
		TR_62 = RG_rl_154 ;
	7'h6a :
		TR_62 = RG_rl_154 ;
	7'h6b :
		TR_62 = RG_rl_154 ;
	7'h6c :
		TR_62 = RG_rl_154 ;
	7'h6d :
		TR_62 = RG_rl_154 ;
	7'h6e :
		TR_62 = RG_rl_154 ;
	7'h6f :
		TR_62 = RG_rl_154 ;
	7'h70 :
		TR_62 = RG_rl_154 ;
	7'h71 :
		TR_62 = RG_rl_154 ;
	7'h72 :
		TR_62 = RG_rl_154 ;
	7'h73 :
		TR_62 = RG_rl_154 ;
	7'h74 :
		TR_62 = RG_rl_154 ;
	7'h75 :
		TR_62 = RG_rl_154 ;
	7'h76 :
		TR_62 = RG_rl_154 ;
	7'h77 :
		TR_62 = RG_rl_154 ;
	7'h78 :
		TR_62 = RG_rl_154 ;
	7'h79 :
		TR_62 = RG_rl_154 ;
	7'h7a :
		TR_62 = RG_rl_154 ;
	7'h7b :
		TR_62 = RG_rl_154 ;
	7'h7c :
		TR_62 = RG_rl_154 ;
	7'h7d :
		TR_62 = RG_rl_154 ;
	7'h7e :
		TR_62 = RG_rl_154 ;
	7'h7f :
		TR_62 = RG_rl_154 ;
	default :
		TR_62 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_23 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h01 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h02 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h03 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h04 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h05 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h06 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h07 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h08 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h09 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h0a :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h0b :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h0c :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h0d :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h0e :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h0f :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h10 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h11 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h12 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h13 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h14 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h15 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h16 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h17 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h18 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h19 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h1a :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h1b :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h1c :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h1d :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h1e :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h1f :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h20 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h21 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h22 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h23 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h24 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h25 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h26 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h27 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h28 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h29 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h2a :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h2b :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h2c :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h2d :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h2e :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h2f :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h30 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h31 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h32 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h33 :
		TR_63 = 9'h000 ;	// line#=../rle.cpp:79
	7'h34 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h35 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h36 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h37 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h38 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h39 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h3a :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h3b :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h3c :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h3d :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h3e :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h3f :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h40 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h41 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h42 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h43 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h44 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h45 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h46 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h47 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h48 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h49 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h4a :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h4b :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h4c :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h4d :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h4e :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h4f :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h50 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h51 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h52 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h53 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h54 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h55 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h56 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h57 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h58 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h59 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h5a :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h5b :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h5c :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h5d :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h5e :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h5f :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h60 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h61 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h62 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h63 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h64 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h65 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h66 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h67 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h68 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h69 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h6a :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h6b :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h6c :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h6d :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h6e :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h6f :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h70 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h71 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h72 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h73 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h74 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h75 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h76 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h77 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h78 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h79 :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h7a :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h7b :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h7c :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h7d :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h7e :
		TR_63 = RG_quantized_block_rl_23 ;
	7'h7f :
		TR_63 = RG_quantized_block_rl_23 ;
	default :
		TR_63 = 9'hx ;
	endcase
always @ ( RG_rl_155 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_64 = RG_rl_155 ;
	7'h01 :
		TR_64 = RG_rl_155 ;
	7'h02 :
		TR_64 = RG_rl_155 ;
	7'h03 :
		TR_64 = RG_rl_155 ;
	7'h04 :
		TR_64 = RG_rl_155 ;
	7'h05 :
		TR_64 = RG_rl_155 ;
	7'h06 :
		TR_64 = RG_rl_155 ;
	7'h07 :
		TR_64 = RG_rl_155 ;
	7'h08 :
		TR_64 = RG_rl_155 ;
	7'h09 :
		TR_64 = RG_rl_155 ;
	7'h0a :
		TR_64 = RG_rl_155 ;
	7'h0b :
		TR_64 = RG_rl_155 ;
	7'h0c :
		TR_64 = RG_rl_155 ;
	7'h0d :
		TR_64 = RG_rl_155 ;
	7'h0e :
		TR_64 = RG_rl_155 ;
	7'h0f :
		TR_64 = RG_rl_155 ;
	7'h10 :
		TR_64 = RG_rl_155 ;
	7'h11 :
		TR_64 = RG_rl_155 ;
	7'h12 :
		TR_64 = RG_rl_155 ;
	7'h13 :
		TR_64 = RG_rl_155 ;
	7'h14 :
		TR_64 = RG_rl_155 ;
	7'h15 :
		TR_64 = RG_rl_155 ;
	7'h16 :
		TR_64 = RG_rl_155 ;
	7'h17 :
		TR_64 = RG_rl_155 ;
	7'h18 :
		TR_64 = RG_rl_155 ;
	7'h19 :
		TR_64 = RG_rl_155 ;
	7'h1a :
		TR_64 = RG_rl_155 ;
	7'h1b :
		TR_64 = RG_rl_155 ;
	7'h1c :
		TR_64 = RG_rl_155 ;
	7'h1d :
		TR_64 = RG_rl_155 ;
	7'h1e :
		TR_64 = RG_rl_155 ;
	7'h1f :
		TR_64 = RG_rl_155 ;
	7'h20 :
		TR_64 = RG_rl_155 ;
	7'h21 :
		TR_64 = RG_rl_155 ;
	7'h22 :
		TR_64 = RG_rl_155 ;
	7'h23 :
		TR_64 = RG_rl_155 ;
	7'h24 :
		TR_64 = RG_rl_155 ;
	7'h25 :
		TR_64 = RG_rl_155 ;
	7'h26 :
		TR_64 = RG_rl_155 ;
	7'h27 :
		TR_64 = RG_rl_155 ;
	7'h28 :
		TR_64 = RG_rl_155 ;
	7'h29 :
		TR_64 = RG_rl_155 ;
	7'h2a :
		TR_64 = RG_rl_155 ;
	7'h2b :
		TR_64 = RG_rl_155 ;
	7'h2c :
		TR_64 = RG_rl_155 ;
	7'h2d :
		TR_64 = RG_rl_155 ;
	7'h2e :
		TR_64 = RG_rl_155 ;
	7'h2f :
		TR_64 = RG_rl_155 ;
	7'h30 :
		TR_64 = RG_rl_155 ;
	7'h31 :
		TR_64 = RG_rl_155 ;
	7'h32 :
		TR_64 = RG_rl_155 ;
	7'h33 :
		TR_64 = RG_rl_155 ;
	7'h34 :
		TR_64 = 9'h000 ;	// line#=../rle.cpp:79
	7'h35 :
		TR_64 = RG_rl_155 ;
	7'h36 :
		TR_64 = RG_rl_155 ;
	7'h37 :
		TR_64 = RG_rl_155 ;
	7'h38 :
		TR_64 = RG_rl_155 ;
	7'h39 :
		TR_64 = RG_rl_155 ;
	7'h3a :
		TR_64 = RG_rl_155 ;
	7'h3b :
		TR_64 = RG_rl_155 ;
	7'h3c :
		TR_64 = RG_rl_155 ;
	7'h3d :
		TR_64 = RG_rl_155 ;
	7'h3e :
		TR_64 = RG_rl_155 ;
	7'h3f :
		TR_64 = RG_rl_155 ;
	7'h40 :
		TR_64 = RG_rl_155 ;
	7'h41 :
		TR_64 = RG_rl_155 ;
	7'h42 :
		TR_64 = RG_rl_155 ;
	7'h43 :
		TR_64 = RG_rl_155 ;
	7'h44 :
		TR_64 = RG_rl_155 ;
	7'h45 :
		TR_64 = RG_rl_155 ;
	7'h46 :
		TR_64 = RG_rl_155 ;
	7'h47 :
		TR_64 = RG_rl_155 ;
	7'h48 :
		TR_64 = RG_rl_155 ;
	7'h49 :
		TR_64 = RG_rl_155 ;
	7'h4a :
		TR_64 = RG_rl_155 ;
	7'h4b :
		TR_64 = RG_rl_155 ;
	7'h4c :
		TR_64 = RG_rl_155 ;
	7'h4d :
		TR_64 = RG_rl_155 ;
	7'h4e :
		TR_64 = RG_rl_155 ;
	7'h4f :
		TR_64 = RG_rl_155 ;
	7'h50 :
		TR_64 = RG_rl_155 ;
	7'h51 :
		TR_64 = RG_rl_155 ;
	7'h52 :
		TR_64 = RG_rl_155 ;
	7'h53 :
		TR_64 = RG_rl_155 ;
	7'h54 :
		TR_64 = RG_rl_155 ;
	7'h55 :
		TR_64 = RG_rl_155 ;
	7'h56 :
		TR_64 = RG_rl_155 ;
	7'h57 :
		TR_64 = RG_rl_155 ;
	7'h58 :
		TR_64 = RG_rl_155 ;
	7'h59 :
		TR_64 = RG_rl_155 ;
	7'h5a :
		TR_64 = RG_rl_155 ;
	7'h5b :
		TR_64 = RG_rl_155 ;
	7'h5c :
		TR_64 = RG_rl_155 ;
	7'h5d :
		TR_64 = RG_rl_155 ;
	7'h5e :
		TR_64 = RG_rl_155 ;
	7'h5f :
		TR_64 = RG_rl_155 ;
	7'h60 :
		TR_64 = RG_rl_155 ;
	7'h61 :
		TR_64 = RG_rl_155 ;
	7'h62 :
		TR_64 = RG_rl_155 ;
	7'h63 :
		TR_64 = RG_rl_155 ;
	7'h64 :
		TR_64 = RG_rl_155 ;
	7'h65 :
		TR_64 = RG_rl_155 ;
	7'h66 :
		TR_64 = RG_rl_155 ;
	7'h67 :
		TR_64 = RG_rl_155 ;
	7'h68 :
		TR_64 = RG_rl_155 ;
	7'h69 :
		TR_64 = RG_rl_155 ;
	7'h6a :
		TR_64 = RG_rl_155 ;
	7'h6b :
		TR_64 = RG_rl_155 ;
	7'h6c :
		TR_64 = RG_rl_155 ;
	7'h6d :
		TR_64 = RG_rl_155 ;
	7'h6e :
		TR_64 = RG_rl_155 ;
	7'h6f :
		TR_64 = RG_rl_155 ;
	7'h70 :
		TR_64 = RG_rl_155 ;
	7'h71 :
		TR_64 = RG_rl_155 ;
	7'h72 :
		TR_64 = RG_rl_155 ;
	7'h73 :
		TR_64 = RG_rl_155 ;
	7'h74 :
		TR_64 = RG_rl_155 ;
	7'h75 :
		TR_64 = RG_rl_155 ;
	7'h76 :
		TR_64 = RG_rl_155 ;
	7'h77 :
		TR_64 = RG_rl_155 ;
	7'h78 :
		TR_64 = RG_rl_155 ;
	7'h79 :
		TR_64 = RG_rl_155 ;
	7'h7a :
		TR_64 = RG_rl_155 ;
	7'h7b :
		TR_64 = RG_rl_155 ;
	7'h7c :
		TR_64 = RG_rl_155 ;
	7'h7d :
		TR_64 = RG_rl_155 ;
	7'h7e :
		TR_64 = RG_rl_155 ;
	7'h7f :
		TR_64 = RG_rl_155 ;
	default :
		TR_64 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_24 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h01 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h02 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h03 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h04 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h05 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h06 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h07 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h08 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h09 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h0a :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h0b :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h0c :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h0d :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h0e :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h0f :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h10 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h11 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h12 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h13 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h14 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h15 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h16 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h17 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h18 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h19 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h1a :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h1b :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h1c :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h1d :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h1e :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h1f :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h20 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h21 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h22 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h23 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h24 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h25 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h26 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h27 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h28 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h29 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h2a :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h2b :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h2c :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h2d :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h2e :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h2f :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h30 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h31 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h32 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h33 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h34 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h35 :
		TR_65 = 9'h000 ;	// line#=../rle.cpp:79
	7'h36 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h37 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h38 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h39 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h3a :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h3b :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h3c :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h3d :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h3e :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h3f :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h40 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h41 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h42 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h43 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h44 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h45 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h46 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h47 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h48 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h49 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h4a :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h4b :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h4c :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h4d :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h4e :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h4f :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h50 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h51 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h52 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h53 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h54 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h55 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h56 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h57 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h58 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h59 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h5a :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h5b :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h5c :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h5d :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h5e :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h5f :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h60 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h61 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h62 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h63 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h64 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h65 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h66 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h67 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h68 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h69 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h6a :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h6b :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h6c :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h6d :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h6e :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h6f :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h70 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h71 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h72 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h73 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h74 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h75 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h76 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h77 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h78 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h79 :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h7a :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h7b :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h7c :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h7d :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h7e :
		TR_65 = RG_quantized_block_rl_24 ;
	7'h7f :
		TR_65 = RG_quantized_block_rl_24 ;
	default :
		TR_65 = 9'hx ;
	endcase
always @ ( RG_rl_156 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_66 = RG_rl_156 ;
	7'h01 :
		TR_66 = RG_rl_156 ;
	7'h02 :
		TR_66 = RG_rl_156 ;
	7'h03 :
		TR_66 = RG_rl_156 ;
	7'h04 :
		TR_66 = RG_rl_156 ;
	7'h05 :
		TR_66 = RG_rl_156 ;
	7'h06 :
		TR_66 = RG_rl_156 ;
	7'h07 :
		TR_66 = RG_rl_156 ;
	7'h08 :
		TR_66 = RG_rl_156 ;
	7'h09 :
		TR_66 = RG_rl_156 ;
	7'h0a :
		TR_66 = RG_rl_156 ;
	7'h0b :
		TR_66 = RG_rl_156 ;
	7'h0c :
		TR_66 = RG_rl_156 ;
	7'h0d :
		TR_66 = RG_rl_156 ;
	7'h0e :
		TR_66 = RG_rl_156 ;
	7'h0f :
		TR_66 = RG_rl_156 ;
	7'h10 :
		TR_66 = RG_rl_156 ;
	7'h11 :
		TR_66 = RG_rl_156 ;
	7'h12 :
		TR_66 = RG_rl_156 ;
	7'h13 :
		TR_66 = RG_rl_156 ;
	7'h14 :
		TR_66 = RG_rl_156 ;
	7'h15 :
		TR_66 = RG_rl_156 ;
	7'h16 :
		TR_66 = RG_rl_156 ;
	7'h17 :
		TR_66 = RG_rl_156 ;
	7'h18 :
		TR_66 = RG_rl_156 ;
	7'h19 :
		TR_66 = RG_rl_156 ;
	7'h1a :
		TR_66 = RG_rl_156 ;
	7'h1b :
		TR_66 = RG_rl_156 ;
	7'h1c :
		TR_66 = RG_rl_156 ;
	7'h1d :
		TR_66 = RG_rl_156 ;
	7'h1e :
		TR_66 = RG_rl_156 ;
	7'h1f :
		TR_66 = RG_rl_156 ;
	7'h20 :
		TR_66 = RG_rl_156 ;
	7'h21 :
		TR_66 = RG_rl_156 ;
	7'h22 :
		TR_66 = RG_rl_156 ;
	7'h23 :
		TR_66 = RG_rl_156 ;
	7'h24 :
		TR_66 = RG_rl_156 ;
	7'h25 :
		TR_66 = RG_rl_156 ;
	7'h26 :
		TR_66 = RG_rl_156 ;
	7'h27 :
		TR_66 = RG_rl_156 ;
	7'h28 :
		TR_66 = RG_rl_156 ;
	7'h29 :
		TR_66 = RG_rl_156 ;
	7'h2a :
		TR_66 = RG_rl_156 ;
	7'h2b :
		TR_66 = RG_rl_156 ;
	7'h2c :
		TR_66 = RG_rl_156 ;
	7'h2d :
		TR_66 = RG_rl_156 ;
	7'h2e :
		TR_66 = RG_rl_156 ;
	7'h2f :
		TR_66 = RG_rl_156 ;
	7'h30 :
		TR_66 = RG_rl_156 ;
	7'h31 :
		TR_66 = RG_rl_156 ;
	7'h32 :
		TR_66 = RG_rl_156 ;
	7'h33 :
		TR_66 = RG_rl_156 ;
	7'h34 :
		TR_66 = RG_rl_156 ;
	7'h35 :
		TR_66 = RG_rl_156 ;
	7'h36 :
		TR_66 = 9'h000 ;	// line#=../rle.cpp:79
	7'h37 :
		TR_66 = RG_rl_156 ;
	7'h38 :
		TR_66 = RG_rl_156 ;
	7'h39 :
		TR_66 = RG_rl_156 ;
	7'h3a :
		TR_66 = RG_rl_156 ;
	7'h3b :
		TR_66 = RG_rl_156 ;
	7'h3c :
		TR_66 = RG_rl_156 ;
	7'h3d :
		TR_66 = RG_rl_156 ;
	7'h3e :
		TR_66 = RG_rl_156 ;
	7'h3f :
		TR_66 = RG_rl_156 ;
	7'h40 :
		TR_66 = RG_rl_156 ;
	7'h41 :
		TR_66 = RG_rl_156 ;
	7'h42 :
		TR_66 = RG_rl_156 ;
	7'h43 :
		TR_66 = RG_rl_156 ;
	7'h44 :
		TR_66 = RG_rl_156 ;
	7'h45 :
		TR_66 = RG_rl_156 ;
	7'h46 :
		TR_66 = RG_rl_156 ;
	7'h47 :
		TR_66 = RG_rl_156 ;
	7'h48 :
		TR_66 = RG_rl_156 ;
	7'h49 :
		TR_66 = RG_rl_156 ;
	7'h4a :
		TR_66 = RG_rl_156 ;
	7'h4b :
		TR_66 = RG_rl_156 ;
	7'h4c :
		TR_66 = RG_rl_156 ;
	7'h4d :
		TR_66 = RG_rl_156 ;
	7'h4e :
		TR_66 = RG_rl_156 ;
	7'h4f :
		TR_66 = RG_rl_156 ;
	7'h50 :
		TR_66 = RG_rl_156 ;
	7'h51 :
		TR_66 = RG_rl_156 ;
	7'h52 :
		TR_66 = RG_rl_156 ;
	7'h53 :
		TR_66 = RG_rl_156 ;
	7'h54 :
		TR_66 = RG_rl_156 ;
	7'h55 :
		TR_66 = RG_rl_156 ;
	7'h56 :
		TR_66 = RG_rl_156 ;
	7'h57 :
		TR_66 = RG_rl_156 ;
	7'h58 :
		TR_66 = RG_rl_156 ;
	7'h59 :
		TR_66 = RG_rl_156 ;
	7'h5a :
		TR_66 = RG_rl_156 ;
	7'h5b :
		TR_66 = RG_rl_156 ;
	7'h5c :
		TR_66 = RG_rl_156 ;
	7'h5d :
		TR_66 = RG_rl_156 ;
	7'h5e :
		TR_66 = RG_rl_156 ;
	7'h5f :
		TR_66 = RG_rl_156 ;
	7'h60 :
		TR_66 = RG_rl_156 ;
	7'h61 :
		TR_66 = RG_rl_156 ;
	7'h62 :
		TR_66 = RG_rl_156 ;
	7'h63 :
		TR_66 = RG_rl_156 ;
	7'h64 :
		TR_66 = RG_rl_156 ;
	7'h65 :
		TR_66 = RG_rl_156 ;
	7'h66 :
		TR_66 = RG_rl_156 ;
	7'h67 :
		TR_66 = RG_rl_156 ;
	7'h68 :
		TR_66 = RG_rl_156 ;
	7'h69 :
		TR_66 = RG_rl_156 ;
	7'h6a :
		TR_66 = RG_rl_156 ;
	7'h6b :
		TR_66 = RG_rl_156 ;
	7'h6c :
		TR_66 = RG_rl_156 ;
	7'h6d :
		TR_66 = RG_rl_156 ;
	7'h6e :
		TR_66 = RG_rl_156 ;
	7'h6f :
		TR_66 = RG_rl_156 ;
	7'h70 :
		TR_66 = RG_rl_156 ;
	7'h71 :
		TR_66 = RG_rl_156 ;
	7'h72 :
		TR_66 = RG_rl_156 ;
	7'h73 :
		TR_66 = RG_rl_156 ;
	7'h74 :
		TR_66 = RG_rl_156 ;
	7'h75 :
		TR_66 = RG_rl_156 ;
	7'h76 :
		TR_66 = RG_rl_156 ;
	7'h77 :
		TR_66 = RG_rl_156 ;
	7'h78 :
		TR_66 = RG_rl_156 ;
	7'h79 :
		TR_66 = RG_rl_156 ;
	7'h7a :
		TR_66 = RG_rl_156 ;
	7'h7b :
		TR_66 = RG_rl_156 ;
	7'h7c :
		TR_66 = RG_rl_156 ;
	7'h7d :
		TR_66 = RG_rl_156 ;
	7'h7e :
		TR_66 = RG_rl_156 ;
	7'h7f :
		TR_66 = RG_rl_156 ;
	default :
		TR_66 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_25 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h01 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h02 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h03 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h04 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h05 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h06 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h07 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h08 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h09 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h0a :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h0b :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h0c :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h0d :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h0e :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h0f :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h10 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h11 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h12 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h13 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h14 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h15 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h16 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h17 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h18 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h19 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h1a :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h1b :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h1c :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h1d :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h1e :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h1f :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h20 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h21 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h22 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h23 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h24 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h25 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h26 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h27 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h28 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h29 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h2a :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h2b :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h2c :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h2d :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h2e :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h2f :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h30 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h31 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h32 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h33 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h34 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h35 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h36 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h37 :
		TR_67 = 9'h000 ;	// line#=../rle.cpp:79
	7'h38 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h39 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h3a :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h3b :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h3c :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h3d :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h3e :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h3f :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h40 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h41 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h42 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h43 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h44 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h45 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h46 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h47 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h48 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h49 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h4a :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h4b :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h4c :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h4d :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h4e :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h4f :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h50 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h51 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h52 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h53 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h54 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h55 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h56 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h57 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h58 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h59 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h5a :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h5b :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h5c :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h5d :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h5e :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h5f :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h60 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h61 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h62 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h63 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h64 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h65 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h66 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h67 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h68 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h69 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h6a :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h6b :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h6c :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h6d :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h6e :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h6f :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h70 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h71 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h72 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h73 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h74 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h75 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h76 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h77 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h78 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h79 :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h7a :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h7b :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h7c :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h7d :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h7e :
		TR_67 = RG_quantized_block_rl_25 ;
	7'h7f :
		TR_67 = RG_quantized_block_rl_25 ;
	default :
		TR_67 = 9'hx ;
	endcase
always @ ( RG_rl_157 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_68 = RG_rl_157 ;
	7'h01 :
		TR_68 = RG_rl_157 ;
	7'h02 :
		TR_68 = RG_rl_157 ;
	7'h03 :
		TR_68 = RG_rl_157 ;
	7'h04 :
		TR_68 = RG_rl_157 ;
	7'h05 :
		TR_68 = RG_rl_157 ;
	7'h06 :
		TR_68 = RG_rl_157 ;
	7'h07 :
		TR_68 = RG_rl_157 ;
	7'h08 :
		TR_68 = RG_rl_157 ;
	7'h09 :
		TR_68 = RG_rl_157 ;
	7'h0a :
		TR_68 = RG_rl_157 ;
	7'h0b :
		TR_68 = RG_rl_157 ;
	7'h0c :
		TR_68 = RG_rl_157 ;
	7'h0d :
		TR_68 = RG_rl_157 ;
	7'h0e :
		TR_68 = RG_rl_157 ;
	7'h0f :
		TR_68 = RG_rl_157 ;
	7'h10 :
		TR_68 = RG_rl_157 ;
	7'h11 :
		TR_68 = RG_rl_157 ;
	7'h12 :
		TR_68 = RG_rl_157 ;
	7'h13 :
		TR_68 = RG_rl_157 ;
	7'h14 :
		TR_68 = RG_rl_157 ;
	7'h15 :
		TR_68 = RG_rl_157 ;
	7'h16 :
		TR_68 = RG_rl_157 ;
	7'h17 :
		TR_68 = RG_rl_157 ;
	7'h18 :
		TR_68 = RG_rl_157 ;
	7'h19 :
		TR_68 = RG_rl_157 ;
	7'h1a :
		TR_68 = RG_rl_157 ;
	7'h1b :
		TR_68 = RG_rl_157 ;
	7'h1c :
		TR_68 = RG_rl_157 ;
	7'h1d :
		TR_68 = RG_rl_157 ;
	7'h1e :
		TR_68 = RG_rl_157 ;
	7'h1f :
		TR_68 = RG_rl_157 ;
	7'h20 :
		TR_68 = RG_rl_157 ;
	7'h21 :
		TR_68 = RG_rl_157 ;
	7'h22 :
		TR_68 = RG_rl_157 ;
	7'h23 :
		TR_68 = RG_rl_157 ;
	7'h24 :
		TR_68 = RG_rl_157 ;
	7'h25 :
		TR_68 = RG_rl_157 ;
	7'h26 :
		TR_68 = RG_rl_157 ;
	7'h27 :
		TR_68 = RG_rl_157 ;
	7'h28 :
		TR_68 = RG_rl_157 ;
	7'h29 :
		TR_68 = RG_rl_157 ;
	7'h2a :
		TR_68 = RG_rl_157 ;
	7'h2b :
		TR_68 = RG_rl_157 ;
	7'h2c :
		TR_68 = RG_rl_157 ;
	7'h2d :
		TR_68 = RG_rl_157 ;
	7'h2e :
		TR_68 = RG_rl_157 ;
	7'h2f :
		TR_68 = RG_rl_157 ;
	7'h30 :
		TR_68 = RG_rl_157 ;
	7'h31 :
		TR_68 = RG_rl_157 ;
	7'h32 :
		TR_68 = RG_rl_157 ;
	7'h33 :
		TR_68 = RG_rl_157 ;
	7'h34 :
		TR_68 = RG_rl_157 ;
	7'h35 :
		TR_68 = RG_rl_157 ;
	7'h36 :
		TR_68 = RG_rl_157 ;
	7'h37 :
		TR_68 = RG_rl_157 ;
	7'h38 :
		TR_68 = 9'h000 ;	// line#=../rle.cpp:79
	7'h39 :
		TR_68 = RG_rl_157 ;
	7'h3a :
		TR_68 = RG_rl_157 ;
	7'h3b :
		TR_68 = RG_rl_157 ;
	7'h3c :
		TR_68 = RG_rl_157 ;
	7'h3d :
		TR_68 = RG_rl_157 ;
	7'h3e :
		TR_68 = RG_rl_157 ;
	7'h3f :
		TR_68 = RG_rl_157 ;
	7'h40 :
		TR_68 = RG_rl_157 ;
	7'h41 :
		TR_68 = RG_rl_157 ;
	7'h42 :
		TR_68 = RG_rl_157 ;
	7'h43 :
		TR_68 = RG_rl_157 ;
	7'h44 :
		TR_68 = RG_rl_157 ;
	7'h45 :
		TR_68 = RG_rl_157 ;
	7'h46 :
		TR_68 = RG_rl_157 ;
	7'h47 :
		TR_68 = RG_rl_157 ;
	7'h48 :
		TR_68 = RG_rl_157 ;
	7'h49 :
		TR_68 = RG_rl_157 ;
	7'h4a :
		TR_68 = RG_rl_157 ;
	7'h4b :
		TR_68 = RG_rl_157 ;
	7'h4c :
		TR_68 = RG_rl_157 ;
	7'h4d :
		TR_68 = RG_rl_157 ;
	7'h4e :
		TR_68 = RG_rl_157 ;
	7'h4f :
		TR_68 = RG_rl_157 ;
	7'h50 :
		TR_68 = RG_rl_157 ;
	7'h51 :
		TR_68 = RG_rl_157 ;
	7'h52 :
		TR_68 = RG_rl_157 ;
	7'h53 :
		TR_68 = RG_rl_157 ;
	7'h54 :
		TR_68 = RG_rl_157 ;
	7'h55 :
		TR_68 = RG_rl_157 ;
	7'h56 :
		TR_68 = RG_rl_157 ;
	7'h57 :
		TR_68 = RG_rl_157 ;
	7'h58 :
		TR_68 = RG_rl_157 ;
	7'h59 :
		TR_68 = RG_rl_157 ;
	7'h5a :
		TR_68 = RG_rl_157 ;
	7'h5b :
		TR_68 = RG_rl_157 ;
	7'h5c :
		TR_68 = RG_rl_157 ;
	7'h5d :
		TR_68 = RG_rl_157 ;
	7'h5e :
		TR_68 = RG_rl_157 ;
	7'h5f :
		TR_68 = RG_rl_157 ;
	7'h60 :
		TR_68 = RG_rl_157 ;
	7'h61 :
		TR_68 = RG_rl_157 ;
	7'h62 :
		TR_68 = RG_rl_157 ;
	7'h63 :
		TR_68 = RG_rl_157 ;
	7'h64 :
		TR_68 = RG_rl_157 ;
	7'h65 :
		TR_68 = RG_rl_157 ;
	7'h66 :
		TR_68 = RG_rl_157 ;
	7'h67 :
		TR_68 = RG_rl_157 ;
	7'h68 :
		TR_68 = RG_rl_157 ;
	7'h69 :
		TR_68 = RG_rl_157 ;
	7'h6a :
		TR_68 = RG_rl_157 ;
	7'h6b :
		TR_68 = RG_rl_157 ;
	7'h6c :
		TR_68 = RG_rl_157 ;
	7'h6d :
		TR_68 = RG_rl_157 ;
	7'h6e :
		TR_68 = RG_rl_157 ;
	7'h6f :
		TR_68 = RG_rl_157 ;
	7'h70 :
		TR_68 = RG_rl_157 ;
	7'h71 :
		TR_68 = RG_rl_157 ;
	7'h72 :
		TR_68 = RG_rl_157 ;
	7'h73 :
		TR_68 = RG_rl_157 ;
	7'h74 :
		TR_68 = RG_rl_157 ;
	7'h75 :
		TR_68 = RG_rl_157 ;
	7'h76 :
		TR_68 = RG_rl_157 ;
	7'h77 :
		TR_68 = RG_rl_157 ;
	7'h78 :
		TR_68 = RG_rl_157 ;
	7'h79 :
		TR_68 = RG_rl_157 ;
	7'h7a :
		TR_68 = RG_rl_157 ;
	7'h7b :
		TR_68 = RG_rl_157 ;
	7'h7c :
		TR_68 = RG_rl_157 ;
	7'h7d :
		TR_68 = RG_rl_157 ;
	7'h7e :
		TR_68 = RG_rl_157 ;
	7'h7f :
		TR_68 = RG_rl_157 ;
	default :
		TR_68 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_26 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h01 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h02 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h03 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h04 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h05 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h06 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h07 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h08 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h09 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h0a :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h0b :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h0c :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h0d :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h0e :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h0f :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h10 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h11 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h12 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h13 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h14 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h15 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h16 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h17 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h18 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h19 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h1a :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h1b :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h1c :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h1d :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h1e :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h1f :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h20 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h21 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h22 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h23 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h24 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h25 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h26 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h27 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h28 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h29 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h2a :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h2b :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h2c :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h2d :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h2e :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h2f :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h30 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h31 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h32 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h33 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h34 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h35 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h36 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h37 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h38 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h39 :
		TR_69 = 9'h000 ;	// line#=../rle.cpp:79
	7'h3a :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h3b :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h3c :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h3d :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h3e :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h3f :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h40 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h41 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h42 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h43 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h44 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h45 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h46 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h47 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h48 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h49 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h4a :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h4b :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h4c :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h4d :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h4e :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h4f :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h50 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h51 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h52 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h53 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h54 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h55 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h56 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h57 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h58 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h59 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h5a :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h5b :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h5c :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h5d :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h5e :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h5f :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h60 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h61 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h62 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h63 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h64 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h65 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h66 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h67 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h68 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h69 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h6a :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h6b :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h6c :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h6d :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h6e :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h6f :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h70 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h71 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h72 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h73 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h74 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h75 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h76 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h77 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h78 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h79 :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h7a :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h7b :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h7c :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h7d :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h7e :
		TR_69 = RG_quantized_block_rl_26 ;
	7'h7f :
		TR_69 = RG_quantized_block_rl_26 ;
	default :
		TR_69 = 9'hx ;
	endcase
always @ ( RG_rl_158 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_70 = RG_rl_158 ;
	7'h01 :
		TR_70 = RG_rl_158 ;
	7'h02 :
		TR_70 = RG_rl_158 ;
	7'h03 :
		TR_70 = RG_rl_158 ;
	7'h04 :
		TR_70 = RG_rl_158 ;
	7'h05 :
		TR_70 = RG_rl_158 ;
	7'h06 :
		TR_70 = RG_rl_158 ;
	7'h07 :
		TR_70 = RG_rl_158 ;
	7'h08 :
		TR_70 = RG_rl_158 ;
	7'h09 :
		TR_70 = RG_rl_158 ;
	7'h0a :
		TR_70 = RG_rl_158 ;
	7'h0b :
		TR_70 = RG_rl_158 ;
	7'h0c :
		TR_70 = RG_rl_158 ;
	7'h0d :
		TR_70 = RG_rl_158 ;
	7'h0e :
		TR_70 = RG_rl_158 ;
	7'h0f :
		TR_70 = RG_rl_158 ;
	7'h10 :
		TR_70 = RG_rl_158 ;
	7'h11 :
		TR_70 = RG_rl_158 ;
	7'h12 :
		TR_70 = RG_rl_158 ;
	7'h13 :
		TR_70 = RG_rl_158 ;
	7'h14 :
		TR_70 = RG_rl_158 ;
	7'h15 :
		TR_70 = RG_rl_158 ;
	7'h16 :
		TR_70 = RG_rl_158 ;
	7'h17 :
		TR_70 = RG_rl_158 ;
	7'h18 :
		TR_70 = RG_rl_158 ;
	7'h19 :
		TR_70 = RG_rl_158 ;
	7'h1a :
		TR_70 = RG_rl_158 ;
	7'h1b :
		TR_70 = RG_rl_158 ;
	7'h1c :
		TR_70 = RG_rl_158 ;
	7'h1d :
		TR_70 = RG_rl_158 ;
	7'h1e :
		TR_70 = RG_rl_158 ;
	7'h1f :
		TR_70 = RG_rl_158 ;
	7'h20 :
		TR_70 = RG_rl_158 ;
	7'h21 :
		TR_70 = RG_rl_158 ;
	7'h22 :
		TR_70 = RG_rl_158 ;
	7'h23 :
		TR_70 = RG_rl_158 ;
	7'h24 :
		TR_70 = RG_rl_158 ;
	7'h25 :
		TR_70 = RG_rl_158 ;
	7'h26 :
		TR_70 = RG_rl_158 ;
	7'h27 :
		TR_70 = RG_rl_158 ;
	7'h28 :
		TR_70 = RG_rl_158 ;
	7'h29 :
		TR_70 = RG_rl_158 ;
	7'h2a :
		TR_70 = RG_rl_158 ;
	7'h2b :
		TR_70 = RG_rl_158 ;
	7'h2c :
		TR_70 = RG_rl_158 ;
	7'h2d :
		TR_70 = RG_rl_158 ;
	7'h2e :
		TR_70 = RG_rl_158 ;
	7'h2f :
		TR_70 = RG_rl_158 ;
	7'h30 :
		TR_70 = RG_rl_158 ;
	7'h31 :
		TR_70 = RG_rl_158 ;
	7'h32 :
		TR_70 = RG_rl_158 ;
	7'h33 :
		TR_70 = RG_rl_158 ;
	7'h34 :
		TR_70 = RG_rl_158 ;
	7'h35 :
		TR_70 = RG_rl_158 ;
	7'h36 :
		TR_70 = RG_rl_158 ;
	7'h37 :
		TR_70 = RG_rl_158 ;
	7'h38 :
		TR_70 = RG_rl_158 ;
	7'h39 :
		TR_70 = RG_rl_158 ;
	7'h3a :
		TR_70 = 9'h000 ;	// line#=../rle.cpp:79
	7'h3b :
		TR_70 = RG_rl_158 ;
	7'h3c :
		TR_70 = RG_rl_158 ;
	7'h3d :
		TR_70 = RG_rl_158 ;
	7'h3e :
		TR_70 = RG_rl_158 ;
	7'h3f :
		TR_70 = RG_rl_158 ;
	7'h40 :
		TR_70 = RG_rl_158 ;
	7'h41 :
		TR_70 = RG_rl_158 ;
	7'h42 :
		TR_70 = RG_rl_158 ;
	7'h43 :
		TR_70 = RG_rl_158 ;
	7'h44 :
		TR_70 = RG_rl_158 ;
	7'h45 :
		TR_70 = RG_rl_158 ;
	7'h46 :
		TR_70 = RG_rl_158 ;
	7'h47 :
		TR_70 = RG_rl_158 ;
	7'h48 :
		TR_70 = RG_rl_158 ;
	7'h49 :
		TR_70 = RG_rl_158 ;
	7'h4a :
		TR_70 = RG_rl_158 ;
	7'h4b :
		TR_70 = RG_rl_158 ;
	7'h4c :
		TR_70 = RG_rl_158 ;
	7'h4d :
		TR_70 = RG_rl_158 ;
	7'h4e :
		TR_70 = RG_rl_158 ;
	7'h4f :
		TR_70 = RG_rl_158 ;
	7'h50 :
		TR_70 = RG_rl_158 ;
	7'h51 :
		TR_70 = RG_rl_158 ;
	7'h52 :
		TR_70 = RG_rl_158 ;
	7'h53 :
		TR_70 = RG_rl_158 ;
	7'h54 :
		TR_70 = RG_rl_158 ;
	7'h55 :
		TR_70 = RG_rl_158 ;
	7'h56 :
		TR_70 = RG_rl_158 ;
	7'h57 :
		TR_70 = RG_rl_158 ;
	7'h58 :
		TR_70 = RG_rl_158 ;
	7'h59 :
		TR_70 = RG_rl_158 ;
	7'h5a :
		TR_70 = RG_rl_158 ;
	7'h5b :
		TR_70 = RG_rl_158 ;
	7'h5c :
		TR_70 = RG_rl_158 ;
	7'h5d :
		TR_70 = RG_rl_158 ;
	7'h5e :
		TR_70 = RG_rl_158 ;
	7'h5f :
		TR_70 = RG_rl_158 ;
	7'h60 :
		TR_70 = RG_rl_158 ;
	7'h61 :
		TR_70 = RG_rl_158 ;
	7'h62 :
		TR_70 = RG_rl_158 ;
	7'h63 :
		TR_70 = RG_rl_158 ;
	7'h64 :
		TR_70 = RG_rl_158 ;
	7'h65 :
		TR_70 = RG_rl_158 ;
	7'h66 :
		TR_70 = RG_rl_158 ;
	7'h67 :
		TR_70 = RG_rl_158 ;
	7'h68 :
		TR_70 = RG_rl_158 ;
	7'h69 :
		TR_70 = RG_rl_158 ;
	7'h6a :
		TR_70 = RG_rl_158 ;
	7'h6b :
		TR_70 = RG_rl_158 ;
	7'h6c :
		TR_70 = RG_rl_158 ;
	7'h6d :
		TR_70 = RG_rl_158 ;
	7'h6e :
		TR_70 = RG_rl_158 ;
	7'h6f :
		TR_70 = RG_rl_158 ;
	7'h70 :
		TR_70 = RG_rl_158 ;
	7'h71 :
		TR_70 = RG_rl_158 ;
	7'h72 :
		TR_70 = RG_rl_158 ;
	7'h73 :
		TR_70 = RG_rl_158 ;
	7'h74 :
		TR_70 = RG_rl_158 ;
	7'h75 :
		TR_70 = RG_rl_158 ;
	7'h76 :
		TR_70 = RG_rl_158 ;
	7'h77 :
		TR_70 = RG_rl_158 ;
	7'h78 :
		TR_70 = RG_rl_158 ;
	7'h79 :
		TR_70 = RG_rl_158 ;
	7'h7a :
		TR_70 = RG_rl_158 ;
	7'h7b :
		TR_70 = RG_rl_158 ;
	7'h7c :
		TR_70 = RG_rl_158 ;
	7'h7d :
		TR_70 = RG_rl_158 ;
	7'h7e :
		TR_70 = RG_rl_158 ;
	7'h7f :
		TR_70 = RG_rl_158 ;
	default :
		TR_70 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_27 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h01 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h02 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h03 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h04 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h05 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h06 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h07 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h08 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h09 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h0a :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h0b :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h0c :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h0d :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h0e :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h0f :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h10 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h11 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h12 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h13 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h14 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h15 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h16 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h17 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h18 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h19 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h1a :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h1b :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h1c :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h1d :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h1e :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h1f :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h20 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h21 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h22 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h23 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h24 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h25 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h26 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h27 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h28 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h29 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h2a :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h2b :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h2c :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h2d :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h2e :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h2f :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h30 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h31 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h32 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h33 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h34 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h35 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h36 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h37 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h38 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h39 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h3a :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h3b :
		TR_71 = 9'h000 ;	// line#=../rle.cpp:79
	7'h3c :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h3d :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h3e :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h3f :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h40 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h41 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h42 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h43 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h44 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h45 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h46 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h47 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h48 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h49 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h4a :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h4b :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h4c :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h4d :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h4e :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h4f :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h50 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h51 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h52 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h53 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h54 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h55 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h56 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h57 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h58 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h59 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h5a :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h5b :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h5c :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h5d :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h5e :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h5f :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h60 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h61 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h62 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h63 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h64 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h65 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h66 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h67 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h68 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h69 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h6a :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h6b :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h6c :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h6d :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h6e :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h6f :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h70 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h71 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h72 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h73 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h74 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h75 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h76 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h77 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h78 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h79 :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h7a :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h7b :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h7c :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h7d :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h7e :
		TR_71 = RG_quantized_block_rl_27 ;
	7'h7f :
		TR_71 = RG_quantized_block_rl_27 ;
	default :
		TR_71 = 9'hx ;
	endcase
always @ ( RG_rl_159 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_72 = RG_rl_159 ;
	7'h01 :
		TR_72 = RG_rl_159 ;
	7'h02 :
		TR_72 = RG_rl_159 ;
	7'h03 :
		TR_72 = RG_rl_159 ;
	7'h04 :
		TR_72 = RG_rl_159 ;
	7'h05 :
		TR_72 = RG_rl_159 ;
	7'h06 :
		TR_72 = RG_rl_159 ;
	7'h07 :
		TR_72 = RG_rl_159 ;
	7'h08 :
		TR_72 = RG_rl_159 ;
	7'h09 :
		TR_72 = RG_rl_159 ;
	7'h0a :
		TR_72 = RG_rl_159 ;
	7'h0b :
		TR_72 = RG_rl_159 ;
	7'h0c :
		TR_72 = RG_rl_159 ;
	7'h0d :
		TR_72 = RG_rl_159 ;
	7'h0e :
		TR_72 = RG_rl_159 ;
	7'h0f :
		TR_72 = RG_rl_159 ;
	7'h10 :
		TR_72 = RG_rl_159 ;
	7'h11 :
		TR_72 = RG_rl_159 ;
	7'h12 :
		TR_72 = RG_rl_159 ;
	7'h13 :
		TR_72 = RG_rl_159 ;
	7'h14 :
		TR_72 = RG_rl_159 ;
	7'h15 :
		TR_72 = RG_rl_159 ;
	7'h16 :
		TR_72 = RG_rl_159 ;
	7'h17 :
		TR_72 = RG_rl_159 ;
	7'h18 :
		TR_72 = RG_rl_159 ;
	7'h19 :
		TR_72 = RG_rl_159 ;
	7'h1a :
		TR_72 = RG_rl_159 ;
	7'h1b :
		TR_72 = RG_rl_159 ;
	7'h1c :
		TR_72 = RG_rl_159 ;
	7'h1d :
		TR_72 = RG_rl_159 ;
	7'h1e :
		TR_72 = RG_rl_159 ;
	7'h1f :
		TR_72 = RG_rl_159 ;
	7'h20 :
		TR_72 = RG_rl_159 ;
	7'h21 :
		TR_72 = RG_rl_159 ;
	7'h22 :
		TR_72 = RG_rl_159 ;
	7'h23 :
		TR_72 = RG_rl_159 ;
	7'h24 :
		TR_72 = RG_rl_159 ;
	7'h25 :
		TR_72 = RG_rl_159 ;
	7'h26 :
		TR_72 = RG_rl_159 ;
	7'h27 :
		TR_72 = RG_rl_159 ;
	7'h28 :
		TR_72 = RG_rl_159 ;
	7'h29 :
		TR_72 = RG_rl_159 ;
	7'h2a :
		TR_72 = RG_rl_159 ;
	7'h2b :
		TR_72 = RG_rl_159 ;
	7'h2c :
		TR_72 = RG_rl_159 ;
	7'h2d :
		TR_72 = RG_rl_159 ;
	7'h2e :
		TR_72 = RG_rl_159 ;
	7'h2f :
		TR_72 = RG_rl_159 ;
	7'h30 :
		TR_72 = RG_rl_159 ;
	7'h31 :
		TR_72 = RG_rl_159 ;
	7'h32 :
		TR_72 = RG_rl_159 ;
	7'h33 :
		TR_72 = RG_rl_159 ;
	7'h34 :
		TR_72 = RG_rl_159 ;
	7'h35 :
		TR_72 = RG_rl_159 ;
	7'h36 :
		TR_72 = RG_rl_159 ;
	7'h37 :
		TR_72 = RG_rl_159 ;
	7'h38 :
		TR_72 = RG_rl_159 ;
	7'h39 :
		TR_72 = RG_rl_159 ;
	7'h3a :
		TR_72 = RG_rl_159 ;
	7'h3b :
		TR_72 = RG_rl_159 ;
	7'h3c :
		TR_72 = 9'h000 ;	// line#=../rle.cpp:79
	7'h3d :
		TR_72 = RG_rl_159 ;
	7'h3e :
		TR_72 = RG_rl_159 ;
	7'h3f :
		TR_72 = RG_rl_159 ;
	7'h40 :
		TR_72 = RG_rl_159 ;
	7'h41 :
		TR_72 = RG_rl_159 ;
	7'h42 :
		TR_72 = RG_rl_159 ;
	7'h43 :
		TR_72 = RG_rl_159 ;
	7'h44 :
		TR_72 = RG_rl_159 ;
	7'h45 :
		TR_72 = RG_rl_159 ;
	7'h46 :
		TR_72 = RG_rl_159 ;
	7'h47 :
		TR_72 = RG_rl_159 ;
	7'h48 :
		TR_72 = RG_rl_159 ;
	7'h49 :
		TR_72 = RG_rl_159 ;
	7'h4a :
		TR_72 = RG_rl_159 ;
	7'h4b :
		TR_72 = RG_rl_159 ;
	7'h4c :
		TR_72 = RG_rl_159 ;
	7'h4d :
		TR_72 = RG_rl_159 ;
	7'h4e :
		TR_72 = RG_rl_159 ;
	7'h4f :
		TR_72 = RG_rl_159 ;
	7'h50 :
		TR_72 = RG_rl_159 ;
	7'h51 :
		TR_72 = RG_rl_159 ;
	7'h52 :
		TR_72 = RG_rl_159 ;
	7'h53 :
		TR_72 = RG_rl_159 ;
	7'h54 :
		TR_72 = RG_rl_159 ;
	7'h55 :
		TR_72 = RG_rl_159 ;
	7'h56 :
		TR_72 = RG_rl_159 ;
	7'h57 :
		TR_72 = RG_rl_159 ;
	7'h58 :
		TR_72 = RG_rl_159 ;
	7'h59 :
		TR_72 = RG_rl_159 ;
	7'h5a :
		TR_72 = RG_rl_159 ;
	7'h5b :
		TR_72 = RG_rl_159 ;
	7'h5c :
		TR_72 = RG_rl_159 ;
	7'h5d :
		TR_72 = RG_rl_159 ;
	7'h5e :
		TR_72 = RG_rl_159 ;
	7'h5f :
		TR_72 = RG_rl_159 ;
	7'h60 :
		TR_72 = RG_rl_159 ;
	7'h61 :
		TR_72 = RG_rl_159 ;
	7'h62 :
		TR_72 = RG_rl_159 ;
	7'h63 :
		TR_72 = RG_rl_159 ;
	7'h64 :
		TR_72 = RG_rl_159 ;
	7'h65 :
		TR_72 = RG_rl_159 ;
	7'h66 :
		TR_72 = RG_rl_159 ;
	7'h67 :
		TR_72 = RG_rl_159 ;
	7'h68 :
		TR_72 = RG_rl_159 ;
	7'h69 :
		TR_72 = RG_rl_159 ;
	7'h6a :
		TR_72 = RG_rl_159 ;
	7'h6b :
		TR_72 = RG_rl_159 ;
	7'h6c :
		TR_72 = RG_rl_159 ;
	7'h6d :
		TR_72 = RG_rl_159 ;
	7'h6e :
		TR_72 = RG_rl_159 ;
	7'h6f :
		TR_72 = RG_rl_159 ;
	7'h70 :
		TR_72 = RG_rl_159 ;
	7'h71 :
		TR_72 = RG_rl_159 ;
	7'h72 :
		TR_72 = RG_rl_159 ;
	7'h73 :
		TR_72 = RG_rl_159 ;
	7'h74 :
		TR_72 = RG_rl_159 ;
	7'h75 :
		TR_72 = RG_rl_159 ;
	7'h76 :
		TR_72 = RG_rl_159 ;
	7'h77 :
		TR_72 = RG_rl_159 ;
	7'h78 :
		TR_72 = RG_rl_159 ;
	7'h79 :
		TR_72 = RG_rl_159 ;
	7'h7a :
		TR_72 = RG_rl_159 ;
	7'h7b :
		TR_72 = RG_rl_159 ;
	7'h7c :
		TR_72 = RG_rl_159 ;
	7'h7d :
		TR_72 = RG_rl_159 ;
	7'h7e :
		TR_72 = RG_rl_159 ;
	7'h7f :
		TR_72 = RG_rl_159 ;
	default :
		TR_72 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_28 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h01 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h02 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h03 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h04 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h05 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h06 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h07 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h08 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h09 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h0a :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h0b :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h0c :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h0d :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h0e :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h0f :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h10 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h11 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h12 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h13 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h14 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h15 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h16 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h17 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h18 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h19 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h1a :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h1b :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h1c :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h1d :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h1e :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h1f :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h20 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h21 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h22 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h23 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h24 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h25 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h26 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h27 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h28 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h29 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h2a :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h2b :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h2c :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h2d :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h2e :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h2f :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h30 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h31 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h32 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h33 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h34 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h35 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h36 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h37 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h38 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h39 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h3a :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h3b :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h3c :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h3d :
		TR_73 = 9'h000 ;	// line#=../rle.cpp:79
	7'h3e :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h3f :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h40 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h41 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h42 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h43 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h44 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h45 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h46 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h47 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h48 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h49 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h4a :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h4b :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h4c :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h4d :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h4e :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h4f :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h50 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h51 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h52 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h53 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h54 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h55 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h56 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h57 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h58 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h59 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h5a :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h5b :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h5c :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h5d :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h5e :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h5f :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h60 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h61 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h62 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h63 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h64 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h65 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h66 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h67 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h68 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h69 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h6a :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h6b :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h6c :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h6d :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h6e :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h6f :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h70 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h71 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h72 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h73 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h74 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h75 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h76 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h77 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h78 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h79 :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h7a :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h7b :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h7c :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h7d :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h7e :
		TR_73 = RG_quantized_block_rl_28 ;
	7'h7f :
		TR_73 = RG_quantized_block_rl_28 ;
	default :
		TR_73 = 9'hx ;
	endcase
always @ ( RG_rl_160 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_74 = RG_rl_160 ;
	7'h01 :
		TR_74 = RG_rl_160 ;
	7'h02 :
		TR_74 = RG_rl_160 ;
	7'h03 :
		TR_74 = RG_rl_160 ;
	7'h04 :
		TR_74 = RG_rl_160 ;
	7'h05 :
		TR_74 = RG_rl_160 ;
	7'h06 :
		TR_74 = RG_rl_160 ;
	7'h07 :
		TR_74 = RG_rl_160 ;
	7'h08 :
		TR_74 = RG_rl_160 ;
	7'h09 :
		TR_74 = RG_rl_160 ;
	7'h0a :
		TR_74 = RG_rl_160 ;
	7'h0b :
		TR_74 = RG_rl_160 ;
	7'h0c :
		TR_74 = RG_rl_160 ;
	7'h0d :
		TR_74 = RG_rl_160 ;
	7'h0e :
		TR_74 = RG_rl_160 ;
	7'h0f :
		TR_74 = RG_rl_160 ;
	7'h10 :
		TR_74 = RG_rl_160 ;
	7'h11 :
		TR_74 = RG_rl_160 ;
	7'h12 :
		TR_74 = RG_rl_160 ;
	7'h13 :
		TR_74 = RG_rl_160 ;
	7'h14 :
		TR_74 = RG_rl_160 ;
	7'h15 :
		TR_74 = RG_rl_160 ;
	7'h16 :
		TR_74 = RG_rl_160 ;
	7'h17 :
		TR_74 = RG_rl_160 ;
	7'h18 :
		TR_74 = RG_rl_160 ;
	7'h19 :
		TR_74 = RG_rl_160 ;
	7'h1a :
		TR_74 = RG_rl_160 ;
	7'h1b :
		TR_74 = RG_rl_160 ;
	7'h1c :
		TR_74 = RG_rl_160 ;
	7'h1d :
		TR_74 = RG_rl_160 ;
	7'h1e :
		TR_74 = RG_rl_160 ;
	7'h1f :
		TR_74 = RG_rl_160 ;
	7'h20 :
		TR_74 = RG_rl_160 ;
	7'h21 :
		TR_74 = RG_rl_160 ;
	7'h22 :
		TR_74 = RG_rl_160 ;
	7'h23 :
		TR_74 = RG_rl_160 ;
	7'h24 :
		TR_74 = RG_rl_160 ;
	7'h25 :
		TR_74 = RG_rl_160 ;
	7'h26 :
		TR_74 = RG_rl_160 ;
	7'h27 :
		TR_74 = RG_rl_160 ;
	7'h28 :
		TR_74 = RG_rl_160 ;
	7'h29 :
		TR_74 = RG_rl_160 ;
	7'h2a :
		TR_74 = RG_rl_160 ;
	7'h2b :
		TR_74 = RG_rl_160 ;
	7'h2c :
		TR_74 = RG_rl_160 ;
	7'h2d :
		TR_74 = RG_rl_160 ;
	7'h2e :
		TR_74 = RG_rl_160 ;
	7'h2f :
		TR_74 = RG_rl_160 ;
	7'h30 :
		TR_74 = RG_rl_160 ;
	7'h31 :
		TR_74 = RG_rl_160 ;
	7'h32 :
		TR_74 = RG_rl_160 ;
	7'h33 :
		TR_74 = RG_rl_160 ;
	7'h34 :
		TR_74 = RG_rl_160 ;
	7'h35 :
		TR_74 = RG_rl_160 ;
	7'h36 :
		TR_74 = RG_rl_160 ;
	7'h37 :
		TR_74 = RG_rl_160 ;
	7'h38 :
		TR_74 = RG_rl_160 ;
	7'h39 :
		TR_74 = RG_rl_160 ;
	7'h3a :
		TR_74 = RG_rl_160 ;
	7'h3b :
		TR_74 = RG_rl_160 ;
	7'h3c :
		TR_74 = RG_rl_160 ;
	7'h3d :
		TR_74 = RG_rl_160 ;
	7'h3e :
		TR_74 = 9'h000 ;	// line#=../rle.cpp:79
	7'h3f :
		TR_74 = RG_rl_160 ;
	7'h40 :
		TR_74 = RG_rl_160 ;
	7'h41 :
		TR_74 = RG_rl_160 ;
	7'h42 :
		TR_74 = RG_rl_160 ;
	7'h43 :
		TR_74 = RG_rl_160 ;
	7'h44 :
		TR_74 = RG_rl_160 ;
	7'h45 :
		TR_74 = RG_rl_160 ;
	7'h46 :
		TR_74 = RG_rl_160 ;
	7'h47 :
		TR_74 = RG_rl_160 ;
	7'h48 :
		TR_74 = RG_rl_160 ;
	7'h49 :
		TR_74 = RG_rl_160 ;
	7'h4a :
		TR_74 = RG_rl_160 ;
	7'h4b :
		TR_74 = RG_rl_160 ;
	7'h4c :
		TR_74 = RG_rl_160 ;
	7'h4d :
		TR_74 = RG_rl_160 ;
	7'h4e :
		TR_74 = RG_rl_160 ;
	7'h4f :
		TR_74 = RG_rl_160 ;
	7'h50 :
		TR_74 = RG_rl_160 ;
	7'h51 :
		TR_74 = RG_rl_160 ;
	7'h52 :
		TR_74 = RG_rl_160 ;
	7'h53 :
		TR_74 = RG_rl_160 ;
	7'h54 :
		TR_74 = RG_rl_160 ;
	7'h55 :
		TR_74 = RG_rl_160 ;
	7'h56 :
		TR_74 = RG_rl_160 ;
	7'h57 :
		TR_74 = RG_rl_160 ;
	7'h58 :
		TR_74 = RG_rl_160 ;
	7'h59 :
		TR_74 = RG_rl_160 ;
	7'h5a :
		TR_74 = RG_rl_160 ;
	7'h5b :
		TR_74 = RG_rl_160 ;
	7'h5c :
		TR_74 = RG_rl_160 ;
	7'h5d :
		TR_74 = RG_rl_160 ;
	7'h5e :
		TR_74 = RG_rl_160 ;
	7'h5f :
		TR_74 = RG_rl_160 ;
	7'h60 :
		TR_74 = RG_rl_160 ;
	7'h61 :
		TR_74 = RG_rl_160 ;
	7'h62 :
		TR_74 = RG_rl_160 ;
	7'h63 :
		TR_74 = RG_rl_160 ;
	7'h64 :
		TR_74 = RG_rl_160 ;
	7'h65 :
		TR_74 = RG_rl_160 ;
	7'h66 :
		TR_74 = RG_rl_160 ;
	7'h67 :
		TR_74 = RG_rl_160 ;
	7'h68 :
		TR_74 = RG_rl_160 ;
	7'h69 :
		TR_74 = RG_rl_160 ;
	7'h6a :
		TR_74 = RG_rl_160 ;
	7'h6b :
		TR_74 = RG_rl_160 ;
	7'h6c :
		TR_74 = RG_rl_160 ;
	7'h6d :
		TR_74 = RG_rl_160 ;
	7'h6e :
		TR_74 = RG_rl_160 ;
	7'h6f :
		TR_74 = RG_rl_160 ;
	7'h70 :
		TR_74 = RG_rl_160 ;
	7'h71 :
		TR_74 = RG_rl_160 ;
	7'h72 :
		TR_74 = RG_rl_160 ;
	7'h73 :
		TR_74 = RG_rl_160 ;
	7'h74 :
		TR_74 = RG_rl_160 ;
	7'h75 :
		TR_74 = RG_rl_160 ;
	7'h76 :
		TR_74 = RG_rl_160 ;
	7'h77 :
		TR_74 = RG_rl_160 ;
	7'h78 :
		TR_74 = RG_rl_160 ;
	7'h79 :
		TR_74 = RG_rl_160 ;
	7'h7a :
		TR_74 = RG_rl_160 ;
	7'h7b :
		TR_74 = RG_rl_160 ;
	7'h7c :
		TR_74 = RG_rl_160 ;
	7'h7d :
		TR_74 = RG_rl_160 ;
	7'h7e :
		TR_74 = RG_rl_160 ;
	7'h7f :
		TR_74 = RG_rl_160 ;
	default :
		TR_74 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_29 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h01 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h02 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h03 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h04 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h05 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h06 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h07 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h08 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h09 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h0a :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h0b :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h0c :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h0d :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h0e :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h0f :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h10 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h11 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h12 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h13 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h14 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h15 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h16 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h17 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h18 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h19 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h1a :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h1b :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h1c :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h1d :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h1e :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h1f :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h20 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h21 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h22 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h23 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h24 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h25 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h26 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h27 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h28 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h29 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h2a :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h2b :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h2c :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h2d :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h2e :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h2f :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h30 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h31 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h32 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h33 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h34 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h35 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h36 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h37 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h38 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h39 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h3a :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h3b :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h3c :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h3d :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h3e :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h3f :
		TR_75 = 9'h000 ;	// line#=../rle.cpp:79
	7'h40 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h41 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h42 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h43 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h44 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h45 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h46 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h47 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h48 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h49 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h4a :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h4b :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h4c :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h4d :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h4e :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h4f :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h50 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h51 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h52 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h53 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h54 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h55 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h56 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h57 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h58 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h59 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h5a :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h5b :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h5c :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h5d :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h5e :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h5f :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h60 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h61 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h62 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h63 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h64 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h65 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h66 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h67 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h68 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h69 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h6a :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h6b :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h6c :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h6d :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h6e :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h6f :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h70 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h71 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h72 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h73 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h74 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h75 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h76 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h77 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h78 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h79 :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h7a :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h7b :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h7c :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h7d :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h7e :
		TR_75 = RG_quantized_block_rl_29 ;
	7'h7f :
		TR_75 = RG_quantized_block_rl_29 ;
	default :
		TR_75 = 9'hx ;
	endcase
always @ ( RG_rl_161 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_76 = RG_rl_161 ;
	7'h01 :
		TR_76 = RG_rl_161 ;
	7'h02 :
		TR_76 = RG_rl_161 ;
	7'h03 :
		TR_76 = RG_rl_161 ;
	7'h04 :
		TR_76 = RG_rl_161 ;
	7'h05 :
		TR_76 = RG_rl_161 ;
	7'h06 :
		TR_76 = RG_rl_161 ;
	7'h07 :
		TR_76 = RG_rl_161 ;
	7'h08 :
		TR_76 = RG_rl_161 ;
	7'h09 :
		TR_76 = RG_rl_161 ;
	7'h0a :
		TR_76 = RG_rl_161 ;
	7'h0b :
		TR_76 = RG_rl_161 ;
	7'h0c :
		TR_76 = RG_rl_161 ;
	7'h0d :
		TR_76 = RG_rl_161 ;
	7'h0e :
		TR_76 = RG_rl_161 ;
	7'h0f :
		TR_76 = RG_rl_161 ;
	7'h10 :
		TR_76 = RG_rl_161 ;
	7'h11 :
		TR_76 = RG_rl_161 ;
	7'h12 :
		TR_76 = RG_rl_161 ;
	7'h13 :
		TR_76 = RG_rl_161 ;
	7'h14 :
		TR_76 = RG_rl_161 ;
	7'h15 :
		TR_76 = RG_rl_161 ;
	7'h16 :
		TR_76 = RG_rl_161 ;
	7'h17 :
		TR_76 = RG_rl_161 ;
	7'h18 :
		TR_76 = RG_rl_161 ;
	7'h19 :
		TR_76 = RG_rl_161 ;
	7'h1a :
		TR_76 = RG_rl_161 ;
	7'h1b :
		TR_76 = RG_rl_161 ;
	7'h1c :
		TR_76 = RG_rl_161 ;
	7'h1d :
		TR_76 = RG_rl_161 ;
	7'h1e :
		TR_76 = RG_rl_161 ;
	7'h1f :
		TR_76 = RG_rl_161 ;
	7'h20 :
		TR_76 = RG_rl_161 ;
	7'h21 :
		TR_76 = RG_rl_161 ;
	7'h22 :
		TR_76 = RG_rl_161 ;
	7'h23 :
		TR_76 = RG_rl_161 ;
	7'h24 :
		TR_76 = RG_rl_161 ;
	7'h25 :
		TR_76 = RG_rl_161 ;
	7'h26 :
		TR_76 = RG_rl_161 ;
	7'h27 :
		TR_76 = RG_rl_161 ;
	7'h28 :
		TR_76 = RG_rl_161 ;
	7'h29 :
		TR_76 = RG_rl_161 ;
	7'h2a :
		TR_76 = RG_rl_161 ;
	7'h2b :
		TR_76 = RG_rl_161 ;
	7'h2c :
		TR_76 = RG_rl_161 ;
	7'h2d :
		TR_76 = RG_rl_161 ;
	7'h2e :
		TR_76 = RG_rl_161 ;
	7'h2f :
		TR_76 = RG_rl_161 ;
	7'h30 :
		TR_76 = RG_rl_161 ;
	7'h31 :
		TR_76 = RG_rl_161 ;
	7'h32 :
		TR_76 = RG_rl_161 ;
	7'h33 :
		TR_76 = RG_rl_161 ;
	7'h34 :
		TR_76 = RG_rl_161 ;
	7'h35 :
		TR_76 = RG_rl_161 ;
	7'h36 :
		TR_76 = RG_rl_161 ;
	7'h37 :
		TR_76 = RG_rl_161 ;
	7'h38 :
		TR_76 = RG_rl_161 ;
	7'h39 :
		TR_76 = RG_rl_161 ;
	7'h3a :
		TR_76 = RG_rl_161 ;
	7'h3b :
		TR_76 = RG_rl_161 ;
	7'h3c :
		TR_76 = RG_rl_161 ;
	7'h3d :
		TR_76 = RG_rl_161 ;
	7'h3e :
		TR_76 = RG_rl_161 ;
	7'h3f :
		TR_76 = RG_rl_161 ;
	7'h40 :
		TR_76 = 9'h000 ;	// line#=../rle.cpp:79
	7'h41 :
		TR_76 = RG_rl_161 ;
	7'h42 :
		TR_76 = RG_rl_161 ;
	7'h43 :
		TR_76 = RG_rl_161 ;
	7'h44 :
		TR_76 = RG_rl_161 ;
	7'h45 :
		TR_76 = RG_rl_161 ;
	7'h46 :
		TR_76 = RG_rl_161 ;
	7'h47 :
		TR_76 = RG_rl_161 ;
	7'h48 :
		TR_76 = RG_rl_161 ;
	7'h49 :
		TR_76 = RG_rl_161 ;
	7'h4a :
		TR_76 = RG_rl_161 ;
	7'h4b :
		TR_76 = RG_rl_161 ;
	7'h4c :
		TR_76 = RG_rl_161 ;
	7'h4d :
		TR_76 = RG_rl_161 ;
	7'h4e :
		TR_76 = RG_rl_161 ;
	7'h4f :
		TR_76 = RG_rl_161 ;
	7'h50 :
		TR_76 = RG_rl_161 ;
	7'h51 :
		TR_76 = RG_rl_161 ;
	7'h52 :
		TR_76 = RG_rl_161 ;
	7'h53 :
		TR_76 = RG_rl_161 ;
	7'h54 :
		TR_76 = RG_rl_161 ;
	7'h55 :
		TR_76 = RG_rl_161 ;
	7'h56 :
		TR_76 = RG_rl_161 ;
	7'h57 :
		TR_76 = RG_rl_161 ;
	7'h58 :
		TR_76 = RG_rl_161 ;
	7'h59 :
		TR_76 = RG_rl_161 ;
	7'h5a :
		TR_76 = RG_rl_161 ;
	7'h5b :
		TR_76 = RG_rl_161 ;
	7'h5c :
		TR_76 = RG_rl_161 ;
	7'h5d :
		TR_76 = RG_rl_161 ;
	7'h5e :
		TR_76 = RG_rl_161 ;
	7'h5f :
		TR_76 = RG_rl_161 ;
	7'h60 :
		TR_76 = RG_rl_161 ;
	7'h61 :
		TR_76 = RG_rl_161 ;
	7'h62 :
		TR_76 = RG_rl_161 ;
	7'h63 :
		TR_76 = RG_rl_161 ;
	7'h64 :
		TR_76 = RG_rl_161 ;
	7'h65 :
		TR_76 = RG_rl_161 ;
	7'h66 :
		TR_76 = RG_rl_161 ;
	7'h67 :
		TR_76 = RG_rl_161 ;
	7'h68 :
		TR_76 = RG_rl_161 ;
	7'h69 :
		TR_76 = RG_rl_161 ;
	7'h6a :
		TR_76 = RG_rl_161 ;
	7'h6b :
		TR_76 = RG_rl_161 ;
	7'h6c :
		TR_76 = RG_rl_161 ;
	7'h6d :
		TR_76 = RG_rl_161 ;
	7'h6e :
		TR_76 = RG_rl_161 ;
	7'h6f :
		TR_76 = RG_rl_161 ;
	7'h70 :
		TR_76 = RG_rl_161 ;
	7'h71 :
		TR_76 = RG_rl_161 ;
	7'h72 :
		TR_76 = RG_rl_161 ;
	7'h73 :
		TR_76 = RG_rl_161 ;
	7'h74 :
		TR_76 = RG_rl_161 ;
	7'h75 :
		TR_76 = RG_rl_161 ;
	7'h76 :
		TR_76 = RG_rl_161 ;
	7'h77 :
		TR_76 = RG_rl_161 ;
	7'h78 :
		TR_76 = RG_rl_161 ;
	7'h79 :
		TR_76 = RG_rl_161 ;
	7'h7a :
		TR_76 = RG_rl_161 ;
	7'h7b :
		TR_76 = RG_rl_161 ;
	7'h7c :
		TR_76 = RG_rl_161 ;
	7'h7d :
		TR_76 = RG_rl_161 ;
	7'h7e :
		TR_76 = RG_rl_161 ;
	7'h7f :
		TR_76 = RG_rl_161 ;
	default :
		TR_76 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_30 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h01 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h02 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h03 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h04 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h05 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h06 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h07 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h08 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h09 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h0a :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h0b :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h0c :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h0d :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h0e :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h0f :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h10 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h11 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h12 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h13 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h14 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h15 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h16 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h17 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h18 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h19 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h1a :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h1b :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h1c :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h1d :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h1e :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h1f :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h20 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h21 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h22 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h23 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h24 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h25 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h26 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h27 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h28 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h29 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h2a :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h2b :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h2c :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h2d :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h2e :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h2f :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h30 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h31 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h32 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h33 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h34 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h35 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h36 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h37 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h38 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h39 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h3a :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h3b :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h3c :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h3d :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h3e :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h3f :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h40 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h41 :
		TR_77 = 9'h000 ;	// line#=../rle.cpp:79
	7'h42 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h43 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h44 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h45 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h46 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h47 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h48 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h49 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h4a :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h4b :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h4c :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h4d :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h4e :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h4f :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h50 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h51 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h52 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h53 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h54 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h55 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h56 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h57 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h58 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h59 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h5a :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h5b :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h5c :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h5d :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h5e :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h5f :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h60 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h61 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h62 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h63 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h64 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h65 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h66 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h67 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h68 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h69 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h6a :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h6b :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h6c :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h6d :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h6e :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h6f :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h70 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h71 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h72 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h73 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h74 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h75 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h76 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h77 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h78 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h79 :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h7a :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h7b :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h7c :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h7d :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h7e :
		TR_77 = RG_quantized_block_rl_30 ;
	7'h7f :
		TR_77 = RG_quantized_block_rl_30 ;
	default :
		TR_77 = 9'hx ;
	endcase
always @ ( RG_rl_162 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_78 = RG_rl_162 ;
	7'h01 :
		TR_78 = RG_rl_162 ;
	7'h02 :
		TR_78 = RG_rl_162 ;
	7'h03 :
		TR_78 = RG_rl_162 ;
	7'h04 :
		TR_78 = RG_rl_162 ;
	7'h05 :
		TR_78 = RG_rl_162 ;
	7'h06 :
		TR_78 = RG_rl_162 ;
	7'h07 :
		TR_78 = RG_rl_162 ;
	7'h08 :
		TR_78 = RG_rl_162 ;
	7'h09 :
		TR_78 = RG_rl_162 ;
	7'h0a :
		TR_78 = RG_rl_162 ;
	7'h0b :
		TR_78 = RG_rl_162 ;
	7'h0c :
		TR_78 = RG_rl_162 ;
	7'h0d :
		TR_78 = RG_rl_162 ;
	7'h0e :
		TR_78 = RG_rl_162 ;
	7'h0f :
		TR_78 = RG_rl_162 ;
	7'h10 :
		TR_78 = RG_rl_162 ;
	7'h11 :
		TR_78 = RG_rl_162 ;
	7'h12 :
		TR_78 = RG_rl_162 ;
	7'h13 :
		TR_78 = RG_rl_162 ;
	7'h14 :
		TR_78 = RG_rl_162 ;
	7'h15 :
		TR_78 = RG_rl_162 ;
	7'h16 :
		TR_78 = RG_rl_162 ;
	7'h17 :
		TR_78 = RG_rl_162 ;
	7'h18 :
		TR_78 = RG_rl_162 ;
	7'h19 :
		TR_78 = RG_rl_162 ;
	7'h1a :
		TR_78 = RG_rl_162 ;
	7'h1b :
		TR_78 = RG_rl_162 ;
	7'h1c :
		TR_78 = RG_rl_162 ;
	7'h1d :
		TR_78 = RG_rl_162 ;
	7'h1e :
		TR_78 = RG_rl_162 ;
	7'h1f :
		TR_78 = RG_rl_162 ;
	7'h20 :
		TR_78 = RG_rl_162 ;
	7'h21 :
		TR_78 = RG_rl_162 ;
	7'h22 :
		TR_78 = RG_rl_162 ;
	7'h23 :
		TR_78 = RG_rl_162 ;
	7'h24 :
		TR_78 = RG_rl_162 ;
	7'h25 :
		TR_78 = RG_rl_162 ;
	7'h26 :
		TR_78 = RG_rl_162 ;
	7'h27 :
		TR_78 = RG_rl_162 ;
	7'h28 :
		TR_78 = RG_rl_162 ;
	7'h29 :
		TR_78 = RG_rl_162 ;
	7'h2a :
		TR_78 = RG_rl_162 ;
	7'h2b :
		TR_78 = RG_rl_162 ;
	7'h2c :
		TR_78 = RG_rl_162 ;
	7'h2d :
		TR_78 = RG_rl_162 ;
	7'h2e :
		TR_78 = RG_rl_162 ;
	7'h2f :
		TR_78 = RG_rl_162 ;
	7'h30 :
		TR_78 = RG_rl_162 ;
	7'h31 :
		TR_78 = RG_rl_162 ;
	7'h32 :
		TR_78 = RG_rl_162 ;
	7'h33 :
		TR_78 = RG_rl_162 ;
	7'h34 :
		TR_78 = RG_rl_162 ;
	7'h35 :
		TR_78 = RG_rl_162 ;
	7'h36 :
		TR_78 = RG_rl_162 ;
	7'h37 :
		TR_78 = RG_rl_162 ;
	7'h38 :
		TR_78 = RG_rl_162 ;
	7'h39 :
		TR_78 = RG_rl_162 ;
	7'h3a :
		TR_78 = RG_rl_162 ;
	7'h3b :
		TR_78 = RG_rl_162 ;
	7'h3c :
		TR_78 = RG_rl_162 ;
	7'h3d :
		TR_78 = RG_rl_162 ;
	7'h3e :
		TR_78 = RG_rl_162 ;
	7'h3f :
		TR_78 = RG_rl_162 ;
	7'h40 :
		TR_78 = RG_rl_162 ;
	7'h41 :
		TR_78 = RG_rl_162 ;
	7'h42 :
		TR_78 = 9'h000 ;	// line#=../rle.cpp:79
	7'h43 :
		TR_78 = RG_rl_162 ;
	7'h44 :
		TR_78 = RG_rl_162 ;
	7'h45 :
		TR_78 = RG_rl_162 ;
	7'h46 :
		TR_78 = RG_rl_162 ;
	7'h47 :
		TR_78 = RG_rl_162 ;
	7'h48 :
		TR_78 = RG_rl_162 ;
	7'h49 :
		TR_78 = RG_rl_162 ;
	7'h4a :
		TR_78 = RG_rl_162 ;
	7'h4b :
		TR_78 = RG_rl_162 ;
	7'h4c :
		TR_78 = RG_rl_162 ;
	7'h4d :
		TR_78 = RG_rl_162 ;
	7'h4e :
		TR_78 = RG_rl_162 ;
	7'h4f :
		TR_78 = RG_rl_162 ;
	7'h50 :
		TR_78 = RG_rl_162 ;
	7'h51 :
		TR_78 = RG_rl_162 ;
	7'h52 :
		TR_78 = RG_rl_162 ;
	7'h53 :
		TR_78 = RG_rl_162 ;
	7'h54 :
		TR_78 = RG_rl_162 ;
	7'h55 :
		TR_78 = RG_rl_162 ;
	7'h56 :
		TR_78 = RG_rl_162 ;
	7'h57 :
		TR_78 = RG_rl_162 ;
	7'h58 :
		TR_78 = RG_rl_162 ;
	7'h59 :
		TR_78 = RG_rl_162 ;
	7'h5a :
		TR_78 = RG_rl_162 ;
	7'h5b :
		TR_78 = RG_rl_162 ;
	7'h5c :
		TR_78 = RG_rl_162 ;
	7'h5d :
		TR_78 = RG_rl_162 ;
	7'h5e :
		TR_78 = RG_rl_162 ;
	7'h5f :
		TR_78 = RG_rl_162 ;
	7'h60 :
		TR_78 = RG_rl_162 ;
	7'h61 :
		TR_78 = RG_rl_162 ;
	7'h62 :
		TR_78 = RG_rl_162 ;
	7'h63 :
		TR_78 = RG_rl_162 ;
	7'h64 :
		TR_78 = RG_rl_162 ;
	7'h65 :
		TR_78 = RG_rl_162 ;
	7'h66 :
		TR_78 = RG_rl_162 ;
	7'h67 :
		TR_78 = RG_rl_162 ;
	7'h68 :
		TR_78 = RG_rl_162 ;
	7'h69 :
		TR_78 = RG_rl_162 ;
	7'h6a :
		TR_78 = RG_rl_162 ;
	7'h6b :
		TR_78 = RG_rl_162 ;
	7'h6c :
		TR_78 = RG_rl_162 ;
	7'h6d :
		TR_78 = RG_rl_162 ;
	7'h6e :
		TR_78 = RG_rl_162 ;
	7'h6f :
		TR_78 = RG_rl_162 ;
	7'h70 :
		TR_78 = RG_rl_162 ;
	7'h71 :
		TR_78 = RG_rl_162 ;
	7'h72 :
		TR_78 = RG_rl_162 ;
	7'h73 :
		TR_78 = RG_rl_162 ;
	7'h74 :
		TR_78 = RG_rl_162 ;
	7'h75 :
		TR_78 = RG_rl_162 ;
	7'h76 :
		TR_78 = RG_rl_162 ;
	7'h77 :
		TR_78 = RG_rl_162 ;
	7'h78 :
		TR_78 = RG_rl_162 ;
	7'h79 :
		TR_78 = RG_rl_162 ;
	7'h7a :
		TR_78 = RG_rl_162 ;
	7'h7b :
		TR_78 = RG_rl_162 ;
	7'h7c :
		TR_78 = RG_rl_162 ;
	7'h7d :
		TR_78 = RG_rl_162 ;
	7'h7e :
		TR_78 = RG_rl_162 ;
	7'h7f :
		TR_78 = RG_rl_162 ;
	default :
		TR_78 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_31 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h01 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h02 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h03 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h04 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h05 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h06 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h07 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h08 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h09 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h0a :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h0b :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h0c :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h0d :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h0e :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h0f :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h10 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h11 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h12 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h13 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h14 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h15 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h16 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h17 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h18 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h19 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h1a :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h1b :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h1c :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h1d :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h1e :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h1f :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h20 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h21 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h22 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h23 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h24 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h25 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h26 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h27 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h28 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h29 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h2a :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h2b :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h2c :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h2d :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h2e :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h2f :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h30 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h31 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h32 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h33 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h34 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h35 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h36 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h37 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h38 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h39 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h3a :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h3b :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h3c :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h3d :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h3e :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h3f :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h40 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h41 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h42 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h43 :
		TR_79 = 9'h000 ;	// line#=../rle.cpp:79
	7'h44 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h45 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h46 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h47 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h48 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h49 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h4a :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h4b :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h4c :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h4d :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h4e :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h4f :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h50 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h51 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h52 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h53 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h54 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h55 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h56 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h57 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h58 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h59 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h5a :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h5b :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h5c :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h5d :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h5e :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h5f :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h60 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h61 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h62 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h63 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h64 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h65 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h66 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h67 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h68 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h69 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h6a :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h6b :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h6c :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h6d :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h6e :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h6f :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h70 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h71 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h72 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h73 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h74 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h75 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h76 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h77 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h78 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h79 :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h7a :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h7b :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h7c :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h7d :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h7e :
		TR_79 = RG_quantized_block_rl_31 ;
	7'h7f :
		TR_79 = RG_quantized_block_rl_31 ;
	default :
		TR_79 = 9'hx ;
	endcase
always @ ( RG_rl_163 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_80 = RG_rl_163 ;
	7'h01 :
		TR_80 = RG_rl_163 ;
	7'h02 :
		TR_80 = RG_rl_163 ;
	7'h03 :
		TR_80 = RG_rl_163 ;
	7'h04 :
		TR_80 = RG_rl_163 ;
	7'h05 :
		TR_80 = RG_rl_163 ;
	7'h06 :
		TR_80 = RG_rl_163 ;
	7'h07 :
		TR_80 = RG_rl_163 ;
	7'h08 :
		TR_80 = RG_rl_163 ;
	7'h09 :
		TR_80 = RG_rl_163 ;
	7'h0a :
		TR_80 = RG_rl_163 ;
	7'h0b :
		TR_80 = RG_rl_163 ;
	7'h0c :
		TR_80 = RG_rl_163 ;
	7'h0d :
		TR_80 = RG_rl_163 ;
	7'h0e :
		TR_80 = RG_rl_163 ;
	7'h0f :
		TR_80 = RG_rl_163 ;
	7'h10 :
		TR_80 = RG_rl_163 ;
	7'h11 :
		TR_80 = RG_rl_163 ;
	7'h12 :
		TR_80 = RG_rl_163 ;
	7'h13 :
		TR_80 = RG_rl_163 ;
	7'h14 :
		TR_80 = RG_rl_163 ;
	7'h15 :
		TR_80 = RG_rl_163 ;
	7'h16 :
		TR_80 = RG_rl_163 ;
	7'h17 :
		TR_80 = RG_rl_163 ;
	7'h18 :
		TR_80 = RG_rl_163 ;
	7'h19 :
		TR_80 = RG_rl_163 ;
	7'h1a :
		TR_80 = RG_rl_163 ;
	7'h1b :
		TR_80 = RG_rl_163 ;
	7'h1c :
		TR_80 = RG_rl_163 ;
	7'h1d :
		TR_80 = RG_rl_163 ;
	7'h1e :
		TR_80 = RG_rl_163 ;
	7'h1f :
		TR_80 = RG_rl_163 ;
	7'h20 :
		TR_80 = RG_rl_163 ;
	7'h21 :
		TR_80 = RG_rl_163 ;
	7'h22 :
		TR_80 = RG_rl_163 ;
	7'h23 :
		TR_80 = RG_rl_163 ;
	7'h24 :
		TR_80 = RG_rl_163 ;
	7'h25 :
		TR_80 = RG_rl_163 ;
	7'h26 :
		TR_80 = RG_rl_163 ;
	7'h27 :
		TR_80 = RG_rl_163 ;
	7'h28 :
		TR_80 = RG_rl_163 ;
	7'h29 :
		TR_80 = RG_rl_163 ;
	7'h2a :
		TR_80 = RG_rl_163 ;
	7'h2b :
		TR_80 = RG_rl_163 ;
	7'h2c :
		TR_80 = RG_rl_163 ;
	7'h2d :
		TR_80 = RG_rl_163 ;
	7'h2e :
		TR_80 = RG_rl_163 ;
	7'h2f :
		TR_80 = RG_rl_163 ;
	7'h30 :
		TR_80 = RG_rl_163 ;
	7'h31 :
		TR_80 = RG_rl_163 ;
	7'h32 :
		TR_80 = RG_rl_163 ;
	7'h33 :
		TR_80 = RG_rl_163 ;
	7'h34 :
		TR_80 = RG_rl_163 ;
	7'h35 :
		TR_80 = RG_rl_163 ;
	7'h36 :
		TR_80 = RG_rl_163 ;
	7'h37 :
		TR_80 = RG_rl_163 ;
	7'h38 :
		TR_80 = RG_rl_163 ;
	7'h39 :
		TR_80 = RG_rl_163 ;
	7'h3a :
		TR_80 = RG_rl_163 ;
	7'h3b :
		TR_80 = RG_rl_163 ;
	7'h3c :
		TR_80 = RG_rl_163 ;
	7'h3d :
		TR_80 = RG_rl_163 ;
	7'h3e :
		TR_80 = RG_rl_163 ;
	7'h3f :
		TR_80 = RG_rl_163 ;
	7'h40 :
		TR_80 = RG_rl_163 ;
	7'h41 :
		TR_80 = RG_rl_163 ;
	7'h42 :
		TR_80 = RG_rl_163 ;
	7'h43 :
		TR_80 = RG_rl_163 ;
	7'h44 :
		TR_80 = 9'h000 ;	// line#=../rle.cpp:79
	7'h45 :
		TR_80 = RG_rl_163 ;
	7'h46 :
		TR_80 = RG_rl_163 ;
	7'h47 :
		TR_80 = RG_rl_163 ;
	7'h48 :
		TR_80 = RG_rl_163 ;
	7'h49 :
		TR_80 = RG_rl_163 ;
	7'h4a :
		TR_80 = RG_rl_163 ;
	7'h4b :
		TR_80 = RG_rl_163 ;
	7'h4c :
		TR_80 = RG_rl_163 ;
	7'h4d :
		TR_80 = RG_rl_163 ;
	7'h4e :
		TR_80 = RG_rl_163 ;
	7'h4f :
		TR_80 = RG_rl_163 ;
	7'h50 :
		TR_80 = RG_rl_163 ;
	7'h51 :
		TR_80 = RG_rl_163 ;
	7'h52 :
		TR_80 = RG_rl_163 ;
	7'h53 :
		TR_80 = RG_rl_163 ;
	7'h54 :
		TR_80 = RG_rl_163 ;
	7'h55 :
		TR_80 = RG_rl_163 ;
	7'h56 :
		TR_80 = RG_rl_163 ;
	7'h57 :
		TR_80 = RG_rl_163 ;
	7'h58 :
		TR_80 = RG_rl_163 ;
	7'h59 :
		TR_80 = RG_rl_163 ;
	7'h5a :
		TR_80 = RG_rl_163 ;
	7'h5b :
		TR_80 = RG_rl_163 ;
	7'h5c :
		TR_80 = RG_rl_163 ;
	7'h5d :
		TR_80 = RG_rl_163 ;
	7'h5e :
		TR_80 = RG_rl_163 ;
	7'h5f :
		TR_80 = RG_rl_163 ;
	7'h60 :
		TR_80 = RG_rl_163 ;
	7'h61 :
		TR_80 = RG_rl_163 ;
	7'h62 :
		TR_80 = RG_rl_163 ;
	7'h63 :
		TR_80 = RG_rl_163 ;
	7'h64 :
		TR_80 = RG_rl_163 ;
	7'h65 :
		TR_80 = RG_rl_163 ;
	7'h66 :
		TR_80 = RG_rl_163 ;
	7'h67 :
		TR_80 = RG_rl_163 ;
	7'h68 :
		TR_80 = RG_rl_163 ;
	7'h69 :
		TR_80 = RG_rl_163 ;
	7'h6a :
		TR_80 = RG_rl_163 ;
	7'h6b :
		TR_80 = RG_rl_163 ;
	7'h6c :
		TR_80 = RG_rl_163 ;
	7'h6d :
		TR_80 = RG_rl_163 ;
	7'h6e :
		TR_80 = RG_rl_163 ;
	7'h6f :
		TR_80 = RG_rl_163 ;
	7'h70 :
		TR_80 = RG_rl_163 ;
	7'h71 :
		TR_80 = RG_rl_163 ;
	7'h72 :
		TR_80 = RG_rl_163 ;
	7'h73 :
		TR_80 = RG_rl_163 ;
	7'h74 :
		TR_80 = RG_rl_163 ;
	7'h75 :
		TR_80 = RG_rl_163 ;
	7'h76 :
		TR_80 = RG_rl_163 ;
	7'h77 :
		TR_80 = RG_rl_163 ;
	7'h78 :
		TR_80 = RG_rl_163 ;
	7'h79 :
		TR_80 = RG_rl_163 ;
	7'h7a :
		TR_80 = RG_rl_163 ;
	7'h7b :
		TR_80 = RG_rl_163 ;
	7'h7c :
		TR_80 = RG_rl_163 ;
	7'h7d :
		TR_80 = RG_rl_163 ;
	7'h7e :
		TR_80 = RG_rl_163 ;
	7'h7f :
		TR_80 = RG_rl_163 ;
	default :
		TR_80 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_32 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h01 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h02 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h03 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h04 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h05 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h06 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h07 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h08 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h09 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h0a :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h0b :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h0c :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h0d :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h0e :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h0f :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h10 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h11 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h12 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h13 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h14 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h15 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h16 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h17 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h18 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h19 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h1a :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h1b :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h1c :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h1d :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h1e :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h1f :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h20 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h21 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h22 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h23 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h24 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h25 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h26 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h27 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h28 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h29 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h2a :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h2b :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h2c :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h2d :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h2e :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h2f :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h30 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h31 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h32 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h33 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h34 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h35 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h36 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h37 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h38 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h39 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h3a :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h3b :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h3c :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h3d :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h3e :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h3f :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h40 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h41 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h42 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h43 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h44 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h45 :
		TR_81 = 9'h000 ;	// line#=../rle.cpp:79
	7'h46 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h47 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h48 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h49 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h4a :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h4b :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h4c :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h4d :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h4e :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h4f :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h50 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h51 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h52 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h53 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h54 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h55 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h56 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h57 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h58 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h59 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h5a :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h5b :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h5c :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h5d :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h5e :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h5f :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h60 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h61 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h62 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h63 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h64 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h65 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h66 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h67 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h68 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h69 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h6a :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h6b :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h6c :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h6d :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h6e :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h6f :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h70 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h71 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h72 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h73 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h74 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h75 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h76 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h77 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h78 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h79 :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h7a :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h7b :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h7c :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h7d :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h7e :
		TR_81 = RG_quantized_block_rl_32 ;
	7'h7f :
		TR_81 = RG_quantized_block_rl_32 ;
	default :
		TR_81 = 9'hx ;
	endcase
always @ ( RG_rl_164 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_82 = RG_rl_164 ;
	7'h01 :
		TR_82 = RG_rl_164 ;
	7'h02 :
		TR_82 = RG_rl_164 ;
	7'h03 :
		TR_82 = RG_rl_164 ;
	7'h04 :
		TR_82 = RG_rl_164 ;
	7'h05 :
		TR_82 = RG_rl_164 ;
	7'h06 :
		TR_82 = RG_rl_164 ;
	7'h07 :
		TR_82 = RG_rl_164 ;
	7'h08 :
		TR_82 = RG_rl_164 ;
	7'h09 :
		TR_82 = RG_rl_164 ;
	7'h0a :
		TR_82 = RG_rl_164 ;
	7'h0b :
		TR_82 = RG_rl_164 ;
	7'h0c :
		TR_82 = RG_rl_164 ;
	7'h0d :
		TR_82 = RG_rl_164 ;
	7'h0e :
		TR_82 = RG_rl_164 ;
	7'h0f :
		TR_82 = RG_rl_164 ;
	7'h10 :
		TR_82 = RG_rl_164 ;
	7'h11 :
		TR_82 = RG_rl_164 ;
	7'h12 :
		TR_82 = RG_rl_164 ;
	7'h13 :
		TR_82 = RG_rl_164 ;
	7'h14 :
		TR_82 = RG_rl_164 ;
	7'h15 :
		TR_82 = RG_rl_164 ;
	7'h16 :
		TR_82 = RG_rl_164 ;
	7'h17 :
		TR_82 = RG_rl_164 ;
	7'h18 :
		TR_82 = RG_rl_164 ;
	7'h19 :
		TR_82 = RG_rl_164 ;
	7'h1a :
		TR_82 = RG_rl_164 ;
	7'h1b :
		TR_82 = RG_rl_164 ;
	7'h1c :
		TR_82 = RG_rl_164 ;
	7'h1d :
		TR_82 = RG_rl_164 ;
	7'h1e :
		TR_82 = RG_rl_164 ;
	7'h1f :
		TR_82 = RG_rl_164 ;
	7'h20 :
		TR_82 = RG_rl_164 ;
	7'h21 :
		TR_82 = RG_rl_164 ;
	7'h22 :
		TR_82 = RG_rl_164 ;
	7'h23 :
		TR_82 = RG_rl_164 ;
	7'h24 :
		TR_82 = RG_rl_164 ;
	7'h25 :
		TR_82 = RG_rl_164 ;
	7'h26 :
		TR_82 = RG_rl_164 ;
	7'h27 :
		TR_82 = RG_rl_164 ;
	7'h28 :
		TR_82 = RG_rl_164 ;
	7'h29 :
		TR_82 = RG_rl_164 ;
	7'h2a :
		TR_82 = RG_rl_164 ;
	7'h2b :
		TR_82 = RG_rl_164 ;
	7'h2c :
		TR_82 = RG_rl_164 ;
	7'h2d :
		TR_82 = RG_rl_164 ;
	7'h2e :
		TR_82 = RG_rl_164 ;
	7'h2f :
		TR_82 = RG_rl_164 ;
	7'h30 :
		TR_82 = RG_rl_164 ;
	7'h31 :
		TR_82 = RG_rl_164 ;
	7'h32 :
		TR_82 = RG_rl_164 ;
	7'h33 :
		TR_82 = RG_rl_164 ;
	7'h34 :
		TR_82 = RG_rl_164 ;
	7'h35 :
		TR_82 = RG_rl_164 ;
	7'h36 :
		TR_82 = RG_rl_164 ;
	7'h37 :
		TR_82 = RG_rl_164 ;
	7'h38 :
		TR_82 = RG_rl_164 ;
	7'h39 :
		TR_82 = RG_rl_164 ;
	7'h3a :
		TR_82 = RG_rl_164 ;
	7'h3b :
		TR_82 = RG_rl_164 ;
	7'h3c :
		TR_82 = RG_rl_164 ;
	7'h3d :
		TR_82 = RG_rl_164 ;
	7'h3e :
		TR_82 = RG_rl_164 ;
	7'h3f :
		TR_82 = RG_rl_164 ;
	7'h40 :
		TR_82 = RG_rl_164 ;
	7'h41 :
		TR_82 = RG_rl_164 ;
	7'h42 :
		TR_82 = RG_rl_164 ;
	7'h43 :
		TR_82 = RG_rl_164 ;
	7'h44 :
		TR_82 = RG_rl_164 ;
	7'h45 :
		TR_82 = RG_rl_164 ;
	7'h46 :
		TR_82 = 9'h000 ;	// line#=../rle.cpp:79
	7'h47 :
		TR_82 = RG_rl_164 ;
	7'h48 :
		TR_82 = RG_rl_164 ;
	7'h49 :
		TR_82 = RG_rl_164 ;
	7'h4a :
		TR_82 = RG_rl_164 ;
	7'h4b :
		TR_82 = RG_rl_164 ;
	7'h4c :
		TR_82 = RG_rl_164 ;
	7'h4d :
		TR_82 = RG_rl_164 ;
	7'h4e :
		TR_82 = RG_rl_164 ;
	7'h4f :
		TR_82 = RG_rl_164 ;
	7'h50 :
		TR_82 = RG_rl_164 ;
	7'h51 :
		TR_82 = RG_rl_164 ;
	7'h52 :
		TR_82 = RG_rl_164 ;
	7'h53 :
		TR_82 = RG_rl_164 ;
	7'h54 :
		TR_82 = RG_rl_164 ;
	7'h55 :
		TR_82 = RG_rl_164 ;
	7'h56 :
		TR_82 = RG_rl_164 ;
	7'h57 :
		TR_82 = RG_rl_164 ;
	7'h58 :
		TR_82 = RG_rl_164 ;
	7'h59 :
		TR_82 = RG_rl_164 ;
	7'h5a :
		TR_82 = RG_rl_164 ;
	7'h5b :
		TR_82 = RG_rl_164 ;
	7'h5c :
		TR_82 = RG_rl_164 ;
	7'h5d :
		TR_82 = RG_rl_164 ;
	7'h5e :
		TR_82 = RG_rl_164 ;
	7'h5f :
		TR_82 = RG_rl_164 ;
	7'h60 :
		TR_82 = RG_rl_164 ;
	7'h61 :
		TR_82 = RG_rl_164 ;
	7'h62 :
		TR_82 = RG_rl_164 ;
	7'h63 :
		TR_82 = RG_rl_164 ;
	7'h64 :
		TR_82 = RG_rl_164 ;
	7'h65 :
		TR_82 = RG_rl_164 ;
	7'h66 :
		TR_82 = RG_rl_164 ;
	7'h67 :
		TR_82 = RG_rl_164 ;
	7'h68 :
		TR_82 = RG_rl_164 ;
	7'h69 :
		TR_82 = RG_rl_164 ;
	7'h6a :
		TR_82 = RG_rl_164 ;
	7'h6b :
		TR_82 = RG_rl_164 ;
	7'h6c :
		TR_82 = RG_rl_164 ;
	7'h6d :
		TR_82 = RG_rl_164 ;
	7'h6e :
		TR_82 = RG_rl_164 ;
	7'h6f :
		TR_82 = RG_rl_164 ;
	7'h70 :
		TR_82 = RG_rl_164 ;
	7'h71 :
		TR_82 = RG_rl_164 ;
	7'h72 :
		TR_82 = RG_rl_164 ;
	7'h73 :
		TR_82 = RG_rl_164 ;
	7'h74 :
		TR_82 = RG_rl_164 ;
	7'h75 :
		TR_82 = RG_rl_164 ;
	7'h76 :
		TR_82 = RG_rl_164 ;
	7'h77 :
		TR_82 = RG_rl_164 ;
	7'h78 :
		TR_82 = RG_rl_164 ;
	7'h79 :
		TR_82 = RG_rl_164 ;
	7'h7a :
		TR_82 = RG_rl_164 ;
	7'h7b :
		TR_82 = RG_rl_164 ;
	7'h7c :
		TR_82 = RG_rl_164 ;
	7'h7d :
		TR_82 = RG_rl_164 ;
	7'h7e :
		TR_82 = RG_rl_164 ;
	7'h7f :
		TR_82 = RG_rl_164 ;
	default :
		TR_82 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_33 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h01 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h02 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h03 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h04 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h05 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h06 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h07 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h08 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h09 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h0a :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h0b :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h0c :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h0d :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h0e :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h0f :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h10 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h11 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h12 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h13 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h14 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h15 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h16 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h17 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h18 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h19 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h1a :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h1b :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h1c :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h1d :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h1e :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h1f :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h20 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h21 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h22 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h23 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h24 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h25 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h26 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h27 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h28 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h29 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h2a :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h2b :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h2c :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h2d :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h2e :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h2f :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h30 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h31 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h32 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h33 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h34 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h35 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h36 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h37 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h38 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h39 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h3a :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h3b :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h3c :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h3d :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h3e :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h3f :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h40 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h41 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h42 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h43 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h44 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h45 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h46 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h47 :
		TR_83 = 9'h000 ;	// line#=../rle.cpp:79
	7'h48 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h49 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h4a :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h4b :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h4c :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h4d :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h4e :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h4f :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h50 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h51 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h52 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h53 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h54 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h55 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h56 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h57 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h58 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h59 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h5a :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h5b :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h5c :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h5d :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h5e :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h5f :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h60 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h61 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h62 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h63 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h64 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h65 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h66 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h67 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h68 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h69 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h6a :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h6b :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h6c :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h6d :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h6e :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h6f :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h70 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h71 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h72 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h73 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h74 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h75 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h76 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h77 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h78 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h79 :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h7a :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h7b :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h7c :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h7d :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h7e :
		TR_83 = RG_quantized_block_rl_33 ;
	7'h7f :
		TR_83 = RG_quantized_block_rl_33 ;
	default :
		TR_83 = 9'hx ;
	endcase
always @ ( RG_rl_165 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_84 = RG_rl_165 ;
	7'h01 :
		TR_84 = RG_rl_165 ;
	7'h02 :
		TR_84 = RG_rl_165 ;
	7'h03 :
		TR_84 = RG_rl_165 ;
	7'h04 :
		TR_84 = RG_rl_165 ;
	7'h05 :
		TR_84 = RG_rl_165 ;
	7'h06 :
		TR_84 = RG_rl_165 ;
	7'h07 :
		TR_84 = RG_rl_165 ;
	7'h08 :
		TR_84 = RG_rl_165 ;
	7'h09 :
		TR_84 = RG_rl_165 ;
	7'h0a :
		TR_84 = RG_rl_165 ;
	7'h0b :
		TR_84 = RG_rl_165 ;
	7'h0c :
		TR_84 = RG_rl_165 ;
	7'h0d :
		TR_84 = RG_rl_165 ;
	7'h0e :
		TR_84 = RG_rl_165 ;
	7'h0f :
		TR_84 = RG_rl_165 ;
	7'h10 :
		TR_84 = RG_rl_165 ;
	7'h11 :
		TR_84 = RG_rl_165 ;
	7'h12 :
		TR_84 = RG_rl_165 ;
	7'h13 :
		TR_84 = RG_rl_165 ;
	7'h14 :
		TR_84 = RG_rl_165 ;
	7'h15 :
		TR_84 = RG_rl_165 ;
	7'h16 :
		TR_84 = RG_rl_165 ;
	7'h17 :
		TR_84 = RG_rl_165 ;
	7'h18 :
		TR_84 = RG_rl_165 ;
	7'h19 :
		TR_84 = RG_rl_165 ;
	7'h1a :
		TR_84 = RG_rl_165 ;
	7'h1b :
		TR_84 = RG_rl_165 ;
	7'h1c :
		TR_84 = RG_rl_165 ;
	7'h1d :
		TR_84 = RG_rl_165 ;
	7'h1e :
		TR_84 = RG_rl_165 ;
	7'h1f :
		TR_84 = RG_rl_165 ;
	7'h20 :
		TR_84 = RG_rl_165 ;
	7'h21 :
		TR_84 = RG_rl_165 ;
	7'h22 :
		TR_84 = RG_rl_165 ;
	7'h23 :
		TR_84 = RG_rl_165 ;
	7'h24 :
		TR_84 = RG_rl_165 ;
	7'h25 :
		TR_84 = RG_rl_165 ;
	7'h26 :
		TR_84 = RG_rl_165 ;
	7'h27 :
		TR_84 = RG_rl_165 ;
	7'h28 :
		TR_84 = RG_rl_165 ;
	7'h29 :
		TR_84 = RG_rl_165 ;
	7'h2a :
		TR_84 = RG_rl_165 ;
	7'h2b :
		TR_84 = RG_rl_165 ;
	7'h2c :
		TR_84 = RG_rl_165 ;
	7'h2d :
		TR_84 = RG_rl_165 ;
	7'h2e :
		TR_84 = RG_rl_165 ;
	7'h2f :
		TR_84 = RG_rl_165 ;
	7'h30 :
		TR_84 = RG_rl_165 ;
	7'h31 :
		TR_84 = RG_rl_165 ;
	7'h32 :
		TR_84 = RG_rl_165 ;
	7'h33 :
		TR_84 = RG_rl_165 ;
	7'h34 :
		TR_84 = RG_rl_165 ;
	7'h35 :
		TR_84 = RG_rl_165 ;
	7'h36 :
		TR_84 = RG_rl_165 ;
	7'h37 :
		TR_84 = RG_rl_165 ;
	7'h38 :
		TR_84 = RG_rl_165 ;
	7'h39 :
		TR_84 = RG_rl_165 ;
	7'h3a :
		TR_84 = RG_rl_165 ;
	7'h3b :
		TR_84 = RG_rl_165 ;
	7'h3c :
		TR_84 = RG_rl_165 ;
	7'h3d :
		TR_84 = RG_rl_165 ;
	7'h3e :
		TR_84 = RG_rl_165 ;
	7'h3f :
		TR_84 = RG_rl_165 ;
	7'h40 :
		TR_84 = RG_rl_165 ;
	7'h41 :
		TR_84 = RG_rl_165 ;
	7'h42 :
		TR_84 = RG_rl_165 ;
	7'h43 :
		TR_84 = RG_rl_165 ;
	7'h44 :
		TR_84 = RG_rl_165 ;
	7'h45 :
		TR_84 = RG_rl_165 ;
	7'h46 :
		TR_84 = RG_rl_165 ;
	7'h47 :
		TR_84 = RG_rl_165 ;
	7'h48 :
		TR_84 = 9'h000 ;	// line#=../rle.cpp:79
	7'h49 :
		TR_84 = RG_rl_165 ;
	7'h4a :
		TR_84 = RG_rl_165 ;
	7'h4b :
		TR_84 = RG_rl_165 ;
	7'h4c :
		TR_84 = RG_rl_165 ;
	7'h4d :
		TR_84 = RG_rl_165 ;
	7'h4e :
		TR_84 = RG_rl_165 ;
	7'h4f :
		TR_84 = RG_rl_165 ;
	7'h50 :
		TR_84 = RG_rl_165 ;
	7'h51 :
		TR_84 = RG_rl_165 ;
	7'h52 :
		TR_84 = RG_rl_165 ;
	7'h53 :
		TR_84 = RG_rl_165 ;
	7'h54 :
		TR_84 = RG_rl_165 ;
	7'h55 :
		TR_84 = RG_rl_165 ;
	7'h56 :
		TR_84 = RG_rl_165 ;
	7'h57 :
		TR_84 = RG_rl_165 ;
	7'h58 :
		TR_84 = RG_rl_165 ;
	7'h59 :
		TR_84 = RG_rl_165 ;
	7'h5a :
		TR_84 = RG_rl_165 ;
	7'h5b :
		TR_84 = RG_rl_165 ;
	7'h5c :
		TR_84 = RG_rl_165 ;
	7'h5d :
		TR_84 = RG_rl_165 ;
	7'h5e :
		TR_84 = RG_rl_165 ;
	7'h5f :
		TR_84 = RG_rl_165 ;
	7'h60 :
		TR_84 = RG_rl_165 ;
	7'h61 :
		TR_84 = RG_rl_165 ;
	7'h62 :
		TR_84 = RG_rl_165 ;
	7'h63 :
		TR_84 = RG_rl_165 ;
	7'h64 :
		TR_84 = RG_rl_165 ;
	7'h65 :
		TR_84 = RG_rl_165 ;
	7'h66 :
		TR_84 = RG_rl_165 ;
	7'h67 :
		TR_84 = RG_rl_165 ;
	7'h68 :
		TR_84 = RG_rl_165 ;
	7'h69 :
		TR_84 = RG_rl_165 ;
	7'h6a :
		TR_84 = RG_rl_165 ;
	7'h6b :
		TR_84 = RG_rl_165 ;
	7'h6c :
		TR_84 = RG_rl_165 ;
	7'h6d :
		TR_84 = RG_rl_165 ;
	7'h6e :
		TR_84 = RG_rl_165 ;
	7'h6f :
		TR_84 = RG_rl_165 ;
	7'h70 :
		TR_84 = RG_rl_165 ;
	7'h71 :
		TR_84 = RG_rl_165 ;
	7'h72 :
		TR_84 = RG_rl_165 ;
	7'h73 :
		TR_84 = RG_rl_165 ;
	7'h74 :
		TR_84 = RG_rl_165 ;
	7'h75 :
		TR_84 = RG_rl_165 ;
	7'h76 :
		TR_84 = RG_rl_165 ;
	7'h77 :
		TR_84 = RG_rl_165 ;
	7'h78 :
		TR_84 = RG_rl_165 ;
	7'h79 :
		TR_84 = RG_rl_165 ;
	7'h7a :
		TR_84 = RG_rl_165 ;
	7'h7b :
		TR_84 = RG_rl_165 ;
	7'h7c :
		TR_84 = RG_rl_165 ;
	7'h7d :
		TR_84 = RG_rl_165 ;
	7'h7e :
		TR_84 = RG_rl_165 ;
	7'h7f :
		TR_84 = RG_rl_165 ;
	default :
		TR_84 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_34 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h01 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h02 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h03 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h04 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h05 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h06 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h07 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h08 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h09 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h0a :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h0b :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h0c :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h0d :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h0e :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h0f :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h10 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h11 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h12 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h13 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h14 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h15 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h16 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h17 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h18 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h19 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h1a :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h1b :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h1c :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h1d :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h1e :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h1f :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h20 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h21 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h22 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h23 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h24 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h25 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h26 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h27 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h28 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h29 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h2a :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h2b :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h2c :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h2d :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h2e :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h2f :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h30 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h31 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h32 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h33 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h34 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h35 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h36 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h37 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h38 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h39 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h3a :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h3b :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h3c :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h3d :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h3e :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h3f :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h40 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h41 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h42 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h43 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h44 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h45 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h46 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h47 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h48 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h49 :
		TR_85 = 9'h000 ;	// line#=../rle.cpp:79
	7'h4a :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h4b :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h4c :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h4d :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h4e :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h4f :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h50 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h51 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h52 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h53 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h54 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h55 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h56 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h57 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h58 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h59 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h5a :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h5b :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h5c :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h5d :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h5e :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h5f :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h60 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h61 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h62 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h63 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h64 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h65 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h66 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h67 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h68 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h69 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h6a :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h6b :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h6c :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h6d :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h6e :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h6f :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h70 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h71 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h72 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h73 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h74 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h75 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h76 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h77 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h78 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h79 :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h7a :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h7b :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h7c :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h7d :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h7e :
		TR_85 = RG_quantized_block_rl_34 ;
	7'h7f :
		TR_85 = RG_quantized_block_rl_34 ;
	default :
		TR_85 = 9'hx ;
	endcase
always @ ( RG_rl_166 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_86 = RG_rl_166 ;
	7'h01 :
		TR_86 = RG_rl_166 ;
	7'h02 :
		TR_86 = RG_rl_166 ;
	7'h03 :
		TR_86 = RG_rl_166 ;
	7'h04 :
		TR_86 = RG_rl_166 ;
	7'h05 :
		TR_86 = RG_rl_166 ;
	7'h06 :
		TR_86 = RG_rl_166 ;
	7'h07 :
		TR_86 = RG_rl_166 ;
	7'h08 :
		TR_86 = RG_rl_166 ;
	7'h09 :
		TR_86 = RG_rl_166 ;
	7'h0a :
		TR_86 = RG_rl_166 ;
	7'h0b :
		TR_86 = RG_rl_166 ;
	7'h0c :
		TR_86 = RG_rl_166 ;
	7'h0d :
		TR_86 = RG_rl_166 ;
	7'h0e :
		TR_86 = RG_rl_166 ;
	7'h0f :
		TR_86 = RG_rl_166 ;
	7'h10 :
		TR_86 = RG_rl_166 ;
	7'h11 :
		TR_86 = RG_rl_166 ;
	7'h12 :
		TR_86 = RG_rl_166 ;
	7'h13 :
		TR_86 = RG_rl_166 ;
	7'h14 :
		TR_86 = RG_rl_166 ;
	7'h15 :
		TR_86 = RG_rl_166 ;
	7'h16 :
		TR_86 = RG_rl_166 ;
	7'h17 :
		TR_86 = RG_rl_166 ;
	7'h18 :
		TR_86 = RG_rl_166 ;
	7'h19 :
		TR_86 = RG_rl_166 ;
	7'h1a :
		TR_86 = RG_rl_166 ;
	7'h1b :
		TR_86 = RG_rl_166 ;
	7'h1c :
		TR_86 = RG_rl_166 ;
	7'h1d :
		TR_86 = RG_rl_166 ;
	7'h1e :
		TR_86 = RG_rl_166 ;
	7'h1f :
		TR_86 = RG_rl_166 ;
	7'h20 :
		TR_86 = RG_rl_166 ;
	7'h21 :
		TR_86 = RG_rl_166 ;
	7'h22 :
		TR_86 = RG_rl_166 ;
	7'h23 :
		TR_86 = RG_rl_166 ;
	7'h24 :
		TR_86 = RG_rl_166 ;
	7'h25 :
		TR_86 = RG_rl_166 ;
	7'h26 :
		TR_86 = RG_rl_166 ;
	7'h27 :
		TR_86 = RG_rl_166 ;
	7'h28 :
		TR_86 = RG_rl_166 ;
	7'h29 :
		TR_86 = RG_rl_166 ;
	7'h2a :
		TR_86 = RG_rl_166 ;
	7'h2b :
		TR_86 = RG_rl_166 ;
	7'h2c :
		TR_86 = RG_rl_166 ;
	7'h2d :
		TR_86 = RG_rl_166 ;
	7'h2e :
		TR_86 = RG_rl_166 ;
	7'h2f :
		TR_86 = RG_rl_166 ;
	7'h30 :
		TR_86 = RG_rl_166 ;
	7'h31 :
		TR_86 = RG_rl_166 ;
	7'h32 :
		TR_86 = RG_rl_166 ;
	7'h33 :
		TR_86 = RG_rl_166 ;
	7'h34 :
		TR_86 = RG_rl_166 ;
	7'h35 :
		TR_86 = RG_rl_166 ;
	7'h36 :
		TR_86 = RG_rl_166 ;
	7'h37 :
		TR_86 = RG_rl_166 ;
	7'h38 :
		TR_86 = RG_rl_166 ;
	7'h39 :
		TR_86 = RG_rl_166 ;
	7'h3a :
		TR_86 = RG_rl_166 ;
	7'h3b :
		TR_86 = RG_rl_166 ;
	7'h3c :
		TR_86 = RG_rl_166 ;
	7'h3d :
		TR_86 = RG_rl_166 ;
	7'h3e :
		TR_86 = RG_rl_166 ;
	7'h3f :
		TR_86 = RG_rl_166 ;
	7'h40 :
		TR_86 = RG_rl_166 ;
	7'h41 :
		TR_86 = RG_rl_166 ;
	7'h42 :
		TR_86 = RG_rl_166 ;
	7'h43 :
		TR_86 = RG_rl_166 ;
	7'h44 :
		TR_86 = RG_rl_166 ;
	7'h45 :
		TR_86 = RG_rl_166 ;
	7'h46 :
		TR_86 = RG_rl_166 ;
	7'h47 :
		TR_86 = RG_rl_166 ;
	7'h48 :
		TR_86 = RG_rl_166 ;
	7'h49 :
		TR_86 = RG_rl_166 ;
	7'h4a :
		TR_86 = 9'h000 ;	// line#=../rle.cpp:79
	7'h4b :
		TR_86 = RG_rl_166 ;
	7'h4c :
		TR_86 = RG_rl_166 ;
	7'h4d :
		TR_86 = RG_rl_166 ;
	7'h4e :
		TR_86 = RG_rl_166 ;
	7'h4f :
		TR_86 = RG_rl_166 ;
	7'h50 :
		TR_86 = RG_rl_166 ;
	7'h51 :
		TR_86 = RG_rl_166 ;
	7'h52 :
		TR_86 = RG_rl_166 ;
	7'h53 :
		TR_86 = RG_rl_166 ;
	7'h54 :
		TR_86 = RG_rl_166 ;
	7'h55 :
		TR_86 = RG_rl_166 ;
	7'h56 :
		TR_86 = RG_rl_166 ;
	7'h57 :
		TR_86 = RG_rl_166 ;
	7'h58 :
		TR_86 = RG_rl_166 ;
	7'h59 :
		TR_86 = RG_rl_166 ;
	7'h5a :
		TR_86 = RG_rl_166 ;
	7'h5b :
		TR_86 = RG_rl_166 ;
	7'h5c :
		TR_86 = RG_rl_166 ;
	7'h5d :
		TR_86 = RG_rl_166 ;
	7'h5e :
		TR_86 = RG_rl_166 ;
	7'h5f :
		TR_86 = RG_rl_166 ;
	7'h60 :
		TR_86 = RG_rl_166 ;
	7'h61 :
		TR_86 = RG_rl_166 ;
	7'h62 :
		TR_86 = RG_rl_166 ;
	7'h63 :
		TR_86 = RG_rl_166 ;
	7'h64 :
		TR_86 = RG_rl_166 ;
	7'h65 :
		TR_86 = RG_rl_166 ;
	7'h66 :
		TR_86 = RG_rl_166 ;
	7'h67 :
		TR_86 = RG_rl_166 ;
	7'h68 :
		TR_86 = RG_rl_166 ;
	7'h69 :
		TR_86 = RG_rl_166 ;
	7'h6a :
		TR_86 = RG_rl_166 ;
	7'h6b :
		TR_86 = RG_rl_166 ;
	7'h6c :
		TR_86 = RG_rl_166 ;
	7'h6d :
		TR_86 = RG_rl_166 ;
	7'h6e :
		TR_86 = RG_rl_166 ;
	7'h6f :
		TR_86 = RG_rl_166 ;
	7'h70 :
		TR_86 = RG_rl_166 ;
	7'h71 :
		TR_86 = RG_rl_166 ;
	7'h72 :
		TR_86 = RG_rl_166 ;
	7'h73 :
		TR_86 = RG_rl_166 ;
	7'h74 :
		TR_86 = RG_rl_166 ;
	7'h75 :
		TR_86 = RG_rl_166 ;
	7'h76 :
		TR_86 = RG_rl_166 ;
	7'h77 :
		TR_86 = RG_rl_166 ;
	7'h78 :
		TR_86 = RG_rl_166 ;
	7'h79 :
		TR_86 = RG_rl_166 ;
	7'h7a :
		TR_86 = RG_rl_166 ;
	7'h7b :
		TR_86 = RG_rl_166 ;
	7'h7c :
		TR_86 = RG_rl_166 ;
	7'h7d :
		TR_86 = RG_rl_166 ;
	7'h7e :
		TR_86 = RG_rl_166 ;
	7'h7f :
		TR_86 = RG_rl_166 ;
	default :
		TR_86 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_35 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h01 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h02 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h03 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h04 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h05 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h06 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h07 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h08 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h09 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h0a :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h0b :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h0c :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h0d :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h0e :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h0f :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h10 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h11 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h12 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h13 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h14 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h15 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h16 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h17 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h18 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h19 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h1a :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h1b :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h1c :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h1d :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h1e :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h1f :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h20 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h21 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h22 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h23 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h24 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h25 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h26 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h27 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h28 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h29 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h2a :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h2b :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h2c :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h2d :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h2e :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h2f :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h30 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h31 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h32 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h33 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h34 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h35 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h36 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h37 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h38 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h39 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h3a :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h3b :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h3c :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h3d :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h3e :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h3f :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h40 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h41 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h42 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h43 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h44 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h45 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h46 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h47 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h48 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h49 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h4a :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h4b :
		TR_87 = 9'h000 ;	// line#=../rle.cpp:79
	7'h4c :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h4d :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h4e :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h4f :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h50 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h51 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h52 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h53 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h54 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h55 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h56 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h57 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h58 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h59 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h5a :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h5b :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h5c :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h5d :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h5e :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h5f :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h60 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h61 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h62 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h63 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h64 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h65 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h66 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h67 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h68 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h69 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h6a :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h6b :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h6c :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h6d :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h6e :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h6f :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h70 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h71 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h72 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h73 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h74 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h75 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h76 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h77 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h78 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h79 :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h7a :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h7b :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h7c :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h7d :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h7e :
		TR_87 = RG_quantized_block_rl_35 ;
	7'h7f :
		TR_87 = RG_quantized_block_rl_35 ;
	default :
		TR_87 = 9'hx ;
	endcase
always @ ( RG_rl_167 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_88 = RG_rl_167 ;
	7'h01 :
		TR_88 = RG_rl_167 ;
	7'h02 :
		TR_88 = RG_rl_167 ;
	7'h03 :
		TR_88 = RG_rl_167 ;
	7'h04 :
		TR_88 = RG_rl_167 ;
	7'h05 :
		TR_88 = RG_rl_167 ;
	7'h06 :
		TR_88 = RG_rl_167 ;
	7'h07 :
		TR_88 = RG_rl_167 ;
	7'h08 :
		TR_88 = RG_rl_167 ;
	7'h09 :
		TR_88 = RG_rl_167 ;
	7'h0a :
		TR_88 = RG_rl_167 ;
	7'h0b :
		TR_88 = RG_rl_167 ;
	7'h0c :
		TR_88 = RG_rl_167 ;
	7'h0d :
		TR_88 = RG_rl_167 ;
	7'h0e :
		TR_88 = RG_rl_167 ;
	7'h0f :
		TR_88 = RG_rl_167 ;
	7'h10 :
		TR_88 = RG_rl_167 ;
	7'h11 :
		TR_88 = RG_rl_167 ;
	7'h12 :
		TR_88 = RG_rl_167 ;
	7'h13 :
		TR_88 = RG_rl_167 ;
	7'h14 :
		TR_88 = RG_rl_167 ;
	7'h15 :
		TR_88 = RG_rl_167 ;
	7'h16 :
		TR_88 = RG_rl_167 ;
	7'h17 :
		TR_88 = RG_rl_167 ;
	7'h18 :
		TR_88 = RG_rl_167 ;
	7'h19 :
		TR_88 = RG_rl_167 ;
	7'h1a :
		TR_88 = RG_rl_167 ;
	7'h1b :
		TR_88 = RG_rl_167 ;
	7'h1c :
		TR_88 = RG_rl_167 ;
	7'h1d :
		TR_88 = RG_rl_167 ;
	7'h1e :
		TR_88 = RG_rl_167 ;
	7'h1f :
		TR_88 = RG_rl_167 ;
	7'h20 :
		TR_88 = RG_rl_167 ;
	7'h21 :
		TR_88 = RG_rl_167 ;
	7'h22 :
		TR_88 = RG_rl_167 ;
	7'h23 :
		TR_88 = RG_rl_167 ;
	7'h24 :
		TR_88 = RG_rl_167 ;
	7'h25 :
		TR_88 = RG_rl_167 ;
	7'h26 :
		TR_88 = RG_rl_167 ;
	7'h27 :
		TR_88 = RG_rl_167 ;
	7'h28 :
		TR_88 = RG_rl_167 ;
	7'h29 :
		TR_88 = RG_rl_167 ;
	7'h2a :
		TR_88 = RG_rl_167 ;
	7'h2b :
		TR_88 = RG_rl_167 ;
	7'h2c :
		TR_88 = RG_rl_167 ;
	7'h2d :
		TR_88 = RG_rl_167 ;
	7'h2e :
		TR_88 = RG_rl_167 ;
	7'h2f :
		TR_88 = RG_rl_167 ;
	7'h30 :
		TR_88 = RG_rl_167 ;
	7'h31 :
		TR_88 = RG_rl_167 ;
	7'h32 :
		TR_88 = RG_rl_167 ;
	7'h33 :
		TR_88 = RG_rl_167 ;
	7'h34 :
		TR_88 = RG_rl_167 ;
	7'h35 :
		TR_88 = RG_rl_167 ;
	7'h36 :
		TR_88 = RG_rl_167 ;
	7'h37 :
		TR_88 = RG_rl_167 ;
	7'h38 :
		TR_88 = RG_rl_167 ;
	7'h39 :
		TR_88 = RG_rl_167 ;
	7'h3a :
		TR_88 = RG_rl_167 ;
	7'h3b :
		TR_88 = RG_rl_167 ;
	7'h3c :
		TR_88 = RG_rl_167 ;
	7'h3d :
		TR_88 = RG_rl_167 ;
	7'h3e :
		TR_88 = RG_rl_167 ;
	7'h3f :
		TR_88 = RG_rl_167 ;
	7'h40 :
		TR_88 = RG_rl_167 ;
	7'h41 :
		TR_88 = RG_rl_167 ;
	7'h42 :
		TR_88 = RG_rl_167 ;
	7'h43 :
		TR_88 = RG_rl_167 ;
	7'h44 :
		TR_88 = RG_rl_167 ;
	7'h45 :
		TR_88 = RG_rl_167 ;
	7'h46 :
		TR_88 = RG_rl_167 ;
	7'h47 :
		TR_88 = RG_rl_167 ;
	7'h48 :
		TR_88 = RG_rl_167 ;
	7'h49 :
		TR_88 = RG_rl_167 ;
	7'h4a :
		TR_88 = RG_rl_167 ;
	7'h4b :
		TR_88 = RG_rl_167 ;
	7'h4c :
		TR_88 = 9'h000 ;	// line#=../rle.cpp:79
	7'h4d :
		TR_88 = RG_rl_167 ;
	7'h4e :
		TR_88 = RG_rl_167 ;
	7'h4f :
		TR_88 = RG_rl_167 ;
	7'h50 :
		TR_88 = RG_rl_167 ;
	7'h51 :
		TR_88 = RG_rl_167 ;
	7'h52 :
		TR_88 = RG_rl_167 ;
	7'h53 :
		TR_88 = RG_rl_167 ;
	7'h54 :
		TR_88 = RG_rl_167 ;
	7'h55 :
		TR_88 = RG_rl_167 ;
	7'h56 :
		TR_88 = RG_rl_167 ;
	7'h57 :
		TR_88 = RG_rl_167 ;
	7'h58 :
		TR_88 = RG_rl_167 ;
	7'h59 :
		TR_88 = RG_rl_167 ;
	7'h5a :
		TR_88 = RG_rl_167 ;
	7'h5b :
		TR_88 = RG_rl_167 ;
	7'h5c :
		TR_88 = RG_rl_167 ;
	7'h5d :
		TR_88 = RG_rl_167 ;
	7'h5e :
		TR_88 = RG_rl_167 ;
	7'h5f :
		TR_88 = RG_rl_167 ;
	7'h60 :
		TR_88 = RG_rl_167 ;
	7'h61 :
		TR_88 = RG_rl_167 ;
	7'h62 :
		TR_88 = RG_rl_167 ;
	7'h63 :
		TR_88 = RG_rl_167 ;
	7'h64 :
		TR_88 = RG_rl_167 ;
	7'h65 :
		TR_88 = RG_rl_167 ;
	7'h66 :
		TR_88 = RG_rl_167 ;
	7'h67 :
		TR_88 = RG_rl_167 ;
	7'h68 :
		TR_88 = RG_rl_167 ;
	7'h69 :
		TR_88 = RG_rl_167 ;
	7'h6a :
		TR_88 = RG_rl_167 ;
	7'h6b :
		TR_88 = RG_rl_167 ;
	7'h6c :
		TR_88 = RG_rl_167 ;
	7'h6d :
		TR_88 = RG_rl_167 ;
	7'h6e :
		TR_88 = RG_rl_167 ;
	7'h6f :
		TR_88 = RG_rl_167 ;
	7'h70 :
		TR_88 = RG_rl_167 ;
	7'h71 :
		TR_88 = RG_rl_167 ;
	7'h72 :
		TR_88 = RG_rl_167 ;
	7'h73 :
		TR_88 = RG_rl_167 ;
	7'h74 :
		TR_88 = RG_rl_167 ;
	7'h75 :
		TR_88 = RG_rl_167 ;
	7'h76 :
		TR_88 = RG_rl_167 ;
	7'h77 :
		TR_88 = RG_rl_167 ;
	7'h78 :
		TR_88 = RG_rl_167 ;
	7'h79 :
		TR_88 = RG_rl_167 ;
	7'h7a :
		TR_88 = RG_rl_167 ;
	7'h7b :
		TR_88 = RG_rl_167 ;
	7'h7c :
		TR_88 = RG_rl_167 ;
	7'h7d :
		TR_88 = RG_rl_167 ;
	7'h7e :
		TR_88 = RG_rl_167 ;
	7'h7f :
		TR_88 = RG_rl_167 ;
	default :
		TR_88 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_36 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h01 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h02 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h03 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h04 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h05 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h06 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h07 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h08 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h09 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h0a :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h0b :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h0c :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h0d :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h0e :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h0f :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h10 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h11 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h12 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h13 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h14 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h15 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h16 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h17 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h18 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h19 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h1a :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h1b :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h1c :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h1d :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h1e :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h1f :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h20 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h21 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h22 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h23 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h24 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h25 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h26 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h27 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h28 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h29 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h2a :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h2b :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h2c :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h2d :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h2e :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h2f :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h30 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h31 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h32 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h33 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h34 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h35 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h36 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h37 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h38 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h39 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h3a :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h3b :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h3c :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h3d :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h3e :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h3f :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h40 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h41 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h42 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h43 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h44 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h45 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h46 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h47 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h48 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h49 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h4a :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h4b :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h4c :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h4d :
		TR_89 = 9'h000 ;	// line#=../rle.cpp:79
	7'h4e :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h4f :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h50 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h51 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h52 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h53 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h54 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h55 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h56 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h57 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h58 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h59 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h5a :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h5b :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h5c :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h5d :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h5e :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h5f :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h60 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h61 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h62 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h63 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h64 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h65 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h66 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h67 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h68 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h69 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h6a :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h6b :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h6c :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h6d :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h6e :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h6f :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h70 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h71 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h72 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h73 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h74 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h75 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h76 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h77 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h78 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h79 :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h7a :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h7b :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h7c :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h7d :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h7e :
		TR_89 = RG_quantized_block_rl_36 ;
	7'h7f :
		TR_89 = RG_quantized_block_rl_36 ;
	default :
		TR_89 = 9'hx ;
	endcase
always @ ( RG_rl_168 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_90 = RG_rl_168 ;
	7'h01 :
		TR_90 = RG_rl_168 ;
	7'h02 :
		TR_90 = RG_rl_168 ;
	7'h03 :
		TR_90 = RG_rl_168 ;
	7'h04 :
		TR_90 = RG_rl_168 ;
	7'h05 :
		TR_90 = RG_rl_168 ;
	7'h06 :
		TR_90 = RG_rl_168 ;
	7'h07 :
		TR_90 = RG_rl_168 ;
	7'h08 :
		TR_90 = RG_rl_168 ;
	7'h09 :
		TR_90 = RG_rl_168 ;
	7'h0a :
		TR_90 = RG_rl_168 ;
	7'h0b :
		TR_90 = RG_rl_168 ;
	7'h0c :
		TR_90 = RG_rl_168 ;
	7'h0d :
		TR_90 = RG_rl_168 ;
	7'h0e :
		TR_90 = RG_rl_168 ;
	7'h0f :
		TR_90 = RG_rl_168 ;
	7'h10 :
		TR_90 = RG_rl_168 ;
	7'h11 :
		TR_90 = RG_rl_168 ;
	7'h12 :
		TR_90 = RG_rl_168 ;
	7'h13 :
		TR_90 = RG_rl_168 ;
	7'h14 :
		TR_90 = RG_rl_168 ;
	7'h15 :
		TR_90 = RG_rl_168 ;
	7'h16 :
		TR_90 = RG_rl_168 ;
	7'h17 :
		TR_90 = RG_rl_168 ;
	7'h18 :
		TR_90 = RG_rl_168 ;
	7'h19 :
		TR_90 = RG_rl_168 ;
	7'h1a :
		TR_90 = RG_rl_168 ;
	7'h1b :
		TR_90 = RG_rl_168 ;
	7'h1c :
		TR_90 = RG_rl_168 ;
	7'h1d :
		TR_90 = RG_rl_168 ;
	7'h1e :
		TR_90 = RG_rl_168 ;
	7'h1f :
		TR_90 = RG_rl_168 ;
	7'h20 :
		TR_90 = RG_rl_168 ;
	7'h21 :
		TR_90 = RG_rl_168 ;
	7'h22 :
		TR_90 = RG_rl_168 ;
	7'h23 :
		TR_90 = RG_rl_168 ;
	7'h24 :
		TR_90 = RG_rl_168 ;
	7'h25 :
		TR_90 = RG_rl_168 ;
	7'h26 :
		TR_90 = RG_rl_168 ;
	7'h27 :
		TR_90 = RG_rl_168 ;
	7'h28 :
		TR_90 = RG_rl_168 ;
	7'h29 :
		TR_90 = RG_rl_168 ;
	7'h2a :
		TR_90 = RG_rl_168 ;
	7'h2b :
		TR_90 = RG_rl_168 ;
	7'h2c :
		TR_90 = RG_rl_168 ;
	7'h2d :
		TR_90 = RG_rl_168 ;
	7'h2e :
		TR_90 = RG_rl_168 ;
	7'h2f :
		TR_90 = RG_rl_168 ;
	7'h30 :
		TR_90 = RG_rl_168 ;
	7'h31 :
		TR_90 = RG_rl_168 ;
	7'h32 :
		TR_90 = RG_rl_168 ;
	7'h33 :
		TR_90 = RG_rl_168 ;
	7'h34 :
		TR_90 = RG_rl_168 ;
	7'h35 :
		TR_90 = RG_rl_168 ;
	7'h36 :
		TR_90 = RG_rl_168 ;
	7'h37 :
		TR_90 = RG_rl_168 ;
	7'h38 :
		TR_90 = RG_rl_168 ;
	7'h39 :
		TR_90 = RG_rl_168 ;
	7'h3a :
		TR_90 = RG_rl_168 ;
	7'h3b :
		TR_90 = RG_rl_168 ;
	7'h3c :
		TR_90 = RG_rl_168 ;
	7'h3d :
		TR_90 = RG_rl_168 ;
	7'h3e :
		TR_90 = RG_rl_168 ;
	7'h3f :
		TR_90 = RG_rl_168 ;
	7'h40 :
		TR_90 = RG_rl_168 ;
	7'h41 :
		TR_90 = RG_rl_168 ;
	7'h42 :
		TR_90 = RG_rl_168 ;
	7'h43 :
		TR_90 = RG_rl_168 ;
	7'h44 :
		TR_90 = RG_rl_168 ;
	7'h45 :
		TR_90 = RG_rl_168 ;
	7'h46 :
		TR_90 = RG_rl_168 ;
	7'h47 :
		TR_90 = RG_rl_168 ;
	7'h48 :
		TR_90 = RG_rl_168 ;
	7'h49 :
		TR_90 = RG_rl_168 ;
	7'h4a :
		TR_90 = RG_rl_168 ;
	7'h4b :
		TR_90 = RG_rl_168 ;
	7'h4c :
		TR_90 = RG_rl_168 ;
	7'h4d :
		TR_90 = RG_rl_168 ;
	7'h4e :
		TR_90 = 9'h000 ;	// line#=../rle.cpp:79
	7'h4f :
		TR_90 = RG_rl_168 ;
	7'h50 :
		TR_90 = RG_rl_168 ;
	7'h51 :
		TR_90 = RG_rl_168 ;
	7'h52 :
		TR_90 = RG_rl_168 ;
	7'h53 :
		TR_90 = RG_rl_168 ;
	7'h54 :
		TR_90 = RG_rl_168 ;
	7'h55 :
		TR_90 = RG_rl_168 ;
	7'h56 :
		TR_90 = RG_rl_168 ;
	7'h57 :
		TR_90 = RG_rl_168 ;
	7'h58 :
		TR_90 = RG_rl_168 ;
	7'h59 :
		TR_90 = RG_rl_168 ;
	7'h5a :
		TR_90 = RG_rl_168 ;
	7'h5b :
		TR_90 = RG_rl_168 ;
	7'h5c :
		TR_90 = RG_rl_168 ;
	7'h5d :
		TR_90 = RG_rl_168 ;
	7'h5e :
		TR_90 = RG_rl_168 ;
	7'h5f :
		TR_90 = RG_rl_168 ;
	7'h60 :
		TR_90 = RG_rl_168 ;
	7'h61 :
		TR_90 = RG_rl_168 ;
	7'h62 :
		TR_90 = RG_rl_168 ;
	7'h63 :
		TR_90 = RG_rl_168 ;
	7'h64 :
		TR_90 = RG_rl_168 ;
	7'h65 :
		TR_90 = RG_rl_168 ;
	7'h66 :
		TR_90 = RG_rl_168 ;
	7'h67 :
		TR_90 = RG_rl_168 ;
	7'h68 :
		TR_90 = RG_rl_168 ;
	7'h69 :
		TR_90 = RG_rl_168 ;
	7'h6a :
		TR_90 = RG_rl_168 ;
	7'h6b :
		TR_90 = RG_rl_168 ;
	7'h6c :
		TR_90 = RG_rl_168 ;
	7'h6d :
		TR_90 = RG_rl_168 ;
	7'h6e :
		TR_90 = RG_rl_168 ;
	7'h6f :
		TR_90 = RG_rl_168 ;
	7'h70 :
		TR_90 = RG_rl_168 ;
	7'h71 :
		TR_90 = RG_rl_168 ;
	7'h72 :
		TR_90 = RG_rl_168 ;
	7'h73 :
		TR_90 = RG_rl_168 ;
	7'h74 :
		TR_90 = RG_rl_168 ;
	7'h75 :
		TR_90 = RG_rl_168 ;
	7'h76 :
		TR_90 = RG_rl_168 ;
	7'h77 :
		TR_90 = RG_rl_168 ;
	7'h78 :
		TR_90 = RG_rl_168 ;
	7'h79 :
		TR_90 = RG_rl_168 ;
	7'h7a :
		TR_90 = RG_rl_168 ;
	7'h7b :
		TR_90 = RG_rl_168 ;
	7'h7c :
		TR_90 = RG_rl_168 ;
	7'h7d :
		TR_90 = RG_rl_168 ;
	7'h7e :
		TR_90 = RG_rl_168 ;
	7'h7f :
		TR_90 = RG_rl_168 ;
	default :
		TR_90 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_37 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h01 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h02 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h03 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h04 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h05 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h06 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h07 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h08 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h09 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h0a :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h0b :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h0c :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h0d :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h0e :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h0f :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h10 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h11 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h12 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h13 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h14 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h15 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h16 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h17 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h18 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h19 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h1a :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h1b :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h1c :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h1d :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h1e :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h1f :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h20 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h21 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h22 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h23 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h24 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h25 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h26 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h27 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h28 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h29 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h2a :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h2b :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h2c :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h2d :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h2e :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h2f :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h30 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h31 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h32 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h33 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h34 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h35 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h36 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h37 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h38 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h39 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h3a :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h3b :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h3c :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h3d :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h3e :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h3f :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h40 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h41 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h42 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h43 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h44 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h45 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h46 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h47 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h48 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h49 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h4a :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h4b :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h4c :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h4d :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h4e :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h4f :
		TR_91 = 9'h000 ;	// line#=../rle.cpp:79
	7'h50 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h51 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h52 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h53 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h54 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h55 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h56 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h57 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h58 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h59 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h5a :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h5b :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h5c :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h5d :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h5e :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h5f :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h60 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h61 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h62 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h63 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h64 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h65 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h66 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h67 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h68 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h69 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h6a :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h6b :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h6c :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h6d :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h6e :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h6f :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h70 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h71 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h72 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h73 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h74 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h75 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h76 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h77 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h78 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h79 :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h7a :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h7b :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h7c :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h7d :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h7e :
		TR_91 = RG_quantized_block_rl_37 ;
	7'h7f :
		TR_91 = RG_quantized_block_rl_37 ;
	default :
		TR_91 = 9'hx ;
	endcase
always @ ( RG_rl_169 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_92 = RG_rl_169 ;
	7'h01 :
		TR_92 = RG_rl_169 ;
	7'h02 :
		TR_92 = RG_rl_169 ;
	7'h03 :
		TR_92 = RG_rl_169 ;
	7'h04 :
		TR_92 = RG_rl_169 ;
	7'h05 :
		TR_92 = RG_rl_169 ;
	7'h06 :
		TR_92 = RG_rl_169 ;
	7'h07 :
		TR_92 = RG_rl_169 ;
	7'h08 :
		TR_92 = RG_rl_169 ;
	7'h09 :
		TR_92 = RG_rl_169 ;
	7'h0a :
		TR_92 = RG_rl_169 ;
	7'h0b :
		TR_92 = RG_rl_169 ;
	7'h0c :
		TR_92 = RG_rl_169 ;
	7'h0d :
		TR_92 = RG_rl_169 ;
	7'h0e :
		TR_92 = RG_rl_169 ;
	7'h0f :
		TR_92 = RG_rl_169 ;
	7'h10 :
		TR_92 = RG_rl_169 ;
	7'h11 :
		TR_92 = RG_rl_169 ;
	7'h12 :
		TR_92 = RG_rl_169 ;
	7'h13 :
		TR_92 = RG_rl_169 ;
	7'h14 :
		TR_92 = RG_rl_169 ;
	7'h15 :
		TR_92 = RG_rl_169 ;
	7'h16 :
		TR_92 = RG_rl_169 ;
	7'h17 :
		TR_92 = RG_rl_169 ;
	7'h18 :
		TR_92 = RG_rl_169 ;
	7'h19 :
		TR_92 = RG_rl_169 ;
	7'h1a :
		TR_92 = RG_rl_169 ;
	7'h1b :
		TR_92 = RG_rl_169 ;
	7'h1c :
		TR_92 = RG_rl_169 ;
	7'h1d :
		TR_92 = RG_rl_169 ;
	7'h1e :
		TR_92 = RG_rl_169 ;
	7'h1f :
		TR_92 = RG_rl_169 ;
	7'h20 :
		TR_92 = RG_rl_169 ;
	7'h21 :
		TR_92 = RG_rl_169 ;
	7'h22 :
		TR_92 = RG_rl_169 ;
	7'h23 :
		TR_92 = RG_rl_169 ;
	7'h24 :
		TR_92 = RG_rl_169 ;
	7'h25 :
		TR_92 = RG_rl_169 ;
	7'h26 :
		TR_92 = RG_rl_169 ;
	7'h27 :
		TR_92 = RG_rl_169 ;
	7'h28 :
		TR_92 = RG_rl_169 ;
	7'h29 :
		TR_92 = RG_rl_169 ;
	7'h2a :
		TR_92 = RG_rl_169 ;
	7'h2b :
		TR_92 = RG_rl_169 ;
	7'h2c :
		TR_92 = RG_rl_169 ;
	7'h2d :
		TR_92 = RG_rl_169 ;
	7'h2e :
		TR_92 = RG_rl_169 ;
	7'h2f :
		TR_92 = RG_rl_169 ;
	7'h30 :
		TR_92 = RG_rl_169 ;
	7'h31 :
		TR_92 = RG_rl_169 ;
	7'h32 :
		TR_92 = RG_rl_169 ;
	7'h33 :
		TR_92 = RG_rl_169 ;
	7'h34 :
		TR_92 = RG_rl_169 ;
	7'h35 :
		TR_92 = RG_rl_169 ;
	7'h36 :
		TR_92 = RG_rl_169 ;
	7'h37 :
		TR_92 = RG_rl_169 ;
	7'h38 :
		TR_92 = RG_rl_169 ;
	7'h39 :
		TR_92 = RG_rl_169 ;
	7'h3a :
		TR_92 = RG_rl_169 ;
	7'h3b :
		TR_92 = RG_rl_169 ;
	7'h3c :
		TR_92 = RG_rl_169 ;
	7'h3d :
		TR_92 = RG_rl_169 ;
	7'h3e :
		TR_92 = RG_rl_169 ;
	7'h3f :
		TR_92 = RG_rl_169 ;
	7'h40 :
		TR_92 = RG_rl_169 ;
	7'h41 :
		TR_92 = RG_rl_169 ;
	7'h42 :
		TR_92 = RG_rl_169 ;
	7'h43 :
		TR_92 = RG_rl_169 ;
	7'h44 :
		TR_92 = RG_rl_169 ;
	7'h45 :
		TR_92 = RG_rl_169 ;
	7'h46 :
		TR_92 = RG_rl_169 ;
	7'h47 :
		TR_92 = RG_rl_169 ;
	7'h48 :
		TR_92 = RG_rl_169 ;
	7'h49 :
		TR_92 = RG_rl_169 ;
	7'h4a :
		TR_92 = RG_rl_169 ;
	7'h4b :
		TR_92 = RG_rl_169 ;
	7'h4c :
		TR_92 = RG_rl_169 ;
	7'h4d :
		TR_92 = RG_rl_169 ;
	7'h4e :
		TR_92 = RG_rl_169 ;
	7'h4f :
		TR_92 = RG_rl_169 ;
	7'h50 :
		TR_92 = 9'h000 ;	// line#=../rle.cpp:79
	7'h51 :
		TR_92 = RG_rl_169 ;
	7'h52 :
		TR_92 = RG_rl_169 ;
	7'h53 :
		TR_92 = RG_rl_169 ;
	7'h54 :
		TR_92 = RG_rl_169 ;
	7'h55 :
		TR_92 = RG_rl_169 ;
	7'h56 :
		TR_92 = RG_rl_169 ;
	7'h57 :
		TR_92 = RG_rl_169 ;
	7'h58 :
		TR_92 = RG_rl_169 ;
	7'h59 :
		TR_92 = RG_rl_169 ;
	7'h5a :
		TR_92 = RG_rl_169 ;
	7'h5b :
		TR_92 = RG_rl_169 ;
	7'h5c :
		TR_92 = RG_rl_169 ;
	7'h5d :
		TR_92 = RG_rl_169 ;
	7'h5e :
		TR_92 = RG_rl_169 ;
	7'h5f :
		TR_92 = RG_rl_169 ;
	7'h60 :
		TR_92 = RG_rl_169 ;
	7'h61 :
		TR_92 = RG_rl_169 ;
	7'h62 :
		TR_92 = RG_rl_169 ;
	7'h63 :
		TR_92 = RG_rl_169 ;
	7'h64 :
		TR_92 = RG_rl_169 ;
	7'h65 :
		TR_92 = RG_rl_169 ;
	7'h66 :
		TR_92 = RG_rl_169 ;
	7'h67 :
		TR_92 = RG_rl_169 ;
	7'h68 :
		TR_92 = RG_rl_169 ;
	7'h69 :
		TR_92 = RG_rl_169 ;
	7'h6a :
		TR_92 = RG_rl_169 ;
	7'h6b :
		TR_92 = RG_rl_169 ;
	7'h6c :
		TR_92 = RG_rl_169 ;
	7'h6d :
		TR_92 = RG_rl_169 ;
	7'h6e :
		TR_92 = RG_rl_169 ;
	7'h6f :
		TR_92 = RG_rl_169 ;
	7'h70 :
		TR_92 = RG_rl_169 ;
	7'h71 :
		TR_92 = RG_rl_169 ;
	7'h72 :
		TR_92 = RG_rl_169 ;
	7'h73 :
		TR_92 = RG_rl_169 ;
	7'h74 :
		TR_92 = RG_rl_169 ;
	7'h75 :
		TR_92 = RG_rl_169 ;
	7'h76 :
		TR_92 = RG_rl_169 ;
	7'h77 :
		TR_92 = RG_rl_169 ;
	7'h78 :
		TR_92 = RG_rl_169 ;
	7'h79 :
		TR_92 = RG_rl_169 ;
	7'h7a :
		TR_92 = RG_rl_169 ;
	7'h7b :
		TR_92 = RG_rl_169 ;
	7'h7c :
		TR_92 = RG_rl_169 ;
	7'h7d :
		TR_92 = RG_rl_169 ;
	7'h7e :
		TR_92 = RG_rl_169 ;
	7'h7f :
		TR_92 = RG_rl_169 ;
	default :
		TR_92 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_38 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h01 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h02 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h03 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h04 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h05 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h06 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h07 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h08 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h09 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h0a :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h0b :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h0c :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h0d :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h0e :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h0f :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h10 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h11 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h12 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h13 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h14 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h15 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h16 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h17 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h18 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h19 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h1a :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h1b :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h1c :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h1d :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h1e :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h1f :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h20 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h21 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h22 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h23 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h24 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h25 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h26 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h27 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h28 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h29 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h2a :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h2b :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h2c :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h2d :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h2e :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h2f :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h30 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h31 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h32 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h33 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h34 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h35 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h36 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h37 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h38 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h39 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h3a :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h3b :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h3c :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h3d :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h3e :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h3f :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h40 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h41 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h42 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h43 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h44 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h45 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h46 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h47 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h48 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h49 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h4a :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h4b :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h4c :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h4d :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h4e :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h4f :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h50 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h51 :
		TR_93 = 9'h000 ;	// line#=../rle.cpp:79
	7'h52 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h53 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h54 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h55 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h56 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h57 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h58 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h59 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h5a :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h5b :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h5c :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h5d :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h5e :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h5f :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h60 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h61 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h62 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h63 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h64 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h65 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h66 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h67 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h68 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h69 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h6a :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h6b :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h6c :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h6d :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h6e :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h6f :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h70 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h71 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h72 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h73 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h74 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h75 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h76 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h77 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h78 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h79 :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h7a :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h7b :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h7c :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h7d :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h7e :
		TR_93 = RG_quantized_block_rl_38 ;
	7'h7f :
		TR_93 = RG_quantized_block_rl_38 ;
	default :
		TR_93 = 9'hx ;
	endcase
always @ ( RG_rl_170 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_94 = RG_rl_170 ;
	7'h01 :
		TR_94 = RG_rl_170 ;
	7'h02 :
		TR_94 = RG_rl_170 ;
	7'h03 :
		TR_94 = RG_rl_170 ;
	7'h04 :
		TR_94 = RG_rl_170 ;
	7'h05 :
		TR_94 = RG_rl_170 ;
	7'h06 :
		TR_94 = RG_rl_170 ;
	7'h07 :
		TR_94 = RG_rl_170 ;
	7'h08 :
		TR_94 = RG_rl_170 ;
	7'h09 :
		TR_94 = RG_rl_170 ;
	7'h0a :
		TR_94 = RG_rl_170 ;
	7'h0b :
		TR_94 = RG_rl_170 ;
	7'h0c :
		TR_94 = RG_rl_170 ;
	7'h0d :
		TR_94 = RG_rl_170 ;
	7'h0e :
		TR_94 = RG_rl_170 ;
	7'h0f :
		TR_94 = RG_rl_170 ;
	7'h10 :
		TR_94 = RG_rl_170 ;
	7'h11 :
		TR_94 = RG_rl_170 ;
	7'h12 :
		TR_94 = RG_rl_170 ;
	7'h13 :
		TR_94 = RG_rl_170 ;
	7'h14 :
		TR_94 = RG_rl_170 ;
	7'h15 :
		TR_94 = RG_rl_170 ;
	7'h16 :
		TR_94 = RG_rl_170 ;
	7'h17 :
		TR_94 = RG_rl_170 ;
	7'h18 :
		TR_94 = RG_rl_170 ;
	7'h19 :
		TR_94 = RG_rl_170 ;
	7'h1a :
		TR_94 = RG_rl_170 ;
	7'h1b :
		TR_94 = RG_rl_170 ;
	7'h1c :
		TR_94 = RG_rl_170 ;
	7'h1d :
		TR_94 = RG_rl_170 ;
	7'h1e :
		TR_94 = RG_rl_170 ;
	7'h1f :
		TR_94 = RG_rl_170 ;
	7'h20 :
		TR_94 = RG_rl_170 ;
	7'h21 :
		TR_94 = RG_rl_170 ;
	7'h22 :
		TR_94 = RG_rl_170 ;
	7'h23 :
		TR_94 = RG_rl_170 ;
	7'h24 :
		TR_94 = RG_rl_170 ;
	7'h25 :
		TR_94 = RG_rl_170 ;
	7'h26 :
		TR_94 = RG_rl_170 ;
	7'h27 :
		TR_94 = RG_rl_170 ;
	7'h28 :
		TR_94 = RG_rl_170 ;
	7'h29 :
		TR_94 = RG_rl_170 ;
	7'h2a :
		TR_94 = RG_rl_170 ;
	7'h2b :
		TR_94 = RG_rl_170 ;
	7'h2c :
		TR_94 = RG_rl_170 ;
	7'h2d :
		TR_94 = RG_rl_170 ;
	7'h2e :
		TR_94 = RG_rl_170 ;
	7'h2f :
		TR_94 = RG_rl_170 ;
	7'h30 :
		TR_94 = RG_rl_170 ;
	7'h31 :
		TR_94 = RG_rl_170 ;
	7'h32 :
		TR_94 = RG_rl_170 ;
	7'h33 :
		TR_94 = RG_rl_170 ;
	7'h34 :
		TR_94 = RG_rl_170 ;
	7'h35 :
		TR_94 = RG_rl_170 ;
	7'h36 :
		TR_94 = RG_rl_170 ;
	7'h37 :
		TR_94 = RG_rl_170 ;
	7'h38 :
		TR_94 = RG_rl_170 ;
	7'h39 :
		TR_94 = RG_rl_170 ;
	7'h3a :
		TR_94 = RG_rl_170 ;
	7'h3b :
		TR_94 = RG_rl_170 ;
	7'h3c :
		TR_94 = RG_rl_170 ;
	7'h3d :
		TR_94 = RG_rl_170 ;
	7'h3e :
		TR_94 = RG_rl_170 ;
	7'h3f :
		TR_94 = RG_rl_170 ;
	7'h40 :
		TR_94 = RG_rl_170 ;
	7'h41 :
		TR_94 = RG_rl_170 ;
	7'h42 :
		TR_94 = RG_rl_170 ;
	7'h43 :
		TR_94 = RG_rl_170 ;
	7'h44 :
		TR_94 = RG_rl_170 ;
	7'h45 :
		TR_94 = RG_rl_170 ;
	7'h46 :
		TR_94 = RG_rl_170 ;
	7'h47 :
		TR_94 = RG_rl_170 ;
	7'h48 :
		TR_94 = RG_rl_170 ;
	7'h49 :
		TR_94 = RG_rl_170 ;
	7'h4a :
		TR_94 = RG_rl_170 ;
	7'h4b :
		TR_94 = RG_rl_170 ;
	7'h4c :
		TR_94 = RG_rl_170 ;
	7'h4d :
		TR_94 = RG_rl_170 ;
	7'h4e :
		TR_94 = RG_rl_170 ;
	7'h4f :
		TR_94 = RG_rl_170 ;
	7'h50 :
		TR_94 = RG_rl_170 ;
	7'h51 :
		TR_94 = RG_rl_170 ;
	7'h52 :
		TR_94 = 9'h000 ;	// line#=../rle.cpp:79
	7'h53 :
		TR_94 = RG_rl_170 ;
	7'h54 :
		TR_94 = RG_rl_170 ;
	7'h55 :
		TR_94 = RG_rl_170 ;
	7'h56 :
		TR_94 = RG_rl_170 ;
	7'h57 :
		TR_94 = RG_rl_170 ;
	7'h58 :
		TR_94 = RG_rl_170 ;
	7'h59 :
		TR_94 = RG_rl_170 ;
	7'h5a :
		TR_94 = RG_rl_170 ;
	7'h5b :
		TR_94 = RG_rl_170 ;
	7'h5c :
		TR_94 = RG_rl_170 ;
	7'h5d :
		TR_94 = RG_rl_170 ;
	7'h5e :
		TR_94 = RG_rl_170 ;
	7'h5f :
		TR_94 = RG_rl_170 ;
	7'h60 :
		TR_94 = RG_rl_170 ;
	7'h61 :
		TR_94 = RG_rl_170 ;
	7'h62 :
		TR_94 = RG_rl_170 ;
	7'h63 :
		TR_94 = RG_rl_170 ;
	7'h64 :
		TR_94 = RG_rl_170 ;
	7'h65 :
		TR_94 = RG_rl_170 ;
	7'h66 :
		TR_94 = RG_rl_170 ;
	7'h67 :
		TR_94 = RG_rl_170 ;
	7'h68 :
		TR_94 = RG_rl_170 ;
	7'h69 :
		TR_94 = RG_rl_170 ;
	7'h6a :
		TR_94 = RG_rl_170 ;
	7'h6b :
		TR_94 = RG_rl_170 ;
	7'h6c :
		TR_94 = RG_rl_170 ;
	7'h6d :
		TR_94 = RG_rl_170 ;
	7'h6e :
		TR_94 = RG_rl_170 ;
	7'h6f :
		TR_94 = RG_rl_170 ;
	7'h70 :
		TR_94 = RG_rl_170 ;
	7'h71 :
		TR_94 = RG_rl_170 ;
	7'h72 :
		TR_94 = RG_rl_170 ;
	7'h73 :
		TR_94 = RG_rl_170 ;
	7'h74 :
		TR_94 = RG_rl_170 ;
	7'h75 :
		TR_94 = RG_rl_170 ;
	7'h76 :
		TR_94 = RG_rl_170 ;
	7'h77 :
		TR_94 = RG_rl_170 ;
	7'h78 :
		TR_94 = RG_rl_170 ;
	7'h79 :
		TR_94 = RG_rl_170 ;
	7'h7a :
		TR_94 = RG_rl_170 ;
	7'h7b :
		TR_94 = RG_rl_170 ;
	7'h7c :
		TR_94 = RG_rl_170 ;
	7'h7d :
		TR_94 = RG_rl_170 ;
	7'h7e :
		TR_94 = RG_rl_170 ;
	7'h7f :
		TR_94 = RG_rl_170 ;
	default :
		TR_94 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_39 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h01 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h02 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h03 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h04 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h05 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h06 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h07 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h08 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h09 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h0a :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h0b :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h0c :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h0d :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h0e :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h0f :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h10 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h11 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h12 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h13 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h14 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h15 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h16 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h17 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h18 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h19 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h1a :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h1b :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h1c :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h1d :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h1e :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h1f :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h20 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h21 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h22 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h23 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h24 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h25 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h26 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h27 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h28 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h29 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h2a :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h2b :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h2c :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h2d :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h2e :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h2f :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h30 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h31 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h32 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h33 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h34 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h35 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h36 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h37 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h38 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h39 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h3a :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h3b :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h3c :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h3d :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h3e :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h3f :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h40 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h41 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h42 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h43 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h44 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h45 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h46 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h47 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h48 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h49 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h4a :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h4b :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h4c :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h4d :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h4e :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h4f :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h50 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h51 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h52 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h53 :
		TR_95 = 9'h000 ;	// line#=../rle.cpp:79
	7'h54 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h55 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h56 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h57 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h58 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h59 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h5a :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h5b :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h5c :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h5d :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h5e :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h5f :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h60 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h61 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h62 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h63 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h64 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h65 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h66 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h67 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h68 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h69 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h6a :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h6b :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h6c :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h6d :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h6e :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h6f :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h70 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h71 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h72 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h73 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h74 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h75 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h76 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h77 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h78 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h79 :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h7a :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h7b :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h7c :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h7d :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h7e :
		TR_95 = RG_quantized_block_rl_39 ;
	7'h7f :
		TR_95 = RG_quantized_block_rl_39 ;
	default :
		TR_95 = 9'hx ;
	endcase
always @ ( RG_rl_171 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_96 = RG_rl_171 ;
	7'h01 :
		TR_96 = RG_rl_171 ;
	7'h02 :
		TR_96 = RG_rl_171 ;
	7'h03 :
		TR_96 = RG_rl_171 ;
	7'h04 :
		TR_96 = RG_rl_171 ;
	7'h05 :
		TR_96 = RG_rl_171 ;
	7'h06 :
		TR_96 = RG_rl_171 ;
	7'h07 :
		TR_96 = RG_rl_171 ;
	7'h08 :
		TR_96 = RG_rl_171 ;
	7'h09 :
		TR_96 = RG_rl_171 ;
	7'h0a :
		TR_96 = RG_rl_171 ;
	7'h0b :
		TR_96 = RG_rl_171 ;
	7'h0c :
		TR_96 = RG_rl_171 ;
	7'h0d :
		TR_96 = RG_rl_171 ;
	7'h0e :
		TR_96 = RG_rl_171 ;
	7'h0f :
		TR_96 = RG_rl_171 ;
	7'h10 :
		TR_96 = RG_rl_171 ;
	7'h11 :
		TR_96 = RG_rl_171 ;
	7'h12 :
		TR_96 = RG_rl_171 ;
	7'h13 :
		TR_96 = RG_rl_171 ;
	7'h14 :
		TR_96 = RG_rl_171 ;
	7'h15 :
		TR_96 = RG_rl_171 ;
	7'h16 :
		TR_96 = RG_rl_171 ;
	7'h17 :
		TR_96 = RG_rl_171 ;
	7'h18 :
		TR_96 = RG_rl_171 ;
	7'h19 :
		TR_96 = RG_rl_171 ;
	7'h1a :
		TR_96 = RG_rl_171 ;
	7'h1b :
		TR_96 = RG_rl_171 ;
	7'h1c :
		TR_96 = RG_rl_171 ;
	7'h1d :
		TR_96 = RG_rl_171 ;
	7'h1e :
		TR_96 = RG_rl_171 ;
	7'h1f :
		TR_96 = RG_rl_171 ;
	7'h20 :
		TR_96 = RG_rl_171 ;
	7'h21 :
		TR_96 = RG_rl_171 ;
	7'h22 :
		TR_96 = RG_rl_171 ;
	7'h23 :
		TR_96 = RG_rl_171 ;
	7'h24 :
		TR_96 = RG_rl_171 ;
	7'h25 :
		TR_96 = RG_rl_171 ;
	7'h26 :
		TR_96 = RG_rl_171 ;
	7'h27 :
		TR_96 = RG_rl_171 ;
	7'h28 :
		TR_96 = RG_rl_171 ;
	7'h29 :
		TR_96 = RG_rl_171 ;
	7'h2a :
		TR_96 = RG_rl_171 ;
	7'h2b :
		TR_96 = RG_rl_171 ;
	7'h2c :
		TR_96 = RG_rl_171 ;
	7'h2d :
		TR_96 = RG_rl_171 ;
	7'h2e :
		TR_96 = RG_rl_171 ;
	7'h2f :
		TR_96 = RG_rl_171 ;
	7'h30 :
		TR_96 = RG_rl_171 ;
	7'h31 :
		TR_96 = RG_rl_171 ;
	7'h32 :
		TR_96 = RG_rl_171 ;
	7'h33 :
		TR_96 = RG_rl_171 ;
	7'h34 :
		TR_96 = RG_rl_171 ;
	7'h35 :
		TR_96 = RG_rl_171 ;
	7'h36 :
		TR_96 = RG_rl_171 ;
	7'h37 :
		TR_96 = RG_rl_171 ;
	7'h38 :
		TR_96 = RG_rl_171 ;
	7'h39 :
		TR_96 = RG_rl_171 ;
	7'h3a :
		TR_96 = RG_rl_171 ;
	7'h3b :
		TR_96 = RG_rl_171 ;
	7'h3c :
		TR_96 = RG_rl_171 ;
	7'h3d :
		TR_96 = RG_rl_171 ;
	7'h3e :
		TR_96 = RG_rl_171 ;
	7'h3f :
		TR_96 = RG_rl_171 ;
	7'h40 :
		TR_96 = RG_rl_171 ;
	7'h41 :
		TR_96 = RG_rl_171 ;
	7'h42 :
		TR_96 = RG_rl_171 ;
	7'h43 :
		TR_96 = RG_rl_171 ;
	7'h44 :
		TR_96 = RG_rl_171 ;
	7'h45 :
		TR_96 = RG_rl_171 ;
	7'h46 :
		TR_96 = RG_rl_171 ;
	7'h47 :
		TR_96 = RG_rl_171 ;
	7'h48 :
		TR_96 = RG_rl_171 ;
	7'h49 :
		TR_96 = RG_rl_171 ;
	7'h4a :
		TR_96 = RG_rl_171 ;
	7'h4b :
		TR_96 = RG_rl_171 ;
	7'h4c :
		TR_96 = RG_rl_171 ;
	7'h4d :
		TR_96 = RG_rl_171 ;
	7'h4e :
		TR_96 = RG_rl_171 ;
	7'h4f :
		TR_96 = RG_rl_171 ;
	7'h50 :
		TR_96 = RG_rl_171 ;
	7'h51 :
		TR_96 = RG_rl_171 ;
	7'h52 :
		TR_96 = RG_rl_171 ;
	7'h53 :
		TR_96 = RG_rl_171 ;
	7'h54 :
		TR_96 = 9'h000 ;	// line#=../rle.cpp:79
	7'h55 :
		TR_96 = RG_rl_171 ;
	7'h56 :
		TR_96 = RG_rl_171 ;
	7'h57 :
		TR_96 = RG_rl_171 ;
	7'h58 :
		TR_96 = RG_rl_171 ;
	7'h59 :
		TR_96 = RG_rl_171 ;
	7'h5a :
		TR_96 = RG_rl_171 ;
	7'h5b :
		TR_96 = RG_rl_171 ;
	7'h5c :
		TR_96 = RG_rl_171 ;
	7'h5d :
		TR_96 = RG_rl_171 ;
	7'h5e :
		TR_96 = RG_rl_171 ;
	7'h5f :
		TR_96 = RG_rl_171 ;
	7'h60 :
		TR_96 = RG_rl_171 ;
	7'h61 :
		TR_96 = RG_rl_171 ;
	7'h62 :
		TR_96 = RG_rl_171 ;
	7'h63 :
		TR_96 = RG_rl_171 ;
	7'h64 :
		TR_96 = RG_rl_171 ;
	7'h65 :
		TR_96 = RG_rl_171 ;
	7'h66 :
		TR_96 = RG_rl_171 ;
	7'h67 :
		TR_96 = RG_rl_171 ;
	7'h68 :
		TR_96 = RG_rl_171 ;
	7'h69 :
		TR_96 = RG_rl_171 ;
	7'h6a :
		TR_96 = RG_rl_171 ;
	7'h6b :
		TR_96 = RG_rl_171 ;
	7'h6c :
		TR_96 = RG_rl_171 ;
	7'h6d :
		TR_96 = RG_rl_171 ;
	7'h6e :
		TR_96 = RG_rl_171 ;
	7'h6f :
		TR_96 = RG_rl_171 ;
	7'h70 :
		TR_96 = RG_rl_171 ;
	7'h71 :
		TR_96 = RG_rl_171 ;
	7'h72 :
		TR_96 = RG_rl_171 ;
	7'h73 :
		TR_96 = RG_rl_171 ;
	7'h74 :
		TR_96 = RG_rl_171 ;
	7'h75 :
		TR_96 = RG_rl_171 ;
	7'h76 :
		TR_96 = RG_rl_171 ;
	7'h77 :
		TR_96 = RG_rl_171 ;
	7'h78 :
		TR_96 = RG_rl_171 ;
	7'h79 :
		TR_96 = RG_rl_171 ;
	7'h7a :
		TR_96 = RG_rl_171 ;
	7'h7b :
		TR_96 = RG_rl_171 ;
	7'h7c :
		TR_96 = RG_rl_171 ;
	7'h7d :
		TR_96 = RG_rl_171 ;
	7'h7e :
		TR_96 = RG_rl_171 ;
	7'h7f :
		TR_96 = RG_rl_171 ;
	default :
		TR_96 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_40 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h01 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h02 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h03 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h04 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h05 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h06 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h07 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h08 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h09 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h0a :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h0b :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h0c :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h0d :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h0e :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h0f :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h10 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h11 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h12 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h13 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h14 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h15 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h16 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h17 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h18 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h19 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h1a :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h1b :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h1c :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h1d :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h1e :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h1f :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h20 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h21 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h22 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h23 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h24 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h25 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h26 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h27 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h28 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h29 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h2a :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h2b :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h2c :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h2d :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h2e :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h2f :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h30 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h31 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h32 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h33 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h34 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h35 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h36 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h37 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h38 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h39 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h3a :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h3b :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h3c :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h3d :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h3e :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h3f :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h40 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h41 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h42 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h43 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h44 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h45 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h46 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h47 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h48 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h49 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h4a :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h4b :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h4c :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h4d :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h4e :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h4f :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h50 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h51 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h52 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h53 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h54 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h55 :
		TR_97 = 9'h000 ;	// line#=../rle.cpp:79
	7'h56 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h57 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h58 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h59 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h5a :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h5b :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h5c :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h5d :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h5e :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h5f :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h60 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h61 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h62 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h63 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h64 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h65 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h66 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h67 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h68 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h69 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h6a :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h6b :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h6c :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h6d :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h6e :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h6f :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h70 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h71 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h72 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h73 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h74 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h75 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h76 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h77 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h78 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h79 :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h7a :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h7b :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h7c :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h7d :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h7e :
		TR_97 = RG_quantized_block_rl_40 ;
	7'h7f :
		TR_97 = RG_quantized_block_rl_40 ;
	default :
		TR_97 = 9'hx ;
	endcase
always @ ( RG_rl_172 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_98 = RG_rl_172 ;
	7'h01 :
		TR_98 = RG_rl_172 ;
	7'h02 :
		TR_98 = RG_rl_172 ;
	7'h03 :
		TR_98 = RG_rl_172 ;
	7'h04 :
		TR_98 = RG_rl_172 ;
	7'h05 :
		TR_98 = RG_rl_172 ;
	7'h06 :
		TR_98 = RG_rl_172 ;
	7'h07 :
		TR_98 = RG_rl_172 ;
	7'h08 :
		TR_98 = RG_rl_172 ;
	7'h09 :
		TR_98 = RG_rl_172 ;
	7'h0a :
		TR_98 = RG_rl_172 ;
	7'h0b :
		TR_98 = RG_rl_172 ;
	7'h0c :
		TR_98 = RG_rl_172 ;
	7'h0d :
		TR_98 = RG_rl_172 ;
	7'h0e :
		TR_98 = RG_rl_172 ;
	7'h0f :
		TR_98 = RG_rl_172 ;
	7'h10 :
		TR_98 = RG_rl_172 ;
	7'h11 :
		TR_98 = RG_rl_172 ;
	7'h12 :
		TR_98 = RG_rl_172 ;
	7'h13 :
		TR_98 = RG_rl_172 ;
	7'h14 :
		TR_98 = RG_rl_172 ;
	7'h15 :
		TR_98 = RG_rl_172 ;
	7'h16 :
		TR_98 = RG_rl_172 ;
	7'h17 :
		TR_98 = RG_rl_172 ;
	7'h18 :
		TR_98 = RG_rl_172 ;
	7'h19 :
		TR_98 = RG_rl_172 ;
	7'h1a :
		TR_98 = RG_rl_172 ;
	7'h1b :
		TR_98 = RG_rl_172 ;
	7'h1c :
		TR_98 = RG_rl_172 ;
	7'h1d :
		TR_98 = RG_rl_172 ;
	7'h1e :
		TR_98 = RG_rl_172 ;
	7'h1f :
		TR_98 = RG_rl_172 ;
	7'h20 :
		TR_98 = RG_rl_172 ;
	7'h21 :
		TR_98 = RG_rl_172 ;
	7'h22 :
		TR_98 = RG_rl_172 ;
	7'h23 :
		TR_98 = RG_rl_172 ;
	7'h24 :
		TR_98 = RG_rl_172 ;
	7'h25 :
		TR_98 = RG_rl_172 ;
	7'h26 :
		TR_98 = RG_rl_172 ;
	7'h27 :
		TR_98 = RG_rl_172 ;
	7'h28 :
		TR_98 = RG_rl_172 ;
	7'h29 :
		TR_98 = RG_rl_172 ;
	7'h2a :
		TR_98 = RG_rl_172 ;
	7'h2b :
		TR_98 = RG_rl_172 ;
	7'h2c :
		TR_98 = RG_rl_172 ;
	7'h2d :
		TR_98 = RG_rl_172 ;
	7'h2e :
		TR_98 = RG_rl_172 ;
	7'h2f :
		TR_98 = RG_rl_172 ;
	7'h30 :
		TR_98 = RG_rl_172 ;
	7'h31 :
		TR_98 = RG_rl_172 ;
	7'h32 :
		TR_98 = RG_rl_172 ;
	7'h33 :
		TR_98 = RG_rl_172 ;
	7'h34 :
		TR_98 = RG_rl_172 ;
	7'h35 :
		TR_98 = RG_rl_172 ;
	7'h36 :
		TR_98 = RG_rl_172 ;
	7'h37 :
		TR_98 = RG_rl_172 ;
	7'h38 :
		TR_98 = RG_rl_172 ;
	7'h39 :
		TR_98 = RG_rl_172 ;
	7'h3a :
		TR_98 = RG_rl_172 ;
	7'h3b :
		TR_98 = RG_rl_172 ;
	7'h3c :
		TR_98 = RG_rl_172 ;
	7'h3d :
		TR_98 = RG_rl_172 ;
	7'h3e :
		TR_98 = RG_rl_172 ;
	7'h3f :
		TR_98 = RG_rl_172 ;
	7'h40 :
		TR_98 = RG_rl_172 ;
	7'h41 :
		TR_98 = RG_rl_172 ;
	7'h42 :
		TR_98 = RG_rl_172 ;
	7'h43 :
		TR_98 = RG_rl_172 ;
	7'h44 :
		TR_98 = RG_rl_172 ;
	7'h45 :
		TR_98 = RG_rl_172 ;
	7'h46 :
		TR_98 = RG_rl_172 ;
	7'h47 :
		TR_98 = RG_rl_172 ;
	7'h48 :
		TR_98 = RG_rl_172 ;
	7'h49 :
		TR_98 = RG_rl_172 ;
	7'h4a :
		TR_98 = RG_rl_172 ;
	7'h4b :
		TR_98 = RG_rl_172 ;
	7'h4c :
		TR_98 = RG_rl_172 ;
	7'h4d :
		TR_98 = RG_rl_172 ;
	7'h4e :
		TR_98 = RG_rl_172 ;
	7'h4f :
		TR_98 = RG_rl_172 ;
	7'h50 :
		TR_98 = RG_rl_172 ;
	7'h51 :
		TR_98 = RG_rl_172 ;
	7'h52 :
		TR_98 = RG_rl_172 ;
	7'h53 :
		TR_98 = RG_rl_172 ;
	7'h54 :
		TR_98 = RG_rl_172 ;
	7'h55 :
		TR_98 = RG_rl_172 ;
	7'h56 :
		TR_98 = 9'h000 ;	// line#=../rle.cpp:79
	7'h57 :
		TR_98 = RG_rl_172 ;
	7'h58 :
		TR_98 = RG_rl_172 ;
	7'h59 :
		TR_98 = RG_rl_172 ;
	7'h5a :
		TR_98 = RG_rl_172 ;
	7'h5b :
		TR_98 = RG_rl_172 ;
	7'h5c :
		TR_98 = RG_rl_172 ;
	7'h5d :
		TR_98 = RG_rl_172 ;
	7'h5e :
		TR_98 = RG_rl_172 ;
	7'h5f :
		TR_98 = RG_rl_172 ;
	7'h60 :
		TR_98 = RG_rl_172 ;
	7'h61 :
		TR_98 = RG_rl_172 ;
	7'h62 :
		TR_98 = RG_rl_172 ;
	7'h63 :
		TR_98 = RG_rl_172 ;
	7'h64 :
		TR_98 = RG_rl_172 ;
	7'h65 :
		TR_98 = RG_rl_172 ;
	7'h66 :
		TR_98 = RG_rl_172 ;
	7'h67 :
		TR_98 = RG_rl_172 ;
	7'h68 :
		TR_98 = RG_rl_172 ;
	7'h69 :
		TR_98 = RG_rl_172 ;
	7'h6a :
		TR_98 = RG_rl_172 ;
	7'h6b :
		TR_98 = RG_rl_172 ;
	7'h6c :
		TR_98 = RG_rl_172 ;
	7'h6d :
		TR_98 = RG_rl_172 ;
	7'h6e :
		TR_98 = RG_rl_172 ;
	7'h6f :
		TR_98 = RG_rl_172 ;
	7'h70 :
		TR_98 = RG_rl_172 ;
	7'h71 :
		TR_98 = RG_rl_172 ;
	7'h72 :
		TR_98 = RG_rl_172 ;
	7'h73 :
		TR_98 = RG_rl_172 ;
	7'h74 :
		TR_98 = RG_rl_172 ;
	7'h75 :
		TR_98 = RG_rl_172 ;
	7'h76 :
		TR_98 = RG_rl_172 ;
	7'h77 :
		TR_98 = RG_rl_172 ;
	7'h78 :
		TR_98 = RG_rl_172 ;
	7'h79 :
		TR_98 = RG_rl_172 ;
	7'h7a :
		TR_98 = RG_rl_172 ;
	7'h7b :
		TR_98 = RG_rl_172 ;
	7'h7c :
		TR_98 = RG_rl_172 ;
	7'h7d :
		TR_98 = RG_rl_172 ;
	7'h7e :
		TR_98 = RG_rl_172 ;
	7'h7f :
		TR_98 = RG_rl_172 ;
	default :
		TR_98 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_41 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h01 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h02 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h03 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h04 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h05 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h06 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h07 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h08 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h09 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h0a :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h0b :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h0c :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h0d :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h0e :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h0f :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h10 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h11 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h12 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h13 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h14 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h15 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h16 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h17 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h18 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h19 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h1a :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h1b :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h1c :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h1d :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h1e :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h1f :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h20 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h21 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h22 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h23 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h24 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h25 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h26 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h27 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h28 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h29 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h2a :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h2b :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h2c :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h2d :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h2e :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h2f :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h30 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h31 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h32 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h33 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h34 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h35 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h36 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h37 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h38 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h39 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h3a :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h3b :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h3c :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h3d :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h3e :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h3f :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h40 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h41 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h42 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h43 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h44 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h45 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h46 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h47 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h48 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h49 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h4a :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h4b :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h4c :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h4d :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h4e :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h4f :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h50 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h51 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h52 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h53 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h54 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h55 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h56 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h57 :
		TR_99 = 9'h000 ;	// line#=../rle.cpp:79
	7'h58 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h59 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h5a :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h5b :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h5c :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h5d :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h5e :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h5f :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h60 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h61 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h62 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h63 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h64 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h65 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h66 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h67 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h68 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h69 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h6a :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h6b :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h6c :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h6d :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h6e :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h6f :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h70 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h71 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h72 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h73 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h74 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h75 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h76 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h77 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h78 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h79 :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h7a :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h7b :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h7c :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h7d :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h7e :
		TR_99 = RG_quantized_block_rl_41 ;
	7'h7f :
		TR_99 = RG_quantized_block_rl_41 ;
	default :
		TR_99 = 9'hx ;
	endcase
always @ ( RG_rl_173 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_100 = RG_rl_173 ;
	7'h01 :
		TR_100 = RG_rl_173 ;
	7'h02 :
		TR_100 = RG_rl_173 ;
	7'h03 :
		TR_100 = RG_rl_173 ;
	7'h04 :
		TR_100 = RG_rl_173 ;
	7'h05 :
		TR_100 = RG_rl_173 ;
	7'h06 :
		TR_100 = RG_rl_173 ;
	7'h07 :
		TR_100 = RG_rl_173 ;
	7'h08 :
		TR_100 = RG_rl_173 ;
	7'h09 :
		TR_100 = RG_rl_173 ;
	7'h0a :
		TR_100 = RG_rl_173 ;
	7'h0b :
		TR_100 = RG_rl_173 ;
	7'h0c :
		TR_100 = RG_rl_173 ;
	7'h0d :
		TR_100 = RG_rl_173 ;
	7'h0e :
		TR_100 = RG_rl_173 ;
	7'h0f :
		TR_100 = RG_rl_173 ;
	7'h10 :
		TR_100 = RG_rl_173 ;
	7'h11 :
		TR_100 = RG_rl_173 ;
	7'h12 :
		TR_100 = RG_rl_173 ;
	7'h13 :
		TR_100 = RG_rl_173 ;
	7'h14 :
		TR_100 = RG_rl_173 ;
	7'h15 :
		TR_100 = RG_rl_173 ;
	7'h16 :
		TR_100 = RG_rl_173 ;
	7'h17 :
		TR_100 = RG_rl_173 ;
	7'h18 :
		TR_100 = RG_rl_173 ;
	7'h19 :
		TR_100 = RG_rl_173 ;
	7'h1a :
		TR_100 = RG_rl_173 ;
	7'h1b :
		TR_100 = RG_rl_173 ;
	7'h1c :
		TR_100 = RG_rl_173 ;
	7'h1d :
		TR_100 = RG_rl_173 ;
	7'h1e :
		TR_100 = RG_rl_173 ;
	7'h1f :
		TR_100 = RG_rl_173 ;
	7'h20 :
		TR_100 = RG_rl_173 ;
	7'h21 :
		TR_100 = RG_rl_173 ;
	7'h22 :
		TR_100 = RG_rl_173 ;
	7'h23 :
		TR_100 = RG_rl_173 ;
	7'h24 :
		TR_100 = RG_rl_173 ;
	7'h25 :
		TR_100 = RG_rl_173 ;
	7'h26 :
		TR_100 = RG_rl_173 ;
	7'h27 :
		TR_100 = RG_rl_173 ;
	7'h28 :
		TR_100 = RG_rl_173 ;
	7'h29 :
		TR_100 = RG_rl_173 ;
	7'h2a :
		TR_100 = RG_rl_173 ;
	7'h2b :
		TR_100 = RG_rl_173 ;
	7'h2c :
		TR_100 = RG_rl_173 ;
	7'h2d :
		TR_100 = RG_rl_173 ;
	7'h2e :
		TR_100 = RG_rl_173 ;
	7'h2f :
		TR_100 = RG_rl_173 ;
	7'h30 :
		TR_100 = RG_rl_173 ;
	7'h31 :
		TR_100 = RG_rl_173 ;
	7'h32 :
		TR_100 = RG_rl_173 ;
	7'h33 :
		TR_100 = RG_rl_173 ;
	7'h34 :
		TR_100 = RG_rl_173 ;
	7'h35 :
		TR_100 = RG_rl_173 ;
	7'h36 :
		TR_100 = RG_rl_173 ;
	7'h37 :
		TR_100 = RG_rl_173 ;
	7'h38 :
		TR_100 = RG_rl_173 ;
	7'h39 :
		TR_100 = RG_rl_173 ;
	7'h3a :
		TR_100 = RG_rl_173 ;
	7'h3b :
		TR_100 = RG_rl_173 ;
	7'h3c :
		TR_100 = RG_rl_173 ;
	7'h3d :
		TR_100 = RG_rl_173 ;
	7'h3e :
		TR_100 = RG_rl_173 ;
	7'h3f :
		TR_100 = RG_rl_173 ;
	7'h40 :
		TR_100 = RG_rl_173 ;
	7'h41 :
		TR_100 = RG_rl_173 ;
	7'h42 :
		TR_100 = RG_rl_173 ;
	7'h43 :
		TR_100 = RG_rl_173 ;
	7'h44 :
		TR_100 = RG_rl_173 ;
	7'h45 :
		TR_100 = RG_rl_173 ;
	7'h46 :
		TR_100 = RG_rl_173 ;
	7'h47 :
		TR_100 = RG_rl_173 ;
	7'h48 :
		TR_100 = RG_rl_173 ;
	7'h49 :
		TR_100 = RG_rl_173 ;
	7'h4a :
		TR_100 = RG_rl_173 ;
	7'h4b :
		TR_100 = RG_rl_173 ;
	7'h4c :
		TR_100 = RG_rl_173 ;
	7'h4d :
		TR_100 = RG_rl_173 ;
	7'h4e :
		TR_100 = RG_rl_173 ;
	7'h4f :
		TR_100 = RG_rl_173 ;
	7'h50 :
		TR_100 = RG_rl_173 ;
	7'h51 :
		TR_100 = RG_rl_173 ;
	7'h52 :
		TR_100 = RG_rl_173 ;
	7'h53 :
		TR_100 = RG_rl_173 ;
	7'h54 :
		TR_100 = RG_rl_173 ;
	7'h55 :
		TR_100 = RG_rl_173 ;
	7'h56 :
		TR_100 = RG_rl_173 ;
	7'h57 :
		TR_100 = RG_rl_173 ;
	7'h58 :
		TR_100 = 9'h000 ;	// line#=../rle.cpp:79
	7'h59 :
		TR_100 = RG_rl_173 ;
	7'h5a :
		TR_100 = RG_rl_173 ;
	7'h5b :
		TR_100 = RG_rl_173 ;
	7'h5c :
		TR_100 = RG_rl_173 ;
	7'h5d :
		TR_100 = RG_rl_173 ;
	7'h5e :
		TR_100 = RG_rl_173 ;
	7'h5f :
		TR_100 = RG_rl_173 ;
	7'h60 :
		TR_100 = RG_rl_173 ;
	7'h61 :
		TR_100 = RG_rl_173 ;
	7'h62 :
		TR_100 = RG_rl_173 ;
	7'h63 :
		TR_100 = RG_rl_173 ;
	7'h64 :
		TR_100 = RG_rl_173 ;
	7'h65 :
		TR_100 = RG_rl_173 ;
	7'h66 :
		TR_100 = RG_rl_173 ;
	7'h67 :
		TR_100 = RG_rl_173 ;
	7'h68 :
		TR_100 = RG_rl_173 ;
	7'h69 :
		TR_100 = RG_rl_173 ;
	7'h6a :
		TR_100 = RG_rl_173 ;
	7'h6b :
		TR_100 = RG_rl_173 ;
	7'h6c :
		TR_100 = RG_rl_173 ;
	7'h6d :
		TR_100 = RG_rl_173 ;
	7'h6e :
		TR_100 = RG_rl_173 ;
	7'h6f :
		TR_100 = RG_rl_173 ;
	7'h70 :
		TR_100 = RG_rl_173 ;
	7'h71 :
		TR_100 = RG_rl_173 ;
	7'h72 :
		TR_100 = RG_rl_173 ;
	7'h73 :
		TR_100 = RG_rl_173 ;
	7'h74 :
		TR_100 = RG_rl_173 ;
	7'h75 :
		TR_100 = RG_rl_173 ;
	7'h76 :
		TR_100 = RG_rl_173 ;
	7'h77 :
		TR_100 = RG_rl_173 ;
	7'h78 :
		TR_100 = RG_rl_173 ;
	7'h79 :
		TR_100 = RG_rl_173 ;
	7'h7a :
		TR_100 = RG_rl_173 ;
	7'h7b :
		TR_100 = RG_rl_173 ;
	7'h7c :
		TR_100 = RG_rl_173 ;
	7'h7d :
		TR_100 = RG_rl_173 ;
	7'h7e :
		TR_100 = RG_rl_173 ;
	7'h7f :
		TR_100 = RG_rl_173 ;
	default :
		TR_100 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_42 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h01 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h02 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h03 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h04 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h05 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h06 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h07 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h08 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h09 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h0a :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h0b :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h0c :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h0d :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h0e :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h0f :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h10 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h11 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h12 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h13 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h14 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h15 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h16 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h17 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h18 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h19 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h1a :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h1b :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h1c :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h1d :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h1e :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h1f :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h20 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h21 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h22 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h23 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h24 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h25 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h26 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h27 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h28 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h29 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h2a :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h2b :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h2c :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h2d :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h2e :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h2f :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h30 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h31 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h32 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h33 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h34 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h35 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h36 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h37 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h38 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h39 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h3a :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h3b :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h3c :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h3d :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h3e :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h3f :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h40 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h41 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h42 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h43 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h44 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h45 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h46 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h47 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h48 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h49 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h4a :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h4b :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h4c :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h4d :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h4e :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h4f :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h50 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h51 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h52 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h53 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h54 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h55 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h56 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h57 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h58 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h59 :
		TR_101 = 9'h000 ;	// line#=../rle.cpp:79
	7'h5a :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h5b :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h5c :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h5d :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h5e :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h5f :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h60 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h61 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h62 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h63 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h64 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h65 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h66 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h67 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h68 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h69 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h6a :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h6b :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h6c :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h6d :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h6e :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h6f :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h70 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h71 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h72 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h73 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h74 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h75 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h76 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h77 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h78 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h79 :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h7a :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h7b :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h7c :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h7d :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h7e :
		TR_101 = RG_quantized_block_rl_42 ;
	7'h7f :
		TR_101 = RG_quantized_block_rl_42 ;
	default :
		TR_101 = 9'hx ;
	endcase
always @ ( RG_rl_174 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_102 = RG_rl_174 ;
	7'h01 :
		TR_102 = RG_rl_174 ;
	7'h02 :
		TR_102 = RG_rl_174 ;
	7'h03 :
		TR_102 = RG_rl_174 ;
	7'h04 :
		TR_102 = RG_rl_174 ;
	7'h05 :
		TR_102 = RG_rl_174 ;
	7'h06 :
		TR_102 = RG_rl_174 ;
	7'h07 :
		TR_102 = RG_rl_174 ;
	7'h08 :
		TR_102 = RG_rl_174 ;
	7'h09 :
		TR_102 = RG_rl_174 ;
	7'h0a :
		TR_102 = RG_rl_174 ;
	7'h0b :
		TR_102 = RG_rl_174 ;
	7'h0c :
		TR_102 = RG_rl_174 ;
	7'h0d :
		TR_102 = RG_rl_174 ;
	7'h0e :
		TR_102 = RG_rl_174 ;
	7'h0f :
		TR_102 = RG_rl_174 ;
	7'h10 :
		TR_102 = RG_rl_174 ;
	7'h11 :
		TR_102 = RG_rl_174 ;
	7'h12 :
		TR_102 = RG_rl_174 ;
	7'h13 :
		TR_102 = RG_rl_174 ;
	7'h14 :
		TR_102 = RG_rl_174 ;
	7'h15 :
		TR_102 = RG_rl_174 ;
	7'h16 :
		TR_102 = RG_rl_174 ;
	7'h17 :
		TR_102 = RG_rl_174 ;
	7'h18 :
		TR_102 = RG_rl_174 ;
	7'h19 :
		TR_102 = RG_rl_174 ;
	7'h1a :
		TR_102 = RG_rl_174 ;
	7'h1b :
		TR_102 = RG_rl_174 ;
	7'h1c :
		TR_102 = RG_rl_174 ;
	7'h1d :
		TR_102 = RG_rl_174 ;
	7'h1e :
		TR_102 = RG_rl_174 ;
	7'h1f :
		TR_102 = RG_rl_174 ;
	7'h20 :
		TR_102 = RG_rl_174 ;
	7'h21 :
		TR_102 = RG_rl_174 ;
	7'h22 :
		TR_102 = RG_rl_174 ;
	7'h23 :
		TR_102 = RG_rl_174 ;
	7'h24 :
		TR_102 = RG_rl_174 ;
	7'h25 :
		TR_102 = RG_rl_174 ;
	7'h26 :
		TR_102 = RG_rl_174 ;
	7'h27 :
		TR_102 = RG_rl_174 ;
	7'h28 :
		TR_102 = RG_rl_174 ;
	7'h29 :
		TR_102 = RG_rl_174 ;
	7'h2a :
		TR_102 = RG_rl_174 ;
	7'h2b :
		TR_102 = RG_rl_174 ;
	7'h2c :
		TR_102 = RG_rl_174 ;
	7'h2d :
		TR_102 = RG_rl_174 ;
	7'h2e :
		TR_102 = RG_rl_174 ;
	7'h2f :
		TR_102 = RG_rl_174 ;
	7'h30 :
		TR_102 = RG_rl_174 ;
	7'h31 :
		TR_102 = RG_rl_174 ;
	7'h32 :
		TR_102 = RG_rl_174 ;
	7'h33 :
		TR_102 = RG_rl_174 ;
	7'h34 :
		TR_102 = RG_rl_174 ;
	7'h35 :
		TR_102 = RG_rl_174 ;
	7'h36 :
		TR_102 = RG_rl_174 ;
	7'h37 :
		TR_102 = RG_rl_174 ;
	7'h38 :
		TR_102 = RG_rl_174 ;
	7'h39 :
		TR_102 = RG_rl_174 ;
	7'h3a :
		TR_102 = RG_rl_174 ;
	7'h3b :
		TR_102 = RG_rl_174 ;
	7'h3c :
		TR_102 = RG_rl_174 ;
	7'h3d :
		TR_102 = RG_rl_174 ;
	7'h3e :
		TR_102 = RG_rl_174 ;
	7'h3f :
		TR_102 = RG_rl_174 ;
	7'h40 :
		TR_102 = RG_rl_174 ;
	7'h41 :
		TR_102 = RG_rl_174 ;
	7'h42 :
		TR_102 = RG_rl_174 ;
	7'h43 :
		TR_102 = RG_rl_174 ;
	7'h44 :
		TR_102 = RG_rl_174 ;
	7'h45 :
		TR_102 = RG_rl_174 ;
	7'h46 :
		TR_102 = RG_rl_174 ;
	7'h47 :
		TR_102 = RG_rl_174 ;
	7'h48 :
		TR_102 = RG_rl_174 ;
	7'h49 :
		TR_102 = RG_rl_174 ;
	7'h4a :
		TR_102 = RG_rl_174 ;
	7'h4b :
		TR_102 = RG_rl_174 ;
	7'h4c :
		TR_102 = RG_rl_174 ;
	7'h4d :
		TR_102 = RG_rl_174 ;
	7'h4e :
		TR_102 = RG_rl_174 ;
	7'h4f :
		TR_102 = RG_rl_174 ;
	7'h50 :
		TR_102 = RG_rl_174 ;
	7'h51 :
		TR_102 = RG_rl_174 ;
	7'h52 :
		TR_102 = RG_rl_174 ;
	7'h53 :
		TR_102 = RG_rl_174 ;
	7'h54 :
		TR_102 = RG_rl_174 ;
	7'h55 :
		TR_102 = RG_rl_174 ;
	7'h56 :
		TR_102 = RG_rl_174 ;
	7'h57 :
		TR_102 = RG_rl_174 ;
	7'h58 :
		TR_102 = RG_rl_174 ;
	7'h59 :
		TR_102 = RG_rl_174 ;
	7'h5a :
		TR_102 = 9'h000 ;	// line#=../rle.cpp:79
	7'h5b :
		TR_102 = RG_rl_174 ;
	7'h5c :
		TR_102 = RG_rl_174 ;
	7'h5d :
		TR_102 = RG_rl_174 ;
	7'h5e :
		TR_102 = RG_rl_174 ;
	7'h5f :
		TR_102 = RG_rl_174 ;
	7'h60 :
		TR_102 = RG_rl_174 ;
	7'h61 :
		TR_102 = RG_rl_174 ;
	7'h62 :
		TR_102 = RG_rl_174 ;
	7'h63 :
		TR_102 = RG_rl_174 ;
	7'h64 :
		TR_102 = RG_rl_174 ;
	7'h65 :
		TR_102 = RG_rl_174 ;
	7'h66 :
		TR_102 = RG_rl_174 ;
	7'h67 :
		TR_102 = RG_rl_174 ;
	7'h68 :
		TR_102 = RG_rl_174 ;
	7'h69 :
		TR_102 = RG_rl_174 ;
	7'h6a :
		TR_102 = RG_rl_174 ;
	7'h6b :
		TR_102 = RG_rl_174 ;
	7'h6c :
		TR_102 = RG_rl_174 ;
	7'h6d :
		TR_102 = RG_rl_174 ;
	7'h6e :
		TR_102 = RG_rl_174 ;
	7'h6f :
		TR_102 = RG_rl_174 ;
	7'h70 :
		TR_102 = RG_rl_174 ;
	7'h71 :
		TR_102 = RG_rl_174 ;
	7'h72 :
		TR_102 = RG_rl_174 ;
	7'h73 :
		TR_102 = RG_rl_174 ;
	7'h74 :
		TR_102 = RG_rl_174 ;
	7'h75 :
		TR_102 = RG_rl_174 ;
	7'h76 :
		TR_102 = RG_rl_174 ;
	7'h77 :
		TR_102 = RG_rl_174 ;
	7'h78 :
		TR_102 = RG_rl_174 ;
	7'h79 :
		TR_102 = RG_rl_174 ;
	7'h7a :
		TR_102 = RG_rl_174 ;
	7'h7b :
		TR_102 = RG_rl_174 ;
	7'h7c :
		TR_102 = RG_rl_174 ;
	7'h7d :
		TR_102 = RG_rl_174 ;
	7'h7e :
		TR_102 = RG_rl_174 ;
	7'h7f :
		TR_102 = RG_rl_174 ;
	default :
		TR_102 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_43 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h01 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h02 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h03 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h04 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h05 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h06 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h07 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h08 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h09 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h0a :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h0b :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h0c :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h0d :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h0e :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h0f :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h10 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h11 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h12 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h13 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h14 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h15 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h16 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h17 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h18 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h19 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h1a :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h1b :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h1c :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h1d :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h1e :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h1f :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h20 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h21 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h22 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h23 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h24 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h25 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h26 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h27 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h28 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h29 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h2a :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h2b :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h2c :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h2d :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h2e :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h2f :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h30 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h31 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h32 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h33 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h34 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h35 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h36 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h37 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h38 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h39 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h3a :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h3b :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h3c :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h3d :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h3e :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h3f :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h40 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h41 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h42 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h43 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h44 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h45 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h46 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h47 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h48 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h49 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h4a :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h4b :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h4c :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h4d :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h4e :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h4f :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h50 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h51 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h52 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h53 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h54 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h55 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h56 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h57 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h58 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h59 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h5a :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h5b :
		TR_103 = 9'h000 ;	// line#=../rle.cpp:79
	7'h5c :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h5d :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h5e :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h5f :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h60 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h61 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h62 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h63 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h64 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h65 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h66 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h67 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h68 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h69 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h6a :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h6b :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h6c :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h6d :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h6e :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h6f :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h70 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h71 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h72 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h73 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h74 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h75 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h76 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h77 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h78 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h79 :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h7a :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h7b :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h7c :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h7d :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h7e :
		TR_103 = RG_quantized_block_rl_43 ;
	7'h7f :
		TR_103 = RG_quantized_block_rl_43 ;
	default :
		TR_103 = 9'hx ;
	endcase
always @ ( RG_rl_175 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_104 = RG_rl_175 ;
	7'h01 :
		TR_104 = RG_rl_175 ;
	7'h02 :
		TR_104 = RG_rl_175 ;
	7'h03 :
		TR_104 = RG_rl_175 ;
	7'h04 :
		TR_104 = RG_rl_175 ;
	7'h05 :
		TR_104 = RG_rl_175 ;
	7'h06 :
		TR_104 = RG_rl_175 ;
	7'h07 :
		TR_104 = RG_rl_175 ;
	7'h08 :
		TR_104 = RG_rl_175 ;
	7'h09 :
		TR_104 = RG_rl_175 ;
	7'h0a :
		TR_104 = RG_rl_175 ;
	7'h0b :
		TR_104 = RG_rl_175 ;
	7'h0c :
		TR_104 = RG_rl_175 ;
	7'h0d :
		TR_104 = RG_rl_175 ;
	7'h0e :
		TR_104 = RG_rl_175 ;
	7'h0f :
		TR_104 = RG_rl_175 ;
	7'h10 :
		TR_104 = RG_rl_175 ;
	7'h11 :
		TR_104 = RG_rl_175 ;
	7'h12 :
		TR_104 = RG_rl_175 ;
	7'h13 :
		TR_104 = RG_rl_175 ;
	7'h14 :
		TR_104 = RG_rl_175 ;
	7'h15 :
		TR_104 = RG_rl_175 ;
	7'h16 :
		TR_104 = RG_rl_175 ;
	7'h17 :
		TR_104 = RG_rl_175 ;
	7'h18 :
		TR_104 = RG_rl_175 ;
	7'h19 :
		TR_104 = RG_rl_175 ;
	7'h1a :
		TR_104 = RG_rl_175 ;
	7'h1b :
		TR_104 = RG_rl_175 ;
	7'h1c :
		TR_104 = RG_rl_175 ;
	7'h1d :
		TR_104 = RG_rl_175 ;
	7'h1e :
		TR_104 = RG_rl_175 ;
	7'h1f :
		TR_104 = RG_rl_175 ;
	7'h20 :
		TR_104 = RG_rl_175 ;
	7'h21 :
		TR_104 = RG_rl_175 ;
	7'h22 :
		TR_104 = RG_rl_175 ;
	7'h23 :
		TR_104 = RG_rl_175 ;
	7'h24 :
		TR_104 = RG_rl_175 ;
	7'h25 :
		TR_104 = RG_rl_175 ;
	7'h26 :
		TR_104 = RG_rl_175 ;
	7'h27 :
		TR_104 = RG_rl_175 ;
	7'h28 :
		TR_104 = RG_rl_175 ;
	7'h29 :
		TR_104 = RG_rl_175 ;
	7'h2a :
		TR_104 = RG_rl_175 ;
	7'h2b :
		TR_104 = RG_rl_175 ;
	7'h2c :
		TR_104 = RG_rl_175 ;
	7'h2d :
		TR_104 = RG_rl_175 ;
	7'h2e :
		TR_104 = RG_rl_175 ;
	7'h2f :
		TR_104 = RG_rl_175 ;
	7'h30 :
		TR_104 = RG_rl_175 ;
	7'h31 :
		TR_104 = RG_rl_175 ;
	7'h32 :
		TR_104 = RG_rl_175 ;
	7'h33 :
		TR_104 = RG_rl_175 ;
	7'h34 :
		TR_104 = RG_rl_175 ;
	7'h35 :
		TR_104 = RG_rl_175 ;
	7'h36 :
		TR_104 = RG_rl_175 ;
	7'h37 :
		TR_104 = RG_rl_175 ;
	7'h38 :
		TR_104 = RG_rl_175 ;
	7'h39 :
		TR_104 = RG_rl_175 ;
	7'h3a :
		TR_104 = RG_rl_175 ;
	7'h3b :
		TR_104 = RG_rl_175 ;
	7'h3c :
		TR_104 = RG_rl_175 ;
	7'h3d :
		TR_104 = RG_rl_175 ;
	7'h3e :
		TR_104 = RG_rl_175 ;
	7'h3f :
		TR_104 = RG_rl_175 ;
	7'h40 :
		TR_104 = RG_rl_175 ;
	7'h41 :
		TR_104 = RG_rl_175 ;
	7'h42 :
		TR_104 = RG_rl_175 ;
	7'h43 :
		TR_104 = RG_rl_175 ;
	7'h44 :
		TR_104 = RG_rl_175 ;
	7'h45 :
		TR_104 = RG_rl_175 ;
	7'h46 :
		TR_104 = RG_rl_175 ;
	7'h47 :
		TR_104 = RG_rl_175 ;
	7'h48 :
		TR_104 = RG_rl_175 ;
	7'h49 :
		TR_104 = RG_rl_175 ;
	7'h4a :
		TR_104 = RG_rl_175 ;
	7'h4b :
		TR_104 = RG_rl_175 ;
	7'h4c :
		TR_104 = RG_rl_175 ;
	7'h4d :
		TR_104 = RG_rl_175 ;
	7'h4e :
		TR_104 = RG_rl_175 ;
	7'h4f :
		TR_104 = RG_rl_175 ;
	7'h50 :
		TR_104 = RG_rl_175 ;
	7'h51 :
		TR_104 = RG_rl_175 ;
	7'h52 :
		TR_104 = RG_rl_175 ;
	7'h53 :
		TR_104 = RG_rl_175 ;
	7'h54 :
		TR_104 = RG_rl_175 ;
	7'h55 :
		TR_104 = RG_rl_175 ;
	7'h56 :
		TR_104 = RG_rl_175 ;
	7'h57 :
		TR_104 = RG_rl_175 ;
	7'h58 :
		TR_104 = RG_rl_175 ;
	7'h59 :
		TR_104 = RG_rl_175 ;
	7'h5a :
		TR_104 = RG_rl_175 ;
	7'h5b :
		TR_104 = RG_rl_175 ;
	7'h5c :
		TR_104 = 9'h000 ;	// line#=../rle.cpp:79
	7'h5d :
		TR_104 = RG_rl_175 ;
	7'h5e :
		TR_104 = RG_rl_175 ;
	7'h5f :
		TR_104 = RG_rl_175 ;
	7'h60 :
		TR_104 = RG_rl_175 ;
	7'h61 :
		TR_104 = RG_rl_175 ;
	7'h62 :
		TR_104 = RG_rl_175 ;
	7'h63 :
		TR_104 = RG_rl_175 ;
	7'h64 :
		TR_104 = RG_rl_175 ;
	7'h65 :
		TR_104 = RG_rl_175 ;
	7'h66 :
		TR_104 = RG_rl_175 ;
	7'h67 :
		TR_104 = RG_rl_175 ;
	7'h68 :
		TR_104 = RG_rl_175 ;
	7'h69 :
		TR_104 = RG_rl_175 ;
	7'h6a :
		TR_104 = RG_rl_175 ;
	7'h6b :
		TR_104 = RG_rl_175 ;
	7'h6c :
		TR_104 = RG_rl_175 ;
	7'h6d :
		TR_104 = RG_rl_175 ;
	7'h6e :
		TR_104 = RG_rl_175 ;
	7'h6f :
		TR_104 = RG_rl_175 ;
	7'h70 :
		TR_104 = RG_rl_175 ;
	7'h71 :
		TR_104 = RG_rl_175 ;
	7'h72 :
		TR_104 = RG_rl_175 ;
	7'h73 :
		TR_104 = RG_rl_175 ;
	7'h74 :
		TR_104 = RG_rl_175 ;
	7'h75 :
		TR_104 = RG_rl_175 ;
	7'h76 :
		TR_104 = RG_rl_175 ;
	7'h77 :
		TR_104 = RG_rl_175 ;
	7'h78 :
		TR_104 = RG_rl_175 ;
	7'h79 :
		TR_104 = RG_rl_175 ;
	7'h7a :
		TR_104 = RG_rl_175 ;
	7'h7b :
		TR_104 = RG_rl_175 ;
	7'h7c :
		TR_104 = RG_rl_175 ;
	7'h7d :
		TR_104 = RG_rl_175 ;
	7'h7e :
		TR_104 = RG_rl_175 ;
	7'h7f :
		TR_104 = RG_rl_175 ;
	default :
		TR_104 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_44 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h01 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h02 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h03 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h04 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h05 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h06 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h07 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h08 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h09 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h0a :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h0b :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h0c :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h0d :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h0e :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h0f :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h10 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h11 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h12 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h13 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h14 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h15 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h16 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h17 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h18 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h19 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h1a :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h1b :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h1c :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h1d :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h1e :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h1f :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h20 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h21 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h22 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h23 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h24 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h25 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h26 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h27 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h28 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h29 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h2a :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h2b :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h2c :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h2d :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h2e :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h2f :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h30 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h31 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h32 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h33 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h34 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h35 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h36 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h37 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h38 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h39 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h3a :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h3b :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h3c :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h3d :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h3e :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h3f :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h40 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h41 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h42 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h43 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h44 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h45 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h46 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h47 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h48 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h49 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h4a :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h4b :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h4c :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h4d :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h4e :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h4f :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h50 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h51 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h52 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h53 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h54 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h55 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h56 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h57 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h58 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h59 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h5a :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h5b :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h5c :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h5d :
		TR_105 = 9'h000 ;	// line#=../rle.cpp:79
	7'h5e :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h5f :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h60 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h61 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h62 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h63 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h64 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h65 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h66 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h67 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h68 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h69 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h6a :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h6b :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h6c :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h6d :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h6e :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h6f :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h70 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h71 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h72 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h73 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h74 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h75 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h76 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h77 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h78 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h79 :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h7a :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h7b :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h7c :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h7d :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h7e :
		TR_105 = RG_quantized_block_rl_44 ;
	7'h7f :
		TR_105 = RG_quantized_block_rl_44 ;
	default :
		TR_105 = 9'hx ;
	endcase
always @ ( RG_rl_176 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_106 = RG_rl_176 ;
	7'h01 :
		TR_106 = RG_rl_176 ;
	7'h02 :
		TR_106 = RG_rl_176 ;
	7'h03 :
		TR_106 = RG_rl_176 ;
	7'h04 :
		TR_106 = RG_rl_176 ;
	7'h05 :
		TR_106 = RG_rl_176 ;
	7'h06 :
		TR_106 = RG_rl_176 ;
	7'h07 :
		TR_106 = RG_rl_176 ;
	7'h08 :
		TR_106 = RG_rl_176 ;
	7'h09 :
		TR_106 = RG_rl_176 ;
	7'h0a :
		TR_106 = RG_rl_176 ;
	7'h0b :
		TR_106 = RG_rl_176 ;
	7'h0c :
		TR_106 = RG_rl_176 ;
	7'h0d :
		TR_106 = RG_rl_176 ;
	7'h0e :
		TR_106 = RG_rl_176 ;
	7'h0f :
		TR_106 = RG_rl_176 ;
	7'h10 :
		TR_106 = RG_rl_176 ;
	7'h11 :
		TR_106 = RG_rl_176 ;
	7'h12 :
		TR_106 = RG_rl_176 ;
	7'h13 :
		TR_106 = RG_rl_176 ;
	7'h14 :
		TR_106 = RG_rl_176 ;
	7'h15 :
		TR_106 = RG_rl_176 ;
	7'h16 :
		TR_106 = RG_rl_176 ;
	7'h17 :
		TR_106 = RG_rl_176 ;
	7'h18 :
		TR_106 = RG_rl_176 ;
	7'h19 :
		TR_106 = RG_rl_176 ;
	7'h1a :
		TR_106 = RG_rl_176 ;
	7'h1b :
		TR_106 = RG_rl_176 ;
	7'h1c :
		TR_106 = RG_rl_176 ;
	7'h1d :
		TR_106 = RG_rl_176 ;
	7'h1e :
		TR_106 = RG_rl_176 ;
	7'h1f :
		TR_106 = RG_rl_176 ;
	7'h20 :
		TR_106 = RG_rl_176 ;
	7'h21 :
		TR_106 = RG_rl_176 ;
	7'h22 :
		TR_106 = RG_rl_176 ;
	7'h23 :
		TR_106 = RG_rl_176 ;
	7'h24 :
		TR_106 = RG_rl_176 ;
	7'h25 :
		TR_106 = RG_rl_176 ;
	7'h26 :
		TR_106 = RG_rl_176 ;
	7'h27 :
		TR_106 = RG_rl_176 ;
	7'h28 :
		TR_106 = RG_rl_176 ;
	7'h29 :
		TR_106 = RG_rl_176 ;
	7'h2a :
		TR_106 = RG_rl_176 ;
	7'h2b :
		TR_106 = RG_rl_176 ;
	7'h2c :
		TR_106 = RG_rl_176 ;
	7'h2d :
		TR_106 = RG_rl_176 ;
	7'h2e :
		TR_106 = RG_rl_176 ;
	7'h2f :
		TR_106 = RG_rl_176 ;
	7'h30 :
		TR_106 = RG_rl_176 ;
	7'h31 :
		TR_106 = RG_rl_176 ;
	7'h32 :
		TR_106 = RG_rl_176 ;
	7'h33 :
		TR_106 = RG_rl_176 ;
	7'h34 :
		TR_106 = RG_rl_176 ;
	7'h35 :
		TR_106 = RG_rl_176 ;
	7'h36 :
		TR_106 = RG_rl_176 ;
	7'h37 :
		TR_106 = RG_rl_176 ;
	7'h38 :
		TR_106 = RG_rl_176 ;
	7'h39 :
		TR_106 = RG_rl_176 ;
	7'h3a :
		TR_106 = RG_rl_176 ;
	7'h3b :
		TR_106 = RG_rl_176 ;
	7'h3c :
		TR_106 = RG_rl_176 ;
	7'h3d :
		TR_106 = RG_rl_176 ;
	7'h3e :
		TR_106 = RG_rl_176 ;
	7'h3f :
		TR_106 = RG_rl_176 ;
	7'h40 :
		TR_106 = RG_rl_176 ;
	7'h41 :
		TR_106 = RG_rl_176 ;
	7'h42 :
		TR_106 = RG_rl_176 ;
	7'h43 :
		TR_106 = RG_rl_176 ;
	7'h44 :
		TR_106 = RG_rl_176 ;
	7'h45 :
		TR_106 = RG_rl_176 ;
	7'h46 :
		TR_106 = RG_rl_176 ;
	7'h47 :
		TR_106 = RG_rl_176 ;
	7'h48 :
		TR_106 = RG_rl_176 ;
	7'h49 :
		TR_106 = RG_rl_176 ;
	7'h4a :
		TR_106 = RG_rl_176 ;
	7'h4b :
		TR_106 = RG_rl_176 ;
	7'h4c :
		TR_106 = RG_rl_176 ;
	7'h4d :
		TR_106 = RG_rl_176 ;
	7'h4e :
		TR_106 = RG_rl_176 ;
	7'h4f :
		TR_106 = RG_rl_176 ;
	7'h50 :
		TR_106 = RG_rl_176 ;
	7'h51 :
		TR_106 = RG_rl_176 ;
	7'h52 :
		TR_106 = RG_rl_176 ;
	7'h53 :
		TR_106 = RG_rl_176 ;
	7'h54 :
		TR_106 = RG_rl_176 ;
	7'h55 :
		TR_106 = RG_rl_176 ;
	7'h56 :
		TR_106 = RG_rl_176 ;
	7'h57 :
		TR_106 = RG_rl_176 ;
	7'h58 :
		TR_106 = RG_rl_176 ;
	7'h59 :
		TR_106 = RG_rl_176 ;
	7'h5a :
		TR_106 = RG_rl_176 ;
	7'h5b :
		TR_106 = RG_rl_176 ;
	7'h5c :
		TR_106 = RG_rl_176 ;
	7'h5d :
		TR_106 = RG_rl_176 ;
	7'h5e :
		TR_106 = 9'h000 ;	// line#=../rle.cpp:79
	7'h5f :
		TR_106 = RG_rl_176 ;
	7'h60 :
		TR_106 = RG_rl_176 ;
	7'h61 :
		TR_106 = RG_rl_176 ;
	7'h62 :
		TR_106 = RG_rl_176 ;
	7'h63 :
		TR_106 = RG_rl_176 ;
	7'h64 :
		TR_106 = RG_rl_176 ;
	7'h65 :
		TR_106 = RG_rl_176 ;
	7'h66 :
		TR_106 = RG_rl_176 ;
	7'h67 :
		TR_106 = RG_rl_176 ;
	7'h68 :
		TR_106 = RG_rl_176 ;
	7'h69 :
		TR_106 = RG_rl_176 ;
	7'h6a :
		TR_106 = RG_rl_176 ;
	7'h6b :
		TR_106 = RG_rl_176 ;
	7'h6c :
		TR_106 = RG_rl_176 ;
	7'h6d :
		TR_106 = RG_rl_176 ;
	7'h6e :
		TR_106 = RG_rl_176 ;
	7'h6f :
		TR_106 = RG_rl_176 ;
	7'h70 :
		TR_106 = RG_rl_176 ;
	7'h71 :
		TR_106 = RG_rl_176 ;
	7'h72 :
		TR_106 = RG_rl_176 ;
	7'h73 :
		TR_106 = RG_rl_176 ;
	7'h74 :
		TR_106 = RG_rl_176 ;
	7'h75 :
		TR_106 = RG_rl_176 ;
	7'h76 :
		TR_106 = RG_rl_176 ;
	7'h77 :
		TR_106 = RG_rl_176 ;
	7'h78 :
		TR_106 = RG_rl_176 ;
	7'h79 :
		TR_106 = RG_rl_176 ;
	7'h7a :
		TR_106 = RG_rl_176 ;
	7'h7b :
		TR_106 = RG_rl_176 ;
	7'h7c :
		TR_106 = RG_rl_176 ;
	7'h7d :
		TR_106 = RG_rl_176 ;
	7'h7e :
		TR_106 = RG_rl_176 ;
	7'h7f :
		TR_106 = RG_rl_176 ;
	default :
		TR_106 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_45 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h01 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h02 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h03 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h04 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h05 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h06 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h07 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h08 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h09 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h0a :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h0b :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h0c :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h0d :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h0e :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h0f :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h10 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h11 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h12 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h13 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h14 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h15 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h16 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h17 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h18 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h19 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h1a :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h1b :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h1c :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h1d :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h1e :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h1f :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h20 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h21 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h22 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h23 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h24 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h25 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h26 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h27 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h28 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h29 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h2a :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h2b :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h2c :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h2d :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h2e :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h2f :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h30 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h31 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h32 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h33 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h34 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h35 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h36 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h37 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h38 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h39 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h3a :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h3b :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h3c :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h3d :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h3e :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h3f :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h40 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h41 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h42 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h43 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h44 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h45 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h46 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h47 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h48 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h49 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h4a :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h4b :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h4c :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h4d :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h4e :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h4f :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h50 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h51 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h52 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h53 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h54 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h55 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h56 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h57 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h58 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h59 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h5a :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h5b :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h5c :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h5d :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h5e :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h5f :
		TR_107 = 9'h000 ;	// line#=../rle.cpp:79
	7'h60 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h61 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h62 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h63 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h64 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h65 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h66 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h67 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h68 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h69 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h6a :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h6b :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h6c :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h6d :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h6e :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h6f :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h70 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h71 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h72 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h73 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h74 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h75 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h76 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h77 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h78 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h79 :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h7a :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h7b :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h7c :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h7d :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h7e :
		TR_107 = RG_quantized_block_rl_45 ;
	7'h7f :
		TR_107 = RG_quantized_block_rl_45 ;
	default :
		TR_107 = 9'hx ;
	endcase
always @ ( RG_rl_177 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_108 = RG_rl_177 ;
	7'h01 :
		TR_108 = RG_rl_177 ;
	7'h02 :
		TR_108 = RG_rl_177 ;
	7'h03 :
		TR_108 = RG_rl_177 ;
	7'h04 :
		TR_108 = RG_rl_177 ;
	7'h05 :
		TR_108 = RG_rl_177 ;
	7'h06 :
		TR_108 = RG_rl_177 ;
	7'h07 :
		TR_108 = RG_rl_177 ;
	7'h08 :
		TR_108 = RG_rl_177 ;
	7'h09 :
		TR_108 = RG_rl_177 ;
	7'h0a :
		TR_108 = RG_rl_177 ;
	7'h0b :
		TR_108 = RG_rl_177 ;
	7'h0c :
		TR_108 = RG_rl_177 ;
	7'h0d :
		TR_108 = RG_rl_177 ;
	7'h0e :
		TR_108 = RG_rl_177 ;
	7'h0f :
		TR_108 = RG_rl_177 ;
	7'h10 :
		TR_108 = RG_rl_177 ;
	7'h11 :
		TR_108 = RG_rl_177 ;
	7'h12 :
		TR_108 = RG_rl_177 ;
	7'h13 :
		TR_108 = RG_rl_177 ;
	7'h14 :
		TR_108 = RG_rl_177 ;
	7'h15 :
		TR_108 = RG_rl_177 ;
	7'h16 :
		TR_108 = RG_rl_177 ;
	7'h17 :
		TR_108 = RG_rl_177 ;
	7'h18 :
		TR_108 = RG_rl_177 ;
	7'h19 :
		TR_108 = RG_rl_177 ;
	7'h1a :
		TR_108 = RG_rl_177 ;
	7'h1b :
		TR_108 = RG_rl_177 ;
	7'h1c :
		TR_108 = RG_rl_177 ;
	7'h1d :
		TR_108 = RG_rl_177 ;
	7'h1e :
		TR_108 = RG_rl_177 ;
	7'h1f :
		TR_108 = RG_rl_177 ;
	7'h20 :
		TR_108 = RG_rl_177 ;
	7'h21 :
		TR_108 = RG_rl_177 ;
	7'h22 :
		TR_108 = RG_rl_177 ;
	7'h23 :
		TR_108 = RG_rl_177 ;
	7'h24 :
		TR_108 = RG_rl_177 ;
	7'h25 :
		TR_108 = RG_rl_177 ;
	7'h26 :
		TR_108 = RG_rl_177 ;
	7'h27 :
		TR_108 = RG_rl_177 ;
	7'h28 :
		TR_108 = RG_rl_177 ;
	7'h29 :
		TR_108 = RG_rl_177 ;
	7'h2a :
		TR_108 = RG_rl_177 ;
	7'h2b :
		TR_108 = RG_rl_177 ;
	7'h2c :
		TR_108 = RG_rl_177 ;
	7'h2d :
		TR_108 = RG_rl_177 ;
	7'h2e :
		TR_108 = RG_rl_177 ;
	7'h2f :
		TR_108 = RG_rl_177 ;
	7'h30 :
		TR_108 = RG_rl_177 ;
	7'h31 :
		TR_108 = RG_rl_177 ;
	7'h32 :
		TR_108 = RG_rl_177 ;
	7'h33 :
		TR_108 = RG_rl_177 ;
	7'h34 :
		TR_108 = RG_rl_177 ;
	7'h35 :
		TR_108 = RG_rl_177 ;
	7'h36 :
		TR_108 = RG_rl_177 ;
	7'h37 :
		TR_108 = RG_rl_177 ;
	7'h38 :
		TR_108 = RG_rl_177 ;
	7'h39 :
		TR_108 = RG_rl_177 ;
	7'h3a :
		TR_108 = RG_rl_177 ;
	7'h3b :
		TR_108 = RG_rl_177 ;
	7'h3c :
		TR_108 = RG_rl_177 ;
	7'h3d :
		TR_108 = RG_rl_177 ;
	7'h3e :
		TR_108 = RG_rl_177 ;
	7'h3f :
		TR_108 = RG_rl_177 ;
	7'h40 :
		TR_108 = RG_rl_177 ;
	7'h41 :
		TR_108 = RG_rl_177 ;
	7'h42 :
		TR_108 = RG_rl_177 ;
	7'h43 :
		TR_108 = RG_rl_177 ;
	7'h44 :
		TR_108 = RG_rl_177 ;
	7'h45 :
		TR_108 = RG_rl_177 ;
	7'h46 :
		TR_108 = RG_rl_177 ;
	7'h47 :
		TR_108 = RG_rl_177 ;
	7'h48 :
		TR_108 = RG_rl_177 ;
	7'h49 :
		TR_108 = RG_rl_177 ;
	7'h4a :
		TR_108 = RG_rl_177 ;
	7'h4b :
		TR_108 = RG_rl_177 ;
	7'h4c :
		TR_108 = RG_rl_177 ;
	7'h4d :
		TR_108 = RG_rl_177 ;
	7'h4e :
		TR_108 = RG_rl_177 ;
	7'h4f :
		TR_108 = RG_rl_177 ;
	7'h50 :
		TR_108 = RG_rl_177 ;
	7'h51 :
		TR_108 = RG_rl_177 ;
	7'h52 :
		TR_108 = RG_rl_177 ;
	7'h53 :
		TR_108 = RG_rl_177 ;
	7'h54 :
		TR_108 = RG_rl_177 ;
	7'h55 :
		TR_108 = RG_rl_177 ;
	7'h56 :
		TR_108 = RG_rl_177 ;
	7'h57 :
		TR_108 = RG_rl_177 ;
	7'h58 :
		TR_108 = RG_rl_177 ;
	7'h59 :
		TR_108 = RG_rl_177 ;
	7'h5a :
		TR_108 = RG_rl_177 ;
	7'h5b :
		TR_108 = RG_rl_177 ;
	7'h5c :
		TR_108 = RG_rl_177 ;
	7'h5d :
		TR_108 = RG_rl_177 ;
	7'h5e :
		TR_108 = RG_rl_177 ;
	7'h5f :
		TR_108 = RG_rl_177 ;
	7'h60 :
		TR_108 = 9'h000 ;	// line#=../rle.cpp:79
	7'h61 :
		TR_108 = RG_rl_177 ;
	7'h62 :
		TR_108 = RG_rl_177 ;
	7'h63 :
		TR_108 = RG_rl_177 ;
	7'h64 :
		TR_108 = RG_rl_177 ;
	7'h65 :
		TR_108 = RG_rl_177 ;
	7'h66 :
		TR_108 = RG_rl_177 ;
	7'h67 :
		TR_108 = RG_rl_177 ;
	7'h68 :
		TR_108 = RG_rl_177 ;
	7'h69 :
		TR_108 = RG_rl_177 ;
	7'h6a :
		TR_108 = RG_rl_177 ;
	7'h6b :
		TR_108 = RG_rl_177 ;
	7'h6c :
		TR_108 = RG_rl_177 ;
	7'h6d :
		TR_108 = RG_rl_177 ;
	7'h6e :
		TR_108 = RG_rl_177 ;
	7'h6f :
		TR_108 = RG_rl_177 ;
	7'h70 :
		TR_108 = RG_rl_177 ;
	7'h71 :
		TR_108 = RG_rl_177 ;
	7'h72 :
		TR_108 = RG_rl_177 ;
	7'h73 :
		TR_108 = RG_rl_177 ;
	7'h74 :
		TR_108 = RG_rl_177 ;
	7'h75 :
		TR_108 = RG_rl_177 ;
	7'h76 :
		TR_108 = RG_rl_177 ;
	7'h77 :
		TR_108 = RG_rl_177 ;
	7'h78 :
		TR_108 = RG_rl_177 ;
	7'h79 :
		TR_108 = RG_rl_177 ;
	7'h7a :
		TR_108 = RG_rl_177 ;
	7'h7b :
		TR_108 = RG_rl_177 ;
	7'h7c :
		TR_108 = RG_rl_177 ;
	7'h7d :
		TR_108 = RG_rl_177 ;
	7'h7e :
		TR_108 = RG_rl_177 ;
	7'h7f :
		TR_108 = RG_rl_177 ;
	default :
		TR_108 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_46 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h01 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h02 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h03 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h04 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h05 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h06 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h07 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h08 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h09 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h0a :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h0b :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h0c :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h0d :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h0e :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h0f :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h10 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h11 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h12 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h13 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h14 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h15 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h16 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h17 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h18 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h19 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h1a :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h1b :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h1c :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h1d :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h1e :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h1f :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h20 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h21 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h22 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h23 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h24 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h25 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h26 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h27 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h28 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h29 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h2a :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h2b :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h2c :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h2d :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h2e :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h2f :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h30 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h31 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h32 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h33 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h34 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h35 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h36 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h37 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h38 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h39 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h3a :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h3b :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h3c :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h3d :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h3e :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h3f :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h40 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h41 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h42 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h43 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h44 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h45 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h46 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h47 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h48 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h49 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h4a :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h4b :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h4c :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h4d :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h4e :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h4f :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h50 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h51 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h52 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h53 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h54 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h55 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h56 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h57 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h58 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h59 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h5a :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h5b :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h5c :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h5d :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h5e :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h5f :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h60 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h61 :
		TR_109 = 9'h000 ;	// line#=../rle.cpp:79
	7'h62 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h63 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h64 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h65 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h66 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h67 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h68 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h69 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h6a :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h6b :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h6c :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h6d :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h6e :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h6f :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h70 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h71 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h72 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h73 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h74 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h75 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h76 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h77 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h78 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h79 :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h7a :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h7b :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h7c :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h7d :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h7e :
		TR_109 = RG_quantized_block_rl_46 ;
	7'h7f :
		TR_109 = RG_quantized_block_rl_46 ;
	default :
		TR_109 = 9'hx ;
	endcase
always @ ( RG_rl_178 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_110 = RG_rl_178 ;
	7'h01 :
		TR_110 = RG_rl_178 ;
	7'h02 :
		TR_110 = RG_rl_178 ;
	7'h03 :
		TR_110 = RG_rl_178 ;
	7'h04 :
		TR_110 = RG_rl_178 ;
	7'h05 :
		TR_110 = RG_rl_178 ;
	7'h06 :
		TR_110 = RG_rl_178 ;
	7'h07 :
		TR_110 = RG_rl_178 ;
	7'h08 :
		TR_110 = RG_rl_178 ;
	7'h09 :
		TR_110 = RG_rl_178 ;
	7'h0a :
		TR_110 = RG_rl_178 ;
	7'h0b :
		TR_110 = RG_rl_178 ;
	7'h0c :
		TR_110 = RG_rl_178 ;
	7'h0d :
		TR_110 = RG_rl_178 ;
	7'h0e :
		TR_110 = RG_rl_178 ;
	7'h0f :
		TR_110 = RG_rl_178 ;
	7'h10 :
		TR_110 = RG_rl_178 ;
	7'h11 :
		TR_110 = RG_rl_178 ;
	7'h12 :
		TR_110 = RG_rl_178 ;
	7'h13 :
		TR_110 = RG_rl_178 ;
	7'h14 :
		TR_110 = RG_rl_178 ;
	7'h15 :
		TR_110 = RG_rl_178 ;
	7'h16 :
		TR_110 = RG_rl_178 ;
	7'h17 :
		TR_110 = RG_rl_178 ;
	7'h18 :
		TR_110 = RG_rl_178 ;
	7'h19 :
		TR_110 = RG_rl_178 ;
	7'h1a :
		TR_110 = RG_rl_178 ;
	7'h1b :
		TR_110 = RG_rl_178 ;
	7'h1c :
		TR_110 = RG_rl_178 ;
	7'h1d :
		TR_110 = RG_rl_178 ;
	7'h1e :
		TR_110 = RG_rl_178 ;
	7'h1f :
		TR_110 = RG_rl_178 ;
	7'h20 :
		TR_110 = RG_rl_178 ;
	7'h21 :
		TR_110 = RG_rl_178 ;
	7'h22 :
		TR_110 = RG_rl_178 ;
	7'h23 :
		TR_110 = RG_rl_178 ;
	7'h24 :
		TR_110 = RG_rl_178 ;
	7'h25 :
		TR_110 = RG_rl_178 ;
	7'h26 :
		TR_110 = RG_rl_178 ;
	7'h27 :
		TR_110 = RG_rl_178 ;
	7'h28 :
		TR_110 = RG_rl_178 ;
	7'h29 :
		TR_110 = RG_rl_178 ;
	7'h2a :
		TR_110 = RG_rl_178 ;
	7'h2b :
		TR_110 = RG_rl_178 ;
	7'h2c :
		TR_110 = RG_rl_178 ;
	7'h2d :
		TR_110 = RG_rl_178 ;
	7'h2e :
		TR_110 = RG_rl_178 ;
	7'h2f :
		TR_110 = RG_rl_178 ;
	7'h30 :
		TR_110 = RG_rl_178 ;
	7'h31 :
		TR_110 = RG_rl_178 ;
	7'h32 :
		TR_110 = RG_rl_178 ;
	7'h33 :
		TR_110 = RG_rl_178 ;
	7'h34 :
		TR_110 = RG_rl_178 ;
	7'h35 :
		TR_110 = RG_rl_178 ;
	7'h36 :
		TR_110 = RG_rl_178 ;
	7'h37 :
		TR_110 = RG_rl_178 ;
	7'h38 :
		TR_110 = RG_rl_178 ;
	7'h39 :
		TR_110 = RG_rl_178 ;
	7'h3a :
		TR_110 = RG_rl_178 ;
	7'h3b :
		TR_110 = RG_rl_178 ;
	7'h3c :
		TR_110 = RG_rl_178 ;
	7'h3d :
		TR_110 = RG_rl_178 ;
	7'h3e :
		TR_110 = RG_rl_178 ;
	7'h3f :
		TR_110 = RG_rl_178 ;
	7'h40 :
		TR_110 = RG_rl_178 ;
	7'h41 :
		TR_110 = RG_rl_178 ;
	7'h42 :
		TR_110 = RG_rl_178 ;
	7'h43 :
		TR_110 = RG_rl_178 ;
	7'h44 :
		TR_110 = RG_rl_178 ;
	7'h45 :
		TR_110 = RG_rl_178 ;
	7'h46 :
		TR_110 = RG_rl_178 ;
	7'h47 :
		TR_110 = RG_rl_178 ;
	7'h48 :
		TR_110 = RG_rl_178 ;
	7'h49 :
		TR_110 = RG_rl_178 ;
	7'h4a :
		TR_110 = RG_rl_178 ;
	7'h4b :
		TR_110 = RG_rl_178 ;
	7'h4c :
		TR_110 = RG_rl_178 ;
	7'h4d :
		TR_110 = RG_rl_178 ;
	7'h4e :
		TR_110 = RG_rl_178 ;
	7'h4f :
		TR_110 = RG_rl_178 ;
	7'h50 :
		TR_110 = RG_rl_178 ;
	7'h51 :
		TR_110 = RG_rl_178 ;
	7'h52 :
		TR_110 = RG_rl_178 ;
	7'h53 :
		TR_110 = RG_rl_178 ;
	7'h54 :
		TR_110 = RG_rl_178 ;
	7'h55 :
		TR_110 = RG_rl_178 ;
	7'h56 :
		TR_110 = RG_rl_178 ;
	7'h57 :
		TR_110 = RG_rl_178 ;
	7'h58 :
		TR_110 = RG_rl_178 ;
	7'h59 :
		TR_110 = RG_rl_178 ;
	7'h5a :
		TR_110 = RG_rl_178 ;
	7'h5b :
		TR_110 = RG_rl_178 ;
	7'h5c :
		TR_110 = RG_rl_178 ;
	7'h5d :
		TR_110 = RG_rl_178 ;
	7'h5e :
		TR_110 = RG_rl_178 ;
	7'h5f :
		TR_110 = RG_rl_178 ;
	7'h60 :
		TR_110 = RG_rl_178 ;
	7'h61 :
		TR_110 = RG_rl_178 ;
	7'h62 :
		TR_110 = 9'h000 ;	// line#=../rle.cpp:79
	7'h63 :
		TR_110 = RG_rl_178 ;
	7'h64 :
		TR_110 = RG_rl_178 ;
	7'h65 :
		TR_110 = RG_rl_178 ;
	7'h66 :
		TR_110 = RG_rl_178 ;
	7'h67 :
		TR_110 = RG_rl_178 ;
	7'h68 :
		TR_110 = RG_rl_178 ;
	7'h69 :
		TR_110 = RG_rl_178 ;
	7'h6a :
		TR_110 = RG_rl_178 ;
	7'h6b :
		TR_110 = RG_rl_178 ;
	7'h6c :
		TR_110 = RG_rl_178 ;
	7'h6d :
		TR_110 = RG_rl_178 ;
	7'h6e :
		TR_110 = RG_rl_178 ;
	7'h6f :
		TR_110 = RG_rl_178 ;
	7'h70 :
		TR_110 = RG_rl_178 ;
	7'h71 :
		TR_110 = RG_rl_178 ;
	7'h72 :
		TR_110 = RG_rl_178 ;
	7'h73 :
		TR_110 = RG_rl_178 ;
	7'h74 :
		TR_110 = RG_rl_178 ;
	7'h75 :
		TR_110 = RG_rl_178 ;
	7'h76 :
		TR_110 = RG_rl_178 ;
	7'h77 :
		TR_110 = RG_rl_178 ;
	7'h78 :
		TR_110 = RG_rl_178 ;
	7'h79 :
		TR_110 = RG_rl_178 ;
	7'h7a :
		TR_110 = RG_rl_178 ;
	7'h7b :
		TR_110 = RG_rl_178 ;
	7'h7c :
		TR_110 = RG_rl_178 ;
	7'h7d :
		TR_110 = RG_rl_178 ;
	7'h7e :
		TR_110 = RG_rl_178 ;
	7'h7f :
		TR_110 = RG_rl_178 ;
	default :
		TR_110 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_47 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h01 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h02 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h03 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h04 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h05 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h06 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h07 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h08 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h09 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h0a :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h0b :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h0c :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h0d :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h0e :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h0f :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h10 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h11 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h12 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h13 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h14 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h15 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h16 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h17 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h18 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h19 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h1a :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h1b :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h1c :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h1d :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h1e :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h1f :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h20 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h21 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h22 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h23 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h24 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h25 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h26 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h27 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h28 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h29 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h2a :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h2b :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h2c :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h2d :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h2e :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h2f :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h30 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h31 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h32 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h33 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h34 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h35 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h36 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h37 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h38 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h39 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h3a :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h3b :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h3c :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h3d :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h3e :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h3f :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h40 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h41 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h42 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h43 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h44 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h45 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h46 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h47 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h48 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h49 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h4a :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h4b :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h4c :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h4d :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h4e :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h4f :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h50 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h51 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h52 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h53 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h54 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h55 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h56 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h57 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h58 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h59 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h5a :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h5b :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h5c :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h5d :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h5e :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h5f :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h60 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h61 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h62 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h63 :
		TR_111 = 9'h000 ;	// line#=../rle.cpp:79
	7'h64 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h65 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h66 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h67 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h68 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h69 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h6a :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h6b :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h6c :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h6d :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h6e :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h6f :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h70 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h71 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h72 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h73 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h74 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h75 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h76 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h77 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h78 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h79 :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h7a :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h7b :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h7c :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h7d :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h7e :
		TR_111 = RG_quantized_block_rl_47 ;
	7'h7f :
		TR_111 = RG_quantized_block_rl_47 ;
	default :
		TR_111 = 9'hx ;
	endcase
always @ ( RG_rl_179 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_112 = RG_rl_179 ;
	7'h01 :
		TR_112 = RG_rl_179 ;
	7'h02 :
		TR_112 = RG_rl_179 ;
	7'h03 :
		TR_112 = RG_rl_179 ;
	7'h04 :
		TR_112 = RG_rl_179 ;
	7'h05 :
		TR_112 = RG_rl_179 ;
	7'h06 :
		TR_112 = RG_rl_179 ;
	7'h07 :
		TR_112 = RG_rl_179 ;
	7'h08 :
		TR_112 = RG_rl_179 ;
	7'h09 :
		TR_112 = RG_rl_179 ;
	7'h0a :
		TR_112 = RG_rl_179 ;
	7'h0b :
		TR_112 = RG_rl_179 ;
	7'h0c :
		TR_112 = RG_rl_179 ;
	7'h0d :
		TR_112 = RG_rl_179 ;
	7'h0e :
		TR_112 = RG_rl_179 ;
	7'h0f :
		TR_112 = RG_rl_179 ;
	7'h10 :
		TR_112 = RG_rl_179 ;
	7'h11 :
		TR_112 = RG_rl_179 ;
	7'h12 :
		TR_112 = RG_rl_179 ;
	7'h13 :
		TR_112 = RG_rl_179 ;
	7'h14 :
		TR_112 = RG_rl_179 ;
	7'h15 :
		TR_112 = RG_rl_179 ;
	7'h16 :
		TR_112 = RG_rl_179 ;
	7'h17 :
		TR_112 = RG_rl_179 ;
	7'h18 :
		TR_112 = RG_rl_179 ;
	7'h19 :
		TR_112 = RG_rl_179 ;
	7'h1a :
		TR_112 = RG_rl_179 ;
	7'h1b :
		TR_112 = RG_rl_179 ;
	7'h1c :
		TR_112 = RG_rl_179 ;
	7'h1d :
		TR_112 = RG_rl_179 ;
	7'h1e :
		TR_112 = RG_rl_179 ;
	7'h1f :
		TR_112 = RG_rl_179 ;
	7'h20 :
		TR_112 = RG_rl_179 ;
	7'h21 :
		TR_112 = RG_rl_179 ;
	7'h22 :
		TR_112 = RG_rl_179 ;
	7'h23 :
		TR_112 = RG_rl_179 ;
	7'h24 :
		TR_112 = RG_rl_179 ;
	7'h25 :
		TR_112 = RG_rl_179 ;
	7'h26 :
		TR_112 = RG_rl_179 ;
	7'h27 :
		TR_112 = RG_rl_179 ;
	7'h28 :
		TR_112 = RG_rl_179 ;
	7'h29 :
		TR_112 = RG_rl_179 ;
	7'h2a :
		TR_112 = RG_rl_179 ;
	7'h2b :
		TR_112 = RG_rl_179 ;
	7'h2c :
		TR_112 = RG_rl_179 ;
	7'h2d :
		TR_112 = RG_rl_179 ;
	7'h2e :
		TR_112 = RG_rl_179 ;
	7'h2f :
		TR_112 = RG_rl_179 ;
	7'h30 :
		TR_112 = RG_rl_179 ;
	7'h31 :
		TR_112 = RG_rl_179 ;
	7'h32 :
		TR_112 = RG_rl_179 ;
	7'h33 :
		TR_112 = RG_rl_179 ;
	7'h34 :
		TR_112 = RG_rl_179 ;
	7'h35 :
		TR_112 = RG_rl_179 ;
	7'h36 :
		TR_112 = RG_rl_179 ;
	7'h37 :
		TR_112 = RG_rl_179 ;
	7'h38 :
		TR_112 = RG_rl_179 ;
	7'h39 :
		TR_112 = RG_rl_179 ;
	7'h3a :
		TR_112 = RG_rl_179 ;
	7'h3b :
		TR_112 = RG_rl_179 ;
	7'h3c :
		TR_112 = RG_rl_179 ;
	7'h3d :
		TR_112 = RG_rl_179 ;
	7'h3e :
		TR_112 = RG_rl_179 ;
	7'h3f :
		TR_112 = RG_rl_179 ;
	7'h40 :
		TR_112 = RG_rl_179 ;
	7'h41 :
		TR_112 = RG_rl_179 ;
	7'h42 :
		TR_112 = RG_rl_179 ;
	7'h43 :
		TR_112 = RG_rl_179 ;
	7'h44 :
		TR_112 = RG_rl_179 ;
	7'h45 :
		TR_112 = RG_rl_179 ;
	7'h46 :
		TR_112 = RG_rl_179 ;
	7'h47 :
		TR_112 = RG_rl_179 ;
	7'h48 :
		TR_112 = RG_rl_179 ;
	7'h49 :
		TR_112 = RG_rl_179 ;
	7'h4a :
		TR_112 = RG_rl_179 ;
	7'h4b :
		TR_112 = RG_rl_179 ;
	7'h4c :
		TR_112 = RG_rl_179 ;
	7'h4d :
		TR_112 = RG_rl_179 ;
	7'h4e :
		TR_112 = RG_rl_179 ;
	7'h4f :
		TR_112 = RG_rl_179 ;
	7'h50 :
		TR_112 = RG_rl_179 ;
	7'h51 :
		TR_112 = RG_rl_179 ;
	7'h52 :
		TR_112 = RG_rl_179 ;
	7'h53 :
		TR_112 = RG_rl_179 ;
	7'h54 :
		TR_112 = RG_rl_179 ;
	7'h55 :
		TR_112 = RG_rl_179 ;
	7'h56 :
		TR_112 = RG_rl_179 ;
	7'h57 :
		TR_112 = RG_rl_179 ;
	7'h58 :
		TR_112 = RG_rl_179 ;
	7'h59 :
		TR_112 = RG_rl_179 ;
	7'h5a :
		TR_112 = RG_rl_179 ;
	7'h5b :
		TR_112 = RG_rl_179 ;
	7'h5c :
		TR_112 = RG_rl_179 ;
	7'h5d :
		TR_112 = RG_rl_179 ;
	7'h5e :
		TR_112 = RG_rl_179 ;
	7'h5f :
		TR_112 = RG_rl_179 ;
	7'h60 :
		TR_112 = RG_rl_179 ;
	7'h61 :
		TR_112 = RG_rl_179 ;
	7'h62 :
		TR_112 = RG_rl_179 ;
	7'h63 :
		TR_112 = RG_rl_179 ;
	7'h64 :
		TR_112 = 9'h000 ;	// line#=../rle.cpp:79
	7'h65 :
		TR_112 = RG_rl_179 ;
	7'h66 :
		TR_112 = RG_rl_179 ;
	7'h67 :
		TR_112 = RG_rl_179 ;
	7'h68 :
		TR_112 = RG_rl_179 ;
	7'h69 :
		TR_112 = RG_rl_179 ;
	7'h6a :
		TR_112 = RG_rl_179 ;
	7'h6b :
		TR_112 = RG_rl_179 ;
	7'h6c :
		TR_112 = RG_rl_179 ;
	7'h6d :
		TR_112 = RG_rl_179 ;
	7'h6e :
		TR_112 = RG_rl_179 ;
	7'h6f :
		TR_112 = RG_rl_179 ;
	7'h70 :
		TR_112 = RG_rl_179 ;
	7'h71 :
		TR_112 = RG_rl_179 ;
	7'h72 :
		TR_112 = RG_rl_179 ;
	7'h73 :
		TR_112 = RG_rl_179 ;
	7'h74 :
		TR_112 = RG_rl_179 ;
	7'h75 :
		TR_112 = RG_rl_179 ;
	7'h76 :
		TR_112 = RG_rl_179 ;
	7'h77 :
		TR_112 = RG_rl_179 ;
	7'h78 :
		TR_112 = RG_rl_179 ;
	7'h79 :
		TR_112 = RG_rl_179 ;
	7'h7a :
		TR_112 = RG_rl_179 ;
	7'h7b :
		TR_112 = RG_rl_179 ;
	7'h7c :
		TR_112 = RG_rl_179 ;
	7'h7d :
		TR_112 = RG_rl_179 ;
	7'h7e :
		TR_112 = RG_rl_179 ;
	7'h7f :
		TR_112 = RG_rl_179 ;
	default :
		TR_112 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_48 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h01 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h02 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h03 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h04 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h05 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h06 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h07 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h08 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h09 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h0a :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h0b :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h0c :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h0d :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h0e :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h0f :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h10 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h11 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h12 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h13 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h14 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h15 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h16 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h17 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h18 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h19 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h1a :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h1b :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h1c :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h1d :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h1e :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h1f :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h20 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h21 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h22 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h23 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h24 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h25 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h26 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h27 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h28 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h29 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h2a :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h2b :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h2c :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h2d :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h2e :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h2f :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h30 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h31 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h32 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h33 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h34 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h35 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h36 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h37 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h38 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h39 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h3a :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h3b :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h3c :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h3d :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h3e :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h3f :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h40 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h41 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h42 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h43 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h44 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h45 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h46 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h47 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h48 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h49 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h4a :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h4b :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h4c :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h4d :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h4e :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h4f :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h50 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h51 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h52 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h53 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h54 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h55 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h56 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h57 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h58 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h59 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h5a :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h5b :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h5c :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h5d :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h5e :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h5f :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h60 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h61 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h62 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h63 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h64 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h65 :
		TR_113 = 9'h000 ;	// line#=../rle.cpp:79
	7'h66 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h67 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h68 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h69 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h6a :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h6b :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h6c :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h6d :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h6e :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h6f :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h70 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h71 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h72 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h73 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h74 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h75 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h76 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h77 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h78 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h79 :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h7a :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h7b :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h7c :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h7d :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h7e :
		TR_113 = RG_quantized_block_rl_48 ;
	7'h7f :
		TR_113 = RG_quantized_block_rl_48 ;
	default :
		TR_113 = 9'hx ;
	endcase
always @ ( RG_rl_180 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_114 = RG_rl_180 ;
	7'h01 :
		TR_114 = RG_rl_180 ;
	7'h02 :
		TR_114 = RG_rl_180 ;
	7'h03 :
		TR_114 = RG_rl_180 ;
	7'h04 :
		TR_114 = RG_rl_180 ;
	7'h05 :
		TR_114 = RG_rl_180 ;
	7'h06 :
		TR_114 = RG_rl_180 ;
	7'h07 :
		TR_114 = RG_rl_180 ;
	7'h08 :
		TR_114 = RG_rl_180 ;
	7'h09 :
		TR_114 = RG_rl_180 ;
	7'h0a :
		TR_114 = RG_rl_180 ;
	7'h0b :
		TR_114 = RG_rl_180 ;
	7'h0c :
		TR_114 = RG_rl_180 ;
	7'h0d :
		TR_114 = RG_rl_180 ;
	7'h0e :
		TR_114 = RG_rl_180 ;
	7'h0f :
		TR_114 = RG_rl_180 ;
	7'h10 :
		TR_114 = RG_rl_180 ;
	7'h11 :
		TR_114 = RG_rl_180 ;
	7'h12 :
		TR_114 = RG_rl_180 ;
	7'h13 :
		TR_114 = RG_rl_180 ;
	7'h14 :
		TR_114 = RG_rl_180 ;
	7'h15 :
		TR_114 = RG_rl_180 ;
	7'h16 :
		TR_114 = RG_rl_180 ;
	7'h17 :
		TR_114 = RG_rl_180 ;
	7'h18 :
		TR_114 = RG_rl_180 ;
	7'h19 :
		TR_114 = RG_rl_180 ;
	7'h1a :
		TR_114 = RG_rl_180 ;
	7'h1b :
		TR_114 = RG_rl_180 ;
	7'h1c :
		TR_114 = RG_rl_180 ;
	7'h1d :
		TR_114 = RG_rl_180 ;
	7'h1e :
		TR_114 = RG_rl_180 ;
	7'h1f :
		TR_114 = RG_rl_180 ;
	7'h20 :
		TR_114 = RG_rl_180 ;
	7'h21 :
		TR_114 = RG_rl_180 ;
	7'h22 :
		TR_114 = RG_rl_180 ;
	7'h23 :
		TR_114 = RG_rl_180 ;
	7'h24 :
		TR_114 = RG_rl_180 ;
	7'h25 :
		TR_114 = RG_rl_180 ;
	7'h26 :
		TR_114 = RG_rl_180 ;
	7'h27 :
		TR_114 = RG_rl_180 ;
	7'h28 :
		TR_114 = RG_rl_180 ;
	7'h29 :
		TR_114 = RG_rl_180 ;
	7'h2a :
		TR_114 = RG_rl_180 ;
	7'h2b :
		TR_114 = RG_rl_180 ;
	7'h2c :
		TR_114 = RG_rl_180 ;
	7'h2d :
		TR_114 = RG_rl_180 ;
	7'h2e :
		TR_114 = RG_rl_180 ;
	7'h2f :
		TR_114 = RG_rl_180 ;
	7'h30 :
		TR_114 = RG_rl_180 ;
	7'h31 :
		TR_114 = RG_rl_180 ;
	7'h32 :
		TR_114 = RG_rl_180 ;
	7'h33 :
		TR_114 = RG_rl_180 ;
	7'h34 :
		TR_114 = RG_rl_180 ;
	7'h35 :
		TR_114 = RG_rl_180 ;
	7'h36 :
		TR_114 = RG_rl_180 ;
	7'h37 :
		TR_114 = RG_rl_180 ;
	7'h38 :
		TR_114 = RG_rl_180 ;
	7'h39 :
		TR_114 = RG_rl_180 ;
	7'h3a :
		TR_114 = RG_rl_180 ;
	7'h3b :
		TR_114 = RG_rl_180 ;
	7'h3c :
		TR_114 = RG_rl_180 ;
	7'h3d :
		TR_114 = RG_rl_180 ;
	7'h3e :
		TR_114 = RG_rl_180 ;
	7'h3f :
		TR_114 = RG_rl_180 ;
	7'h40 :
		TR_114 = RG_rl_180 ;
	7'h41 :
		TR_114 = RG_rl_180 ;
	7'h42 :
		TR_114 = RG_rl_180 ;
	7'h43 :
		TR_114 = RG_rl_180 ;
	7'h44 :
		TR_114 = RG_rl_180 ;
	7'h45 :
		TR_114 = RG_rl_180 ;
	7'h46 :
		TR_114 = RG_rl_180 ;
	7'h47 :
		TR_114 = RG_rl_180 ;
	7'h48 :
		TR_114 = RG_rl_180 ;
	7'h49 :
		TR_114 = RG_rl_180 ;
	7'h4a :
		TR_114 = RG_rl_180 ;
	7'h4b :
		TR_114 = RG_rl_180 ;
	7'h4c :
		TR_114 = RG_rl_180 ;
	7'h4d :
		TR_114 = RG_rl_180 ;
	7'h4e :
		TR_114 = RG_rl_180 ;
	7'h4f :
		TR_114 = RG_rl_180 ;
	7'h50 :
		TR_114 = RG_rl_180 ;
	7'h51 :
		TR_114 = RG_rl_180 ;
	7'h52 :
		TR_114 = RG_rl_180 ;
	7'h53 :
		TR_114 = RG_rl_180 ;
	7'h54 :
		TR_114 = RG_rl_180 ;
	7'h55 :
		TR_114 = RG_rl_180 ;
	7'h56 :
		TR_114 = RG_rl_180 ;
	7'h57 :
		TR_114 = RG_rl_180 ;
	7'h58 :
		TR_114 = RG_rl_180 ;
	7'h59 :
		TR_114 = RG_rl_180 ;
	7'h5a :
		TR_114 = RG_rl_180 ;
	7'h5b :
		TR_114 = RG_rl_180 ;
	7'h5c :
		TR_114 = RG_rl_180 ;
	7'h5d :
		TR_114 = RG_rl_180 ;
	7'h5e :
		TR_114 = RG_rl_180 ;
	7'h5f :
		TR_114 = RG_rl_180 ;
	7'h60 :
		TR_114 = RG_rl_180 ;
	7'h61 :
		TR_114 = RG_rl_180 ;
	7'h62 :
		TR_114 = RG_rl_180 ;
	7'h63 :
		TR_114 = RG_rl_180 ;
	7'h64 :
		TR_114 = RG_rl_180 ;
	7'h65 :
		TR_114 = RG_rl_180 ;
	7'h66 :
		TR_114 = 9'h000 ;	// line#=../rle.cpp:79
	7'h67 :
		TR_114 = RG_rl_180 ;
	7'h68 :
		TR_114 = RG_rl_180 ;
	7'h69 :
		TR_114 = RG_rl_180 ;
	7'h6a :
		TR_114 = RG_rl_180 ;
	7'h6b :
		TR_114 = RG_rl_180 ;
	7'h6c :
		TR_114 = RG_rl_180 ;
	7'h6d :
		TR_114 = RG_rl_180 ;
	7'h6e :
		TR_114 = RG_rl_180 ;
	7'h6f :
		TR_114 = RG_rl_180 ;
	7'h70 :
		TR_114 = RG_rl_180 ;
	7'h71 :
		TR_114 = RG_rl_180 ;
	7'h72 :
		TR_114 = RG_rl_180 ;
	7'h73 :
		TR_114 = RG_rl_180 ;
	7'h74 :
		TR_114 = RG_rl_180 ;
	7'h75 :
		TR_114 = RG_rl_180 ;
	7'h76 :
		TR_114 = RG_rl_180 ;
	7'h77 :
		TR_114 = RG_rl_180 ;
	7'h78 :
		TR_114 = RG_rl_180 ;
	7'h79 :
		TR_114 = RG_rl_180 ;
	7'h7a :
		TR_114 = RG_rl_180 ;
	7'h7b :
		TR_114 = RG_rl_180 ;
	7'h7c :
		TR_114 = RG_rl_180 ;
	7'h7d :
		TR_114 = RG_rl_180 ;
	7'h7e :
		TR_114 = RG_rl_180 ;
	7'h7f :
		TR_114 = RG_rl_180 ;
	default :
		TR_114 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_49 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h01 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h02 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h03 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h04 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h05 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h06 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h07 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h08 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h09 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h0a :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h0b :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h0c :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h0d :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h0e :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h0f :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h10 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h11 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h12 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h13 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h14 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h15 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h16 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h17 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h18 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h19 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h1a :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h1b :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h1c :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h1d :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h1e :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h1f :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h20 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h21 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h22 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h23 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h24 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h25 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h26 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h27 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h28 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h29 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h2a :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h2b :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h2c :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h2d :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h2e :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h2f :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h30 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h31 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h32 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h33 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h34 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h35 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h36 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h37 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h38 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h39 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h3a :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h3b :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h3c :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h3d :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h3e :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h3f :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h40 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h41 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h42 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h43 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h44 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h45 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h46 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h47 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h48 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h49 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h4a :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h4b :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h4c :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h4d :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h4e :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h4f :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h50 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h51 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h52 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h53 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h54 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h55 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h56 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h57 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h58 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h59 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h5a :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h5b :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h5c :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h5d :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h5e :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h5f :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h60 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h61 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h62 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h63 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h64 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h65 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h66 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h67 :
		TR_115 = 9'h000 ;	// line#=../rle.cpp:79
	7'h68 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h69 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h6a :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h6b :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h6c :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h6d :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h6e :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h6f :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h70 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h71 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h72 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h73 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h74 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h75 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h76 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h77 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h78 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h79 :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h7a :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h7b :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h7c :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h7d :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h7e :
		TR_115 = RG_quantized_block_rl_49 ;
	7'h7f :
		TR_115 = RG_quantized_block_rl_49 ;
	default :
		TR_115 = 9'hx ;
	endcase
always @ ( RG_rl_181 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_116 = RG_rl_181 ;
	7'h01 :
		TR_116 = RG_rl_181 ;
	7'h02 :
		TR_116 = RG_rl_181 ;
	7'h03 :
		TR_116 = RG_rl_181 ;
	7'h04 :
		TR_116 = RG_rl_181 ;
	7'h05 :
		TR_116 = RG_rl_181 ;
	7'h06 :
		TR_116 = RG_rl_181 ;
	7'h07 :
		TR_116 = RG_rl_181 ;
	7'h08 :
		TR_116 = RG_rl_181 ;
	7'h09 :
		TR_116 = RG_rl_181 ;
	7'h0a :
		TR_116 = RG_rl_181 ;
	7'h0b :
		TR_116 = RG_rl_181 ;
	7'h0c :
		TR_116 = RG_rl_181 ;
	7'h0d :
		TR_116 = RG_rl_181 ;
	7'h0e :
		TR_116 = RG_rl_181 ;
	7'h0f :
		TR_116 = RG_rl_181 ;
	7'h10 :
		TR_116 = RG_rl_181 ;
	7'h11 :
		TR_116 = RG_rl_181 ;
	7'h12 :
		TR_116 = RG_rl_181 ;
	7'h13 :
		TR_116 = RG_rl_181 ;
	7'h14 :
		TR_116 = RG_rl_181 ;
	7'h15 :
		TR_116 = RG_rl_181 ;
	7'h16 :
		TR_116 = RG_rl_181 ;
	7'h17 :
		TR_116 = RG_rl_181 ;
	7'h18 :
		TR_116 = RG_rl_181 ;
	7'h19 :
		TR_116 = RG_rl_181 ;
	7'h1a :
		TR_116 = RG_rl_181 ;
	7'h1b :
		TR_116 = RG_rl_181 ;
	7'h1c :
		TR_116 = RG_rl_181 ;
	7'h1d :
		TR_116 = RG_rl_181 ;
	7'h1e :
		TR_116 = RG_rl_181 ;
	7'h1f :
		TR_116 = RG_rl_181 ;
	7'h20 :
		TR_116 = RG_rl_181 ;
	7'h21 :
		TR_116 = RG_rl_181 ;
	7'h22 :
		TR_116 = RG_rl_181 ;
	7'h23 :
		TR_116 = RG_rl_181 ;
	7'h24 :
		TR_116 = RG_rl_181 ;
	7'h25 :
		TR_116 = RG_rl_181 ;
	7'h26 :
		TR_116 = RG_rl_181 ;
	7'h27 :
		TR_116 = RG_rl_181 ;
	7'h28 :
		TR_116 = RG_rl_181 ;
	7'h29 :
		TR_116 = RG_rl_181 ;
	7'h2a :
		TR_116 = RG_rl_181 ;
	7'h2b :
		TR_116 = RG_rl_181 ;
	7'h2c :
		TR_116 = RG_rl_181 ;
	7'h2d :
		TR_116 = RG_rl_181 ;
	7'h2e :
		TR_116 = RG_rl_181 ;
	7'h2f :
		TR_116 = RG_rl_181 ;
	7'h30 :
		TR_116 = RG_rl_181 ;
	7'h31 :
		TR_116 = RG_rl_181 ;
	7'h32 :
		TR_116 = RG_rl_181 ;
	7'h33 :
		TR_116 = RG_rl_181 ;
	7'h34 :
		TR_116 = RG_rl_181 ;
	7'h35 :
		TR_116 = RG_rl_181 ;
	7'h36 :
		TR_116 = RG_rl_181 ;
	7'h37 :
		TR_116 = RG_rl_181 ;
	7'h38 :
		TR_116 = RG_rl_181 ;
	7'h39 :
		TR_116 = RG_rl_181 ;
	7'h3a :
		TR_116 = RG_rl_181 ;
	7'h3b :
		TR_116 = RG_rl_181 ;
	7'h3c :
		TR_116 = RG_rl_181 ;
	7'h3d :
		TR_116 = RG_rl_181 ;
	7'h3e :
		TR_116 = RG_rl_181 ;
	7'h3f :
		TR_116 = RG_rl_181 ;
	7'h40 :
		TR_116 = RG_rl_181 ;
	7'h41 :
		TR_116 = RG_rl_181 ;
	7'h42 :
		TR_116 = RG_rl_181 ;
	7'h43 :
		TR_116 = RG_rl_181 ;
	7'h44 :
		TR_116 = RG_rl_181 ;
	7'h45 :
		TR_116 = RG_rl_181 ;
	7'h46 :
		TR_116 = RG_rl_181 ;
	7'h47 :
		TR_116 = RG_rl_181 ;
	7'h48 :
		TR_116 = RG_rl_181 ;
	7'h49 :
		TR_116 = RG_rl_181 ;
	7'h4a :
		TR_116 = RG_rl_181 ;
	7'h4b :
		TR_116 = RG_rl_181 ;
	7'h4c :
		TR_116 = RG_rl_181 ;
	7'h4d :
		TR_116 = RG_rl_181 ;
	7'h4e :
		TR_116 = RG_rl_181 ;
	7'h4f :
		TR_116 = RG_rl_181 ;
	7'h50 :
		TR_116 = RG_rl_181 ;
	7'h51 :
		TR_116 = RG_rl_181 ;
	7'h52 :
		TR_116 = RG_rl_181 ;
	7'h53 :
		TR_116 = RG_rl_181 ;
	7'h54 :
		TR_116 = RG_rl_181 ;
	7'h55 :
		TR_116 = RG_rl_181 ;
	7'h56 :
		TR_116 = RG_rl_181 ;
	7'h57 :
		TR_116 = RG_rl_181 ;
	7'h58 :
		TR_116 = RG_rl_181 ;
	7'h59 :
		TR_116 = RG_rl_181 ;
	7'h5a :
		TR_116 = RG_rl_181 ;
	7'h5b :
		TR_116 = RG_rl_181 ;
	7'h5c :
		TR_116 = RG_rl_181 ;
	7'h5d :
		TR_116 = RG_rl_181 ;
	7'h5e :
		TR_116 = RG_rl_181 ;
	7'h5f :
		TR_116 = RG_rl_181 ;
	7'h60 :
		TR_116 = RG_rl_181 ;
	7'h61 :
		TR_116 = RG_rl_181 ;
	7'h62 :
		TR_116 = RG_rl_181 ;
	7'h63 :
		TR_116 = RG_rl_181 ;
	7'h64 :
		TR_116 = RG_rl_181 ;
	7'h65 :
		TR_116 = RG_rl_181 ;
	7'h66 :
		TR_116 = RG_rl_181 ;
	7'h67 :
		TR_116 = RG_rl_181 ;
	7'h68 :
		TR_116 = 9'h000 ;	// line#=../rle.cpp:79
	7'h69 :
		TR_116 = RG_rl_181 ;
	7'h6a :
		TR_116 = RG_rl_181 ;
	7'h6b :
		TR_116 = RG_rl_181 ;
	7'h6c :
		TR_116 = RG_rl_181 ;
	7'h6d :
		TR_116 = RG_rl_181 ;
	7'h6e :
		TR_116 = RG_rl_181 ;
	7'h6f :
		TR_116 = RG_rl_181 ;
	7'h70 :
		TR_116 = RG_rl_181 ;
	7'h71 :
		TR_116 = RG_rl_181 ;
	7'h72 :
		TR_116 = RG_rl_181 ;
	7'h73 :
		TR_116 = RG_rl_181 ;
	7'h74 :
		TR_116 = RG_rl_181 ;
	7'h75 :
		TR_116 = RG_rl_181 ;
	7'h76 :
		TR_116 = RG_rl_181 ;
	7'h77 :
		TR_116 = RG_rl_181 ;
	7'h78 :
		TR_116 = RG_rl_181 ;
	7'h79 :
		TR_116 = RG_rl_181 ;
	7'h7a :
		TR_116 = RG_rl_181 ;
	7'h7b :
		TR_116 = RG_rl_181 ;
	7'h7c :
		TR_116 = RG_rl_181 ;
	7'h7d :
		TR_116 = RG_rl_181 ;
	7'h7e :
		TR_116 = RG_rl_181 ;
	7'h7f :
		TR_116 = RG_rl_181 ;
	default :
		TR_116 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_50 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h01 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h02 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h03 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h04 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h05 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h06 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h07 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h08 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h09 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h0a :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h0b :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h0c :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h0d :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h0e :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h0f :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h10 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h11 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h12 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h13 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h14 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h15 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h16 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h17 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h18 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h19 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h1a :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h1b :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h1c :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h1d :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h1e :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h1f :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h20 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h21 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h22 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h23 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h24 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h25 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h26 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h27 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h28 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h29 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h2a :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h2b :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h2c :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h2d :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h2e :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h2f :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h30 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h31 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h32 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h33 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h34 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h35 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h36 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h37 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h38 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h39 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h3a :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h3b :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h3c :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h3d :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h3e :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h3f :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h40 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h41 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h42 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h43 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h44 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h45 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h46 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h47 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h48 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h49 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h4a :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h4b :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h4c :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h4d :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h4e :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h4f :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h50 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h51 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h52 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h53 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h54 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h55 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h56 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h57 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h58 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h59 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h5a :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h5b :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h5c :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h5d :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h5e :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h5f :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h60 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h61 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h62 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h63 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h64 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h65 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h66 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h67 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h68 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h69 :
		TR_117 = 9'h000 ;	// line#=../rle.cpp:79
	7'h6a :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h6b :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h6c :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h6d :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h6e :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h6f :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h70 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h71 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h72 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h73 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h74 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h75 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h76 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h77 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h78 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h79 :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h7a :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h7b :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h7c :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h7d :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h7e :
		TR_117 = RG_quantized_block_rl_50 ;
	7'h7f :
		TR_117 = RG_quantized_block_rl_50 ;
	default :
		TR_117 = 9'hx ;
	endcase
always @ ( RG_rl_182 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_118 = RG_rl_182 ;
	7'h01 :
		TR_118 = RG_rl_182 ;
	7'h02 :
		TR_118 = RG_rl_182 ;
	7'h03 :
		TR_118 = RG_rl_182 ;
	7'h04 :
		TR_118 = RG_rl_182 ;
	7'h05 :
		TR_118 = RG_rl_182 ;
	7'h06 :
		TR_118 = RG_rl_182 ;
	7'h07 :
		TR_118 = RG_rl_182 ;
	7'h08 :
		TR_118 = RG_rl_182 ;
	7'h09 :
		TR_118 = RG_rl_182 ;
	7'h0a :
		TR_118 = RG_rl_182 ;
	7'h0b :
		TR_118 = RG_rl_182 ;
	7'h0c :
		TR_118 = RG_rl_182 ;
	7'h0d :
		TR_118 = RG_rl_182 ;
	7'h0e :
		TR_118 = RG_rl_182 ;
	7'h0f :
		TR_118 = RG_rl_182 ;
	7'h10 :
		TR_118 = RG_rl_182 ;
	7'h11 :
		TR_118 = RG_rl_182 ;
	7'h12 :
		TR_118 = RG_rl_182 ;
	7'h13 :
		TR_118 = RG_rl_182 ;
	7'h14 :
		TR_118 = RG_rl_182 ;
	7'h15 :
		TR_118 = RG_rl_182 ;
	7'h16 :
		TR_118 = RG_rl_182 ;
	7'h17 :
		TR_118 = RG_rl_182 ;
	7'h18 :
		TR_118 = RG_rl_182 ;
	7'h19 :
		TR_118 = RG_rl_182 ;
	7'h1a :
		TR_118 = RG_rl_182 ;
	7'h1b :
		TR_118 = RG_rl_182 ;
	7'h1c :
		TR_118 = RG_rl_182 ;
	7'h1d :
		TR_118 = RG_rl_182 ;
	7'h1e :
		TR_118 = RG_rl_182 ;
	7'h1f :
		TR_118 = RG_rl_182 ;
	7'h20 :
		TR_118 = RG_rl_182 ;
	7'h21 :
		TR_118 = RG_rl_182 ;
	7'h22 :
		TR_118 = RG_rl_182 ;
	7'h23 :
		TR_118 = RG_rl_182 ;
	7'h24 :
		TR_118 = RG_rl_182 ;
	7'h25 :
		TR_118 = RG_rl_182 ;
	7'h26 :
		TR_118 = RG_rl_182 ;
	7'h27 :
		TR_118 = RG_rl_182 ;
	7'h28 :
		TR_118 = RG_rl_182 ;
	7'h29 :
		TR_118 = RG_rl_182 ;
	7'h2a :
		TR_118 = RG_rl_182 ;
	7'h2b :
		TR_118 = RG_rl_182 ;
	7'h2c :
		TR_118 = RG_rl_182 ;
	7'h2d :
		TR_118 = RG_rl_182 ;
	7'h2e :
		TR_118 = RG_rl_182 ;
	7'h2f :
		TR_118 = RG_rl_182 ;
	7'h30 :
		TR_118 = RG_rl_182 ;
	7'h31 :
		TR_118 = RG_rl_182 ;
	7'h32 :
		TR_118 = RG_rl_182 ;
	7'h33 :
		TR_118 = RG_rl_182 ;
	7'h34 :
		TR_118 = RG_rl_182 ;
	7'h35 :
		TR_118 = RG_rl_182 ;
	7'h36 :
		TR_118 = RG_rl_182 ;
	7'h37 :
		TR_118 = RG_rl_182 ;
	7'h38 :
		TR_118 = RG_rl_182 ;
	7'h39 :
		TR_118 = RG_rl_182 ;
	7'h3a :
		TR_118 = RG_rl_182 ;
	7'h3b :
		TR_118 = RG_rl_182 ;
	7'h3c :
		TR_118 = RG_rl_182 ;
	7'h3d :
		TR_118 = RG_rl_182 ;
	7'h3e :
		TR_118 = RG_rl_182 ;
	7'h3f :
		TR_118 = RG_rl_182 ;
	7'h40 :
		TR_118 = RG_rl_182 ;
	7'h41 :
		TR_118 = RG_rl_182 ;
	7'h42 :
		TR_118 = RG_rl_182 ;
	7'h43 :
		TR_118 = RG_rl_182 ;
	7'h44 :
		TR_118 = RG_rl_182 ;
	7'h45 :
		TR_118 = RG_rl_182 ;
	7'h46 :
		TR_118 = RG_rl_182 ;
	7'h47 :
		TR_118 = RG_rl_182 ;
	7'h48 :
		TR_118 = RG_rl_182 ;
	7'h49 :
		TR_118 = RG_rl_182 ;
	7'h4a :
		TR_118 = RG_rl_182 ;
	7'h4b :
		TR_118 = RG_rl_182 ;
	7'h4c :
		TR_118 = RG_rl_182 ;
	7'h4d :
		TR_118 = RG_rl_182 ;
	7'h4e :
		TR_118 = RG_rl_182 ;
	7'h4f :
		TR_118 = RG_rl_182 ;
	7'h50 :
		TR_118 = RG_rl_182 ;
	7'h51 :
		TR_118 = RG_rl_182 ;
	7'h52 :
		TR_118 = RG_rl_182 ;
	7'h53 :
		TR_118 = RG_rl_182 ;
	7'h54 :
		TR_118 = RG_rl_182 ;
	7'h55 :
		TR_118 = RG_rl_182 ;
	7'h56 :
		TR_118 = RG_rl_182 ;
	7'h57 :
		TR_118 = RG_rl_182 ;
	7'h58 :
		TR_118 = RG_rl_182 ;
	7'h59 :
		TR_118 = RG_rl_182 ;
	7'h5a :
		TR_118 = RG_rl_182 ;
	7'h5b :
		TR_118 = RG_rl_182 ;
	7'h5c :
		TR_118 = RG_rl_182 ;
	7'h5d :
		TR_118 = RG_rl_182 ;
	7'h5e :
		TR_118 = RG_rl_182 ;
	7'h5f :
		TR_118 = RG_rl_182 ;
	7'h60 :
		TR_118 = RG_rl_182 ;
	7'h61 :
		TR_118 = RG_rl_182 ;
	7'h62 :
		TR_118 = RG_rl_182 ;
	7'h63 :
		TR_118 = RG_rl_182 ;
	7'h64 :
		TR_118 = RG_rl_182 ;
	7'h65 :
		TR_118 = RG_rl_182 ;
	7'h66 :
		TR_118 = RG_rl_182 ;
	7'h67 :
		TR_118 = RG_rl_182 ;
	7'h68 :
		TR_118 = RG_rl_182 ;
	7'h69 :
		TR_118 = RG_rl_182 ;
	7'h6a :
		TR_118 = 9'h000 ;	// line#=../rle.cpp:79
	7'h6b :
		TR_118 = RG_rl_182 ;
	7'h6c :
		TR_118 = RG_rl_182 ;
	7'h6d :
		TR_118 = RG_rl_182 ;
	7'h6e :
		TR_118 = RG_rl_182 ;
	7'h6f :
		TR_118 = RG_rl_182 ;
	7'h70 :
		TR_118 = RG_rl_182 ;
	7'h71 :
		TR_118 = RG_rl_182 ;
	7'h72 :
		TR_118 = RG_rl_182 ;
	7'h73 :
		TR_118 = RG_rl_182 ;
	7'h74 :
		TR_118 = RG_rl_182 ;
	7'h75 :
		TR_118 = RG_rl_182 ;
	7'h76 :
		TR_118 = RG_rl_182 ;
	7'h77 :
		TR_118 = RG_rl_182 ;
	7'h78 :
		TR_118 = RG_rl_182 ;
	7'h79 :
		TR_118 = RG_rl_182 ;
	7'h7a :
		TR_118 = RG_rl_182 ;
	7'h7b :
		TR_118 = RG_rl_182 ;
	7'h7c :
		TR_118 = RG_rl_182 ;
	7'h7d :
		TR_118 = RG_rl_182 ;
	7'h7e :
		TR_118 = RG_rl_182 ;
	7'h7f :
		TR_118 = RG_rl_182 ;
	default :
		TR_118 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_51 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h01 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h02 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h03 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h04 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h05 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h06 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h07 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h08 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h09 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h0a :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h0b :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h0c :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h0d :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h0e :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h0f :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h10 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h11 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h12 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h13 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h14 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h15 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h16 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h17 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h18 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h19 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h1a :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h1b :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h1c :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h1d :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h1e :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h1f :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h20 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h21 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h22 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h23 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h24 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h25 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h26 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h27 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h28 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h29 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h2a :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h2b :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h2c :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h2d :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h2e :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h2f :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h30 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h31 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h32 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h33 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h34 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h35 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h36 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h37 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h38 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h39 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h3a :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h3b :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h3c :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h3d :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h3e :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h3f :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h40 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h41 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h42 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h43 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h44 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h45 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h46 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h47 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h48 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h49 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h4a :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h4b :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h4c :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h4d :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h4e :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h4f :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h50 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h51 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h52 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h53 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h54 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h55 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h56 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h57 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h58 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h59 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h5a :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h5b :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h5c :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h5d :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h5e :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h5f :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h60 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h61 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h62 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h63 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h64 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h65 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h66 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h67 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h68 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h69 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h6a :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h6b :
		TR_119 = 9'h000 ;	// line#=../rle.cpp:79
	7'h6c :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h6d :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h6e :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h6f :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h70 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h71 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h72 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h73 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h74 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h75 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h76 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h77 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h78 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h79 :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h7a :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h7b :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h7c :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h7d :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h7e :
		TR_119 = RG_quantized_block_rl_51 ;
	7'h7f :
		TR_119 = RG_quantized_block_rl_51 ;
	default :
		TR_119 = 9'hx ;
	endcase
always @ ( RG_rl_183 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_120 = RG_rl_183 ;
	7'h01 :
		TR_120 = RG_rl_183 ;
	7'h02 :
		TR_120 = RG_rl_183 ;
	7'h03 :
		TR_120 = RG_rl_183 ;
	7'h04 :
		TR_120 = RG_rl_183 ;
	7'h05 :
		TR_120 = RG_rl_183 ;
	7'h06 :
		TR_120 = RG_rl_183 ;
	7'h07 :
		TR_120 = RG_rl_183 ;
	7'h08 :
		TR_120 = RG_rl_183 ;
	7'h09 :
		TR_120 = RG_rl_183 ;
	7'h0a :
		TR_120 = RG_rl_183 ;
	7'h0b :
		TR_120 = RG_rl_183 ;
	7'h0c :
		TR_120 = RG_rl_183 ;
	7'h0d :
		TR_120 = RG_rl_183 ;
	7'h0e :
		TR_120 = RG_rl_183 ;
	7'h0f :
		TR_120 = RG_rl_183 ;
	7'h10 :
		TR_120 = RG_rl_183 ;
	7'h11 :
		TR_120 = RG_rl_183 ;
	7'h12 :
		TR_120 = RG_rl_183 ;
	7'h13 :
		TR_120 = RG_rl_183 ;
	7'h14 :
		TR_120 = RG_rl_183 ;
	7'h15 :
		TR_120 = RG_rl_183 ;
	7'h16 :
		TR_120 = RG_rl_183 ;
	7'h17 :
		TR_120 = RG_rl_183 ;
	7'h18 :
		TR_120 = RG_rl_183 ;
	7'h19 :
		TR_120 = RG_rl_183 ;
	7'h1a :
		TR_120 = RG_rl_183 ;
	7'h1b :
		TR_120 = RG_rl_183 ;
	7'h1c :
		TR_120 = RG_rl_183 ;
	7'h1d :
		TR_120 = RG_rl_183 ;
	7'h1e :
		TR_120 = RG_rl_183 ;
	7'h1f :
		TR_120 = RG_rl_183 ;
	7'h20 :
		TR_120 = RG_rl_183 ;
	7'h21 :
		TR_120 = RG_rl_183 ;
	7'h22 :
		TR_120 = RG_rl_183 ;
	7'h23 :
		TR_120 = RG_rl_183 ;
	7'h24 :
		TR_120 = RG_rl_183 ;
	7'h25 :
		TR_120 = RG_rl_183 ;
	7'h26 :
		TR_120 = RG_rl_183 ;
	7'h27 :
		TR_120 = RG_rl_183 ;
	7'h28 :
		TR_120 = RG_rl_183 ;
	7'h29 :
		TR_120 = RG_rl_183 ;
	7'h2a :
		TR_120 = RG_rl_183 ;
	7'h2b :
		TR_120 = RG_rl_183 ;
	7'h2c :
		TR_120 = RG_rl_183 ;
	7'h2d :
		TR_120 = RG_rl_183 ;
	7'h2e :
		TR_120 = RG_rl_183 ;
	7'h2f :
		TR_120 = RG_rl_183 ;
	7'h30 :
		TR_120 = RG_rl_183 ;
	7'h31 :
		TR_120 = RG_rl_183 ;
	7'h32 :
		TR_120 = RG_rl_183 ;
	7'h33 :
		TR_120 = RG_rl_183 ;
	7'h34 :
		TR_120 = RG_rl_183 ;
	7'h35 :
		TR_120 = RG_rl_183 ;
	7'h36 :
		TR_120 = RG_rl_183 ;
	7'h37 :
		TR_120 = RG_rl_183 ;
	7'h38 :
		TR_120 = RG_rl_183 ;
	7'h39 :
		TR_120 = RG_rl_183 ;
	7'h3a :
		TR_120 = RG_rl_183 ;
	7'h3b :
		TR_120 = RG_rl_183 ;
	7'h3c :
		TR_120 = RG_rl_183 ;
	7'h3d :
		TR_120 = RG_rl_183 ;
	7'h3e :
		TR_120 = RG_rl_183 ;
	7'h3f :
		TR_120 = RG_rl_183 ;
	7'h40 :
		TR_120 = RG_rl_183 ;
	7'h41 :
		TR_120 = RG_rl_183 ;
	7'h42 :
		TR_120 = RG_rl_183 ;
	7'h43 :
		TR_120 = RG_rl_183 ;
	7'h44 :
		TR_120 = RG_rl_183 ;
	7'h45 :
		TR_120 = RG_rl_183 ;
	7'h46 :
		TR_120 = RG_rl_183 ;
	7'h47 :
		TR_120 = RG_rl_183 ;
	7'h48 :
		TR_120 = RG_rl_183 ;
	7'h49 :
		TR_120 = RG_rl_183 ;
	7'h4a :
		TR_120 = RG_rl_183 ;
	7'h4b :
		TR_120 = RG_rl_183 ;
	7'h4c :
		TR_120 = RG_rl_183 ;
	7'h4d :
		TR_120 = RG_rl_183 ;
	7'h4e :
		TR_120 = RG_rl_183 ;
	7'h4f :
		TR_120 = RG_rl_183 ;
	7'h50 :
		TR_120 = RG_rl_183 ;
	7'h51 :
		TR_120 = RG_rl_183 ;
	7'h52 :
		TR_120 = RG_rl_183 ;
	7'h53 :
		TR_120 = RG_rl_183 ;
	7'h54 :
		TR_120 = RG_rl_183 ;
	7'h55 :
		TR_120 = RG_rl_183 ;
	7'h56 :
		TR_120 = RG_rl_183 ;
	7'h57 :
		TR_120 = RG_rl_183 ;
	7'h58 :
		TR_120 = RG_rl_183 ;
	7'h59 :
		TR_120 = RG_rl_183 ;
	7'h5a :
		TR_120 = RG_rl_183 ;
	7'h5b :
		TR_120 = RG_rl_183 ;
	7'h5c :
		TR_120 = RG_rl_183 ;
	7'h5d :
		TR_120 = RG_rl_183 ;
	7'h5e :
		TR_120 = RG_rl_183 ;
	7'h5f :
		TR_120 = RG_rl_183 ;
	7'h60 :
		TR_120 = RG_rl_183 ;
	7'h61 :
		TR_120 = RG_rl_183 ;
	7'h62 :
		TR_120 = RG_rl_183 ;
	7'h63 :
		TR_120 = RG_rl_183 ;
	7'h64 :
		TR_120 = RG_rl_183 ;
	7'h65 :
		TR_120 = RG_rl_183 ;
	7'h66 :
		TR_120 = RG_rl_183 ;
	7'h67 :
		TR_120 = RG_rl_183 ;
	7'h68 :
		TR_120 = RG_rl_183 ;
	7'h69 :
		TR_120 = RG_rl_183 ;
	7'h6a :
		TR_120 = RG_rl_183 ;
	7'h6b :
		TR_120 = RG_rl_183 ;
	7'h6c :
		TR_120 = 9'h000 ;	// line#=../rle.cpp:79
	7'h6d :
		TR_120 = RG_rl_183 ;
	7'h6e :
		TR_120 = RG_rl_183 ;
	7'h6f :
		TR_120 = RG_rl_183 ;
	7'h70 :
		TR_120 = RG_rl_183 ;
	7'h71 :
		TR_120 = RG_rl_183 ;
	7'h72 :
		TR_120 = RG_rl_183 ;
	7'h73 :
		TR_120 = RG_rl_183 ;
	7'h74 :
		TR_120 = RG_rl_183 ;
	7'h75 :
		TR_120 = RG_rl_183 ;
	7'h76 :
		TR_120 = RG_rl_183 ;
	7'h77 :
		TR_120 = RG_rl_183 ;
	7'h78 :
		TR_120 = RG_rl_183 ;
	7'h79 :
		TR_120 = RG_rl_183 ;
	7'h7a :
		TR_120 = RG_rl_183 ;
	7'h7b :
		TR_120 = RG_rl_183 ;
	7'h7c :
		TR_120 = RG_rl_183 ;
	7'h7d :
		TR_120 = RG_rl_183 ;
	7'h7e :
		TR_120 = RG_rl_183 ;
	7'h7f :
		TR_120 = RG_rl_183 ;
	default :
		TR_120 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_52 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h01 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h02 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h03 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h04 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h05 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h06 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h07 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h08 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h09 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h0a :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h0b :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h0c :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h0d :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h0e :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h0f :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h10 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h11 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h12 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h13 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h14 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h15 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h16 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h17 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h18 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h19 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h1a :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h1b :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h1c :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h1d :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h1e :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h1f :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h20 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h21 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h22 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h23 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h24 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h25 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h26 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h27 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h28 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h29 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h2a :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h2b :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h2c :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h2d :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h2e :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h2f :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h30 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h31 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h32 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h33 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h34 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h35 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h36 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h37 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h38 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h39 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h3a :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h3b :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h3c :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h3d :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h3e :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h3f :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h40 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h41 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h42 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h43 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h44 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h45 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h46 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h47 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h48 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h49 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h4a :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h4b :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h4c :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h4d :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h4e :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h4f :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h50 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h51 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h52 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h53 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h54 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h55 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h56 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h57 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h58 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h59 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h5a :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h5b :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h5c :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h5d :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h5e :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h5f :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h60 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h61 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h62 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h63 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h64 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h65 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h66 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h67 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h68 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h69 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h6a :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h6b :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h6c :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h6d :
		TR_121 = 9'h000 ;	// line#=../rle.cpp:79
	7'h6e :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h6f :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h70 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h71 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h72 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h73 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h74 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h75 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h76 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h77 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h78 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h79 :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h7a :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h7b :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h7c :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h7d :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h7e :
		TR_121 = RG_quantized_block_rl_52 ;
	7'h7f :
		TR_121 = RG_quantized_block_rl_52 ;
	default :
		TR_121 = 9'hx ;
	endcase
always @ ( RG_rl_184 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_122 = RG_rl_184 ;
	7'h01 :
		TR_122 = RG_rl_184 ;
	7'h02 :
		TR_122 = RG_rl_184 ;
	7'h03 :
		TR_122 = RG_rl_184 ;
	7'h04 :
		TR_122 = RG_rl_184 ;
	7'h05 :
		TR_122 = RG_rl_184 ;
	7'h06 :
		TR_122 = RG_rl_184 ;
	7'h07 :
		TR_122 = RG_rl_184 ;
	7'h08 :
		TR_122 = RG_rl_184 ;
	7'h09 :
		TR_122 = RG_rl_184 ;
	7'h0a :
		TR_122 = RG_rl_184 ;
	7'h0b :
		TR_122 = RG_rl_184 ;
	7'h0c :
		TR_122 = RG_rl_184 ;
	7'h0d :
		TR_122 = RG_rl_184 ;
	7'h0e :
		TR_122 = RG_rl_184 ;
	7'h0f :
		TR_122 = RG_rl_184 ;
	7'h10 :
		TR_122 = RG_rl_184 ;
	7'h11 :
		TR_122 = RG_rl_184 ;
	7'h12 :
		TR_122 = RG_rl_184 ;
	7'h13 :
		TR_122 = RG_rl_184 ;
	7'h14 :
		TR_122 = RG_rl_184 ;
	7'h15 :
		TR_122 = RG_rl_184 ;
	7'h16 :
		TR_122 = RG_rl_184 ;
	7'h17 :
		TR_122 = RG_rl_184 ;
	7'h18 :
		TR_122 = RG_rl_184 ;
	7'h19 :
		TR_122 = RG_rl_184 ;
	7'h1a :
		TR_122 = RG_rl_184 ;
	7'h1b :
		TR_122 = RG_rl_184 ;
	7'h1c :
		TR_122 = RG_rl_184 ;
	7'h1d :
		TR_122 = RG_rl_184 ;
	7'h1e :
		TR_122 = RG_rl_184 ;
	7'h1f :
		TR_122 = RG_rl_184 ;
	7'h20 :
		TR_122 = RG_rl_184 ;
	7'h21 :
		TR_122 = RG_rl_184 ;
	7'h22 :
		TR_122 = RG_rl_184 ;
	7'h23 :
		TR_122 = RG_rl_184 ;
	7'h24 :
		TR_122 = RG_rl_184 ;
	7'h25 :
		TR_122 = RG_rl_184 ;
	7'h26 :
		TR_122 = RG_rl_184 ;
	7'h27 :
		TR_122 = RG_rl_184 ;
	7'h28 :
		TR_122 = RG_rl_184 ;
	7'h29 :
		TR_122 = RG_rl_184 ;
	7'h2a :
		TR_122 = RG_rl_184 ;
	7'h2b :
		TR_122 = RG_rl_184 ;
	7'h2c :
		TR_122 = RG_rl_184 ;
	7'h2d :
		TR_122 = RG_rl_184 ;
	7'h2e :
		TR_122 = RG_rl_184 ;
	7'h2f :
		TR_122 = RG_rl_184 ;
	7'h30 :
		TR_122 = RG_rl_184 ;
	7'h31 :
		TR_122 = RG_rl_184 ;
	7'h32 :
		TR_122 = RG_rl_184 ;
	7'h33 :
		TR_122 = RG_rl_184 ;
	7'h34 :
		TR_122 = RG_rl_184 ;
	7'h35 :
		TR_122 = RG_rl_184 ;
	7'h36 :
		TR_122 = RG_rl_184 ;
	7'h37 :
		TR_122 = RG_rl_184 ;
	7'h38 :
		TR_122 = RG_rl_184 ;
	7'h39 :
		TR_122 = RG_rl_184 ;
	7'h3a :
		TR_122 = RG_rl_184 ;
	7'h3b :
		TR_122 = RG_rl_184 ;
	7'h3c :
		TR_122 = RG_rl_184 ;
	7'h3d :
		TR_122 = RG_rl_184 ;
	7'h3e :
		TR_122 = RG_rl_184 ;
	7'h3f :
		TR_122 = RG_rl_184 ;
	7'h40 :
		TR_122 = RG_rl_184 ;
	7'h41 :
		TR_122 = RG_rl_184 ;
	7'h42 :
		TR_122 = RG_rl_184 ;
	7'h43 :
		TR_122 = RG_rl_184 ;
	7'h44 :
		TR_122 = RG_rl_184 ;
	7'h45 :
		TR_122 = RG_rl_184 ;
	7'h46 :
		TR_122 = RG_rl_184 ;
	7'h47 :
		TR_122 = RG_rl_184 ;
	7'h48 :
		TR_122 = RG_rl_184 ;
	7'h49 :
		TR_122 = RG_rl_184 ;
	7'h4a :
		TR_122 = RG_rl_184 ;
	7'h4b :
		TR_122 = RG_rl_184 ;
	7'h4c :
		TR_122 = RG_rl_184 ;
	7'h4d :
		TR_122 = RG_rl_184 ;
	7'h4e :
		TR_122 = RG_rl_184 ;
	7'h4f :
		TR_122 = RG_rl_184 ;
	7'h50 :
		TR_122 = RG_rl_184 ;
	7'h51 :
		TR_122 = RG_rl_184 ;
	7'h52 :
		TR_122 = RG_rl_184 ;
	7'h53 :
		TR_122 = RG_rl_184 ;
	7'h54 :
		TR_122 = RG_rl_184 ;
	7'h55 :
		TR_122 = RG_rl_184 ;
	7'h56 :
		TR_122 = RG_rl_184 ;
	7'h57 :
		TR_122 = RG_rl_184 ;
	7'h58 :
		TR_122 = RG_rl_184 ;
	7'h59 :
		TR_122 = RG_rl_184 ;
	7'h5a :
		TR_122 = RG_rl_184 ;
	7'h5b :
		TR_122 = RG_rl_184 ;
	7'h5c :
		TR_122 = RG_rl_184 ;
	7'h5d :
		TR_122 = RG_rl_184 ;
	7'h5e :
		TR_122 = RG_rl_184 ;
	7'h5f :
		TR_122 = RG_rl_184 ;
	7'h60 :
		TR_122 = RG_rl_184 ;
	7'h61 :
		TR_122 = RG_rl_184 ;
	7'h62 :
		TR_122 = RG_rl_184 ;
	7'h63 :
		TR_122 = RG_rl_184 ;
	7'h64 :
		TR_122 = RG_rl_184 ;
	7'h65 :
		TR_122 = RG_rl_184 ;
	7'h66 :
		TR_122 = RG_rl_184 ;
	7'h67 :
		TR_122 = RG_rl_184 ;
	7'h68 :
		TR_122 = RG_rl_184 ;
	7'h69 :
		TR_122 = RG_rl_184 ;
	7'h6a :
		TR_122 = RG_rl_184 ;
	7'h6b :
		TR_122 = RG_rl_184 ;
	7'h6c :
		TR_122 = RG_rl_184 ;
	7'h6d :
		TR_122 = RG_rl_184 ;
	7'h6e :
		TR_122 = 9'h000 ;	// line#=../rle.cpp:79
	7'h6f :
		TR_122 = RG_rl_184 ;
	7'h70 :
		TR_122 = RG_rl_184 ;
	7'h71 :
		TR_122 = RG_rl_184 ;
	7'h72 :
		TR_122 = RG_rl_184 ;
	7'h73 :
		TR_122 = RG_rl_184 ;
	7'h74 :
		TR_122 = RG_rl_184 ;
	7'h75 :
		TR_122 = RG_rl_184 ;
	7'h76 :
		TR_122 = RG_rl_184 ;
	7'h77 :
		TR_122 = RG_rl_184 ;
	7'h78 :
		TR_122 = RG_rl_184 ;
	7'h79 :
		TR_122 = RG_rl_184 ;
	7'h7a :
		TR_122 = RG_rl_184 ;
	7'h7b :
		TR_122 = RG_rl_184 ;
	7'h7c :
		TR_122 = RG_rl_184 ;
	7'h7d :
		TR_122 = RG_rl_184 ;
	7'h7e :
		TR_122 = RG_rl_184 ;
	7'h7f :
		TR_122 = RG_rl_184 ;
	default :
		TR_122 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_53 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h01 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h02 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h03 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h04 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h05 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h06 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h07 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h08 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h09 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h0a :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h0b :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h0c :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h0d :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h0e :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h0f :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h10 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h11 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h12 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h13 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h14 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h15 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h16 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h17 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h18 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h19 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h1a :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h1b :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h1c :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h1d :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h1e :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h1f :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h20 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h21 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h22 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h23 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h24 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h25 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h26 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h27 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h28 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h29 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h2a :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h2b :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h2c :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h2d :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h2e :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h2f :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h30 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h31 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h32 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h33 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h34 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h35 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h36 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h37 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h38 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h39 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h3a :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h3b :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h3c :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h3d :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h3e :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h3f :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h40 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h41 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h42 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h43 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h44 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h45 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h46 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h47 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h48 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h49 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h4a :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h4b :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h4c :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h4d :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h4e :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h4f :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h50 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h51 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h52 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h53 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h54 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h55 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h56 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h57 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h58 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h59 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h5a :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h5b :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h5c :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h5d :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h5e :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h5f :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h60 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h61 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h62 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h63 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h64 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h65 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h66 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h67 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h68 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h69 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h6a :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h6b :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h6c :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h6d :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h6e :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h6f :
		TR_123 = 9'h000 ;	// line#=../rle.cpp:79
	7'h70 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h71 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h72 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h73 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h74 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h75 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h76 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h77 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h78 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h79 :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h7a :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h7b :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h7c :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h7d :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h7e :
		TR_123 = RG_quantized_block_rl_53 ;
	7'h7f :
		TR_123 = RG_quantized_block_rl_53 ;
	default :
		TR_123 = 9'hx ;
	endcase
always @ ( RG_rl_185 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_124 = RG_rl_185 ;
	7'h01 :
		TR_124 = RG_rl_185 ;
	7'h02 :
		TR_124 = RG_rl_185 ;
	7'h03 :
		TR_124 = RG_rl_185 ;
	7'h04 :
		TR_124 = RG_rl_185 ;
	7'h05 :
		TR_124 = RG_rl_185 ;
	7'h06 :
		TR_124 = RG_rl_185 ;
	7'h07 :
		TR_124 = RG_rl_185 ;
	7'h08 :
		TR_124 = RG_rl_185 ;
	7'h09 :
		TR_124 = RG_rl_185 ;
	7'h0a :
		TR_124 = RG_rl_185 ;
	7'h0b :
		TR_124 = RG_rl_185 ;
	7'h0c :
		TR_124 = RG_rl_185 ;
	7'h0d :
		TR_124 = RG_rl_185 ;
	7'h0e :
		TR_124 = RG_rl_185 ;
	7'h0f :
		TR_124 = RG_rl_185 ;
	7'h10 :
		TR_124 = RG_rl_185 ;
	7'h11 :
		TR_124 = RG_rl_185 ;
	7'h12 :
		TR_124 = RG_rl_185 ;
	7'h13 :
		TR_124 = RG_rl_185 ;
	7'h14 :
		TR_124 = RG_rl_185 ;
	7'h15 :
		TR_124 = RG_rl_185 ;
	7'h16 :
		TR_124 = RG_rl_185 ;
	7'h17 :
		TR_124 = RG_rl_185 ;
	7'h18 :
		TR_124 = RG_rl_185 ;
	7'h19 :
		TR_124 = RG_rl_185 ;
	7'h1a :
		TR_124 = RG_rl_185 ;
	7'h1b :
		TR_124 = RG_rl_185 ;
	7'h1c :
		TR_124 = RG_rl_185 ;
	7'h1d :
		TR_124 = RG_rl_185 ;
	7'h1e :
		TR_124 = RG_rl_185 ;
	7'h1f :
		TR_124 = RG_rl_185 ;
	7'h20 :
		TR_124 = RG_rl_185 ;
	7'h21 :
		TR_124 = RG_rl_185 ;
	7'h22 :
		TR_124 = RG_rl_185 ;
	7'h23 :
		TR_124 = RG_rl_185 ;
	7'h24 :
		TR_124 = RG_rl_185 ;
	7'h25 :
		TR_124 = RG_rl_185 ;
	7'h26 :
		TR_124 = RG_rl_185 ;
	7'h27 :
		TR_124 = RG_rl_185 ;
	7'h28 :
		TR_124 = RG_rl_185 ;
	7'h29 :
		TR_124 = RG_rl_185 ;
	7'h2a :
		TR_124 = RG_rl_185 ;
	7'h2b :
		TR_124 = RG_rl_185 ;
	7'h2c :
		TR_124 = RG_rl_185 ;
	7'h2d :
		TR_124 = RG_rl_185 ;
	7'h2e :
		TR_124 = RG_rl_185 ;
	7'h2f :
		TR_124 = RG_rl_185 ;
	7'h30 :
		TR_124 = RG_rl_185 ;
	7'h31 :
		TR_124 = RG_rl_185 ;
	7'h32 :
		TR_124 = RG_rl_185 ;
	7'h33 :
		TR_124 = RG_rl_185 ;
	7'h34 :
		TR_124 = RG_rl_185 ;
	7'h35 :
		TR_124 = RG_rl_185 ;
	7'h36 :
		TR_124 = RG_rl_185 ;
	7'h37 :
		TR_124 = RG_rl_185 ;
	7'h38 :
		TR_124 = RG_rl_185 ;
	7'h39 :
		TR_124 = RG_rl_185 ;
	7'h3a :
		TR_124 = RG_rl_185 ;
	7'h3b :
		TR_124 = RG_rl_185 ;
	7'h3c :
		TR_124 = RG_rl_185 ;
	7'h3d :
		TR_124 = RG_rl_185 ;
	7'h3e :
		TR_124 = RG_rl_185 ;
	7'h3f :
		TR_124 = RG_rl_185 ;
	7'h40 :
		TR_124 = RG_rl_185 ;
	7'h41 :
		TR_124 = RG_rl_185 ;
	7'h42 :
		TR_124 = RG_rl_185 ;
	7'h43 :
		TR_124 = RG_rl_185 ;
	7'h44 :
		TR_124 = RG_rl_185 ;
	7'h45 :
		TR_124 = RG_rl_185 ;
	7'h46 :
		TR_124 = RG_rl_185 ;
	7'h47 :
		TR_124 = RG_rl_185 ;
	7'h48 :
		TR_124 = RG_rl_185 ;
	7'h49 :
		TR_124 = RG_rl_185 ;
	7'h4a :
		TR_124 = RG_rl_185 ;
	7'h4b :
		TR_124 = RG_rl_185 ;
	7'h4c :
		TR_124 = RG_rl_185 ;
	7'h4d :
		TR_124 = RG_rl_185 ;
	7'h4e :
		TR_124 = RG_rl_185 ;
	7'h4f :
		TR_124 = RG_rl_185 ;
	7'h50 :
		TR_124 = RG_rl_185 ;
	7'h51 :
		TR_124 = RG_rl_185 ;
	7'h52 :
		TR_124 = RG_rl_185 ;
	7'h53 :
		TR_124 = RG_rl_185 ;
	7'h54 :
		TR_124 = RG_rl_185 ;
	7'h55 :
		TR_124 = RG_rl_185 ;
	7'h56 :
		TR_124 = RG_rl_185 ;
	7'h57 :
		TR_124 = RG_rl_185 ;
	7'h58 :
		TR_124 = RG_rl_185 ;
	7'h59 :
		TR_124 = RG_rl_185 ;
	7'h5a :
		TR_124 = RG_rl_185 ;
	7'h5b :
		TR_124 = RG_rl_185 ;
	7'h5c :
		TR_124 = RG_rl_185 ;
	7'h5d :
		TR_124 = RG_rl_185 ;
	7'h5e :
		TR_124 = RG_rl_185 ;
	7'h5f :
		TR_124 = RG_rl_185 ;
	7'h60 :
		TR_124 = RG_rl_185 ;
	7'h61 :
		TR_124 = RG_rl_185 ;
	7'h62 :
		TR_124 = RG_rl_185 ;
	7'h63 :
		TR_124 = RG_rl_185 ;
	7'h64 :
		TR_124 = RG_rl_185 ;
	7'h65 :
		TR_124 = RG_rl_185 ;
	7'h66 :
		TR_124 = RG_rl_185 ;
	7'h67 :
		TR_124 = RG_rl_185 ;
	7'h68 :
		TR_124 = RG_rl_185 ;
	7'h69 :
		TR_124 = RG_rl_185 ;
	7'h6a :
		TR_124 = RG_rl_185 ;
	7'h6b :
		TR_124 = RG_rl_185 ;
	7'h6c :
		TR_124 = RG_rl_185 ;
	7'h6d :
		TR_124 = RG_rl_185 ;
	7'h6e :
		TR_124 = RG_rl_185 ;
	7'h6f :
		TR_124 = RG_rl_185 ;
	7'h70 :
		TR_124 = 9'h000 ;	// line#=../rle.cpp:79
	7'h71 :
		TR_124 = RG_rl_185 ;
	7'h72 :
		TR_124 = RG_rl_185 ;
	7'h73 :
		TR_124 = RG_rl_185 ;
	7'h74 :
		TR_124 = RG_rl_185 ;
	7'h75 :
		TR_124 = RG_rl_185 ;
	7'h76 :
		TR_124 = RG_rl_185 ;
	7'h77 :
		TR_124 = RG_rl_185 ;
	7'h78 :
		TR_124 = RG_rl_185 ;
	7'h79 :
		TR_124 = RG_rl_185 ;
	7'h7a :
		TR_124 = RG_rl_185 ;
	7'h7b :
		TR_124 = RG_rl_185 ;
	7'h7c :
		TR_124 = RG_rl_185 ;
	7'h7d :
		TR_124 = RG_rl_185 ;
	7'h7e :
		TR_124 = RG_rl_185 ;
	7'h7f :
		TR_124 = RG_rl_185 ;
	default :
		TR_124 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_54 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h01 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h02 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h03 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h04 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h05 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h06 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h07 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h08 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h09 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h10 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h11 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h12 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h13 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h14 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h15 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h16 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h17 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h18 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h19 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h20 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h21 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h22 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h23 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h24 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h25 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h26 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h27 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h28 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h29 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h30 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h31 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h32 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h33 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h34 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h35 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h36 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h37 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h38 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h39 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h40 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h41 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h42 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h43 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h44 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h45 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h46 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h47 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h48 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h49 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h50 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h51 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h52 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h53 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h54 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h55 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h56 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h57 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h58 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h59 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h60 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h61 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h62 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h63 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h64 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h65 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h66 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h67 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h68 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h69 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h70 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h71 :
		TR_125 = 9'h000 ;	// line#=../rle.cpp:79
	7'h72 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h73 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h74 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h75 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h76 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h77 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h78 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h79 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7f :
		TR_125 = RG_quantized_block_rl_54 ;
	default :
		TR_125 = 9'hx ;
	endcase
always @ ( RG_rl_186 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_126 = RG_rl_186 ;
	7'h01 :
		TR_126 = RG_rl_186 ;
	7'h02 :
		TR_126 = RG_rl_186 ;
	7'h03 :
		TR_126 = RG_rl_186 ;
	7'h04 :
		TR_126 = RG_rl_186 ;
	7'h05 :
		TR_126 = RG_rl_186 ;
	7'h06 :
		TR_126 = RG_rl_186 ;
	7'h07 :
		TR_126 = RG_rl_186 ;
	7'h08 :
		TR_126 = RG_rl_186 ;
	7'h09 :
		TR_126 = RG_rl_186 ;
	7'h0a :
		TR_126 = RG_rl_186 ;
	7'h0b :
		TR_126 = RG_rl_186 ;
	7'h0c :
		TR_126 = RG_rl_186 ;
	7'h0d :
		TR_126 = RG_rl_186 ;
	7'h0e :
		TR_126 = RG_rl_186 ;
	7'h0f :
		TR_126 = RG_rl_186 ;
	7'h10 :
		TR_126 = RG_rl_186 ;
	7'h11 :
		TR_126 = RG_rl_186 ;
	7'h12 :
		TR_126 = RG_rl_186 ;
	7'h13 :
		TR_126 = RG_rl_186 ;
	7'h14 :
		TR_126 = RG_rl_186 ;
	7'h15 :
		TR_126 = RG_rl_186 ;
	7'h16 :
		TR_126 = RG_rl_186 ;
	7'h17 :
		TR_126 = RG_rl_186 ;
	7'h18 :
		TR_126 = RG_rl_186 ;
	7'h19 :
		TR_126 = RG_rl_186 ;
	7'h1a :
		TR_126 = RG_rl_186 ;
	7'h1b :
		TR_126 = RG_rl_186 ;
	7'h1c :
		TR_126 = RG_rl_186 ;
	7'h1d :
		TR_126 = RG_rl_186 ;
	7'h1e :
		TR_126 = RG_rl_186 ;
	7'h1f :
		TR_126 = RG_rl_186 ;
	7'h20 :
		TR_126 = RG_rl_186 ;
	7'h21 :
		TR_126 = RG_rl_186 ;
	7'h22 :
		TR_126 = RG_rl_186 ;
	7'h23 :
		TR_126 = RG_rl_186 ;
	7'h24 :
		TR_126 = RG_rl_186 ;
	7'h25 :
		TR_126 = RG_rl_186 ;
	7'h26 :
		TR_126 = RG_rl_186 ;
	7'h27 :
		TR_126 = RG_rl_186 ;
	7'h28 :
		TR_126 = RG_rl_186 ;
	7'h29 :
		TR_126 = RG_rl_186 ;
	7'h2a :
		TR_126 = RG_rl_186 ;
	7'h2b :
		TR_126 = RG_rl_186 ;
	7'h2c :
		TR_126 = RG_rl_186 ;
	7'h2d :
		TR_126 = RG_rl_186 ;
	7'h2e :
		TR_126 = RG_rl_186 ;
	7'h2f :
		TR_126 = RG_rl_186 ;
	7'h30 :
		TR_126 = RG_rl_186 ;
	7'h31 :
		TR_126 = RG_rl_186 ;
	7'h32 :
		TR_126 = RG_rl_186 ;
	7'h33 :
		TR_126 = RG_rl_186 ;
	7'h34 :
		TR_126 = RG_rl_186 ;
	7'h35 :
		TR_126 = RG_rl_186 ;
	7'h36 :
		TR_126 = RG_rl_186 ;
	7'h37 :
		TR_126 = RG_rl_186 ;
	7'h38 :
		TR_126 = RG_rl_186 ;
	7'h39 :
		TR_126 = RG_rl_186 ;
	7'h3a :
		TR_126 = RG_rl_186 ;
	7'h3b :
		TR_126 = RG_rl_186 ;
	7'h3c :
		TR_126 = RG_rl_186 ;
	7'h3d :
		TR_126 = RG_rl_186 ;
	7'h3e :
		TR_126 = RG_rl_186 ;
	7'h3f :
		TR_126 = RG_rl_186 ;
	7'h40 :
		TR_126 = RG_rl_186 ;
	7'h41 :
		TR_126 = RG_rl_186 ;
	7'h42 :
		TR_126 = RG_rl_186 ;
	7'h43 :
		TR_126 = RG_rl_186 ;
	7'h44 :
		TR_126 = RG_rl_186 ;
	7'h45 :
		TR_126 = RG_rl_186 ;
	7'h46 :
		TR_126 = RG_rl_186 ;
	7'h47 :
		TR_126 = RG_rl_186 ;
	7'h48 :
		TR_126 = RG_rl_186 ;
	7'h49 :
		TR_126 = RG_rl_186 ;
	7'h4a :
		TR_126 = RG_rl_186 ;
	7'h4b :
		TR_126 = RG_rl_186 ;
	7'h4c :
		TR_126 = RG_rl_186 ;
	7'h4d :
		TR_126 = RG_rl_186 ;
	7'h4e :
		TR_126 = RG_rl_186 ;
	7'h4f :
		TR_126 = RG_rl_186 ;
	7'h50 :
		TR_126 = RG_rl_186 ;
	7'h51 :
		TR_126 = RG_rl_186 ;
	7'h52 :
		TR_126 = RG_rl_186 ;
	7'h53 :
		TR_126 = RG_rl_186 ;
	7'h54 :
		TR_126 = RG_rl_186 ;
	7'h55 :
		TR_126 = RG_rl_186 ;
	7'h56 :
		TR_126 = RG_rl_186 ;
	7'h57 :
		TR_126 = RG_rl_186 ;
	7'h58 :
		TR_126 = RG_rl_186 ;
	7'h59 :
		TR_126 = RG_rl_186 ;
	7'h5a :
		TR_126 = RG_rl_186 ;
	7'h5b :
		TR_126 = RG_rl_186 ;
	7'h5c :
		TR_126 = RG_rl_186 ;
	7'h5d :
		TR_126 = RG_rl_186 ;
	7'h5e :
		TR_126 = RG_rl_186 ;
	7'h5f :
		TR_126 = RG_rl_186 ;
	7'h60 :
		TR_126 = RG_rl_186 ;
	7'h61 :
		TR_126 = RG_rl_186 ;
	7'h62 :
		TR_126 = RG_rl_186 ;
	7'h63 :
		TR_126 = RG_rl_186 ;
	7'h64 :
		TR_126 = RG_rl_186 ;
	7'h65 :
		TR_126 = RG_rl_186 ;
	7'h66 :
		TR_126 = RG_rl_186 ;
	7'h67 :
		TR_126 = RG_rl_186 ;
	7'h68 :
		TR_126 = RG_rl_186 ;
	7'h69 :
		TR_126 = RG_rl_186 ;
	7'h6a :
		TR_126 = RG_rl_186 ;
	7'h6b :
		TR_126 = RG_rl_186 ;
	7'h6c :
		TR_126 = RG_rl_186 ;
	7'h6d :
		TR_126 = RG_rl_186 ;
	7'h6e :
		TR_126 = RG_rl_186 ;
	7'h6f :
		TR_126 = RG_rl_186 ;
	7'h70 :
		TR_126 = RG_rl_186 ;
	7'h71 :
		TR_126 = RG_rl_186 ;
	7'h72 :
		TR_126 = 9'h000 ;	// line#=../rle.cpp:79
	7'h73 :
		TR_126 = RG_rl_186 ;
	7'h74 :
		TR_126 = RG_rl_186 ;
	7'h75 :
		TR_126 = RG_rl_186 ;
	7'h76 :
		TR_126 = RG_rl_186 ;
	7'h77 :
		TR_126 = RG_rl_186 ;
	7'h78 :
		TR_126 = RG_rl_186 ;
	7'h79 :
		TR_126 = RG_rl_186 ;
	7'h7a :
		TR_126 = RG_rl_186 ;
	7'h7b :
		TR_126 = RG_rl_186 ;
	7'h7c :
		TR_126 = RG_rl_186 ;
	7'h7d :
		TR_126 = RG_rl_186 ;
	7'h7e :
		TR_126 = RG_rl_186 ;
	7'h7f :
		TR_126 = RG_rl_186 ;
	default :
		TR_126 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_55 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h01 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h02 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h03 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h04 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h05 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h06 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h07 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h08 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h09 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h0a :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h0b :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h0c :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h0d :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h0e :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h0f :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h10 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h11 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h12 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h13 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h14 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h15 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h16 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h17 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h18 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h19 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h1a :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h1b :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h1c :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h1d :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h1e :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h1f :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h20 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h21 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h22 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h23 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h24 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h25 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h26 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h27 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h28 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h29 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h2a :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h2b :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h2c :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h2d :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h2e :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h2f :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h30 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h31 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h32 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h33 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h34 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h35 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h36 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h37 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h38 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h39 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h3a :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h3b :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h3c :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h3d :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h3e :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h3f :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h40 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h41 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h42 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h43 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h44 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h45 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h46 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h47 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h48 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h49 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h4a :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h4b :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h4c :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h4d :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h4e :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h4f :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h50 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h51 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h52 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h53 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h54 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h55 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h56 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h57 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h58 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h59 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h5a :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h5b :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h5c :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h5d :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h5e :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h5f :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h60 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h61 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h62 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h63 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h64 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h65 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h66 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h67 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h68 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h69 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h6a :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h6b :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h6c :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h6d :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h6e :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h6f :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h70 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h71 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h72 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h73 :
		TR_127 = 9'h000 ;	// line#=../rle.cpp:79
	7'h74 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h75 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h76 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h77 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h78 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h79 :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h7a :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h7b :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h7c :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h7d :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h7e :
		TR_127 = RG_quantized_block_rl_55 ;
	7'h7f :
		TR_127 = RG_quantized_block_rl_55 ;
	default :
		TR_127 = 9'hx ;
	endcase
always @ ( RG_rl_187 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_128 = RG_rl_187 ;
	7'h01 :
		TR_128 = RG_rl_187 ;
	7'h02 :
		TR_128 = RG_rl_187 ;
	7'h03 :
		TR_128 = RG_rl_187 ;
	7'h04 :
		TR_128 = RG_rl_187 ;
	7'h05 :
		TR_128 = RG_rl_187 ;
	7'h06 :
		TR_128 = RG_rl_187 ;
	7'h07 :
		TR_128 = RG_rl_187 ;
	7'h08 :
		TR_128 = RG_rl_187 ;
	7'h09 :
		TR_128 = RG_rl_187 ;
	7'h0a :
		TR_128 = RG_rl_187 ;
	7'h0b :
		TR_128 = RG_rl_187 ;
	7'h0c :
		TR_128 = RG_rl_187 ;
	7'h0d :
		TR_128 = RG_rl_187 ;
	7'h0e :
		TR_128 = RG_rl_187 ;
	7'h0f :
		TR_128 = RG_rl_187 ;
	7'h10 :
		TR_128 = RG_rl_187 ;
	7'h11 :
		TR_128 = RG_rl_187 ;
	7'h12 :
		TR_128 = RG_rl_187 ;
	7'h13 :
		TR_128 = RG_rl_187 ;
	7'h14 :
		TR_128 = RG_rl_187 ;
	7'h15 :
		TR_128 = RG_rl_187 ;
	7'h16 :
		TR_128 = RG_rl_187 ;
	7'h17 :
		TR_128 = RG_rl_187 ;
	7'h18 :
		TR_128 = RG_rl_187 ;
	7'h19 :
		TR_128 = RG_rl_187 ;
	7'h1a :
		TR_128 = RG_rl_187 ;
	7'h1b :
		TR_128 = RG_rl_187 ;
	7'h1c :
		TR_128 = RG_rl_187 ;
	7'h1d :
		TR_128 = RG_rl_187 ;
	7'h1e :
		TR_128 = RG_rl_187 ;
	7'h1f :
		TR_128 = RG_rl_187 ;
	7'h20 :
		TR_128 = RG_rl_187 ;
	7'h21 :
		TR_128 = RG_rl_187 ;
	7'h22 :
		TR_128 = RG_rl_187 ;
	7'h23 :
		TR_128 = RG_rl_187 ;
	7'h24 :
		TR_128 = RG_rl_187 ;
	7'h25 :
		TR_128 = RG_rl_187 ;
	7'h26 :
		TR_128 = RG_rl_187 ;
	7'h27 :
		TR_128 = RG_rl_187 ;
	7'h28 :
		TR_128 = RG_rl_187 ;
	7'h29 :
		TR_128 = RG_rl_187 ;
	7'h2a :
		TR_128 = RG_rl_187 ;
	7'h2b :
		TR_128 = RG_rl_187 ;
	7'h2c :
		TR_128 = RG_rl_187 ;
	7'h2d :
		TR_128 = RG_rl_187 ;
	7'h2e :
		TR_128 = RG_rl_187 ;
	7'h2f :
		TR_128 = RG_rl_187 ;
	7'h30 :
		TR_128 = RG_rl_187 ;
	7'h31 :
		TR_128 = RG_rl_187 ;
	7'h32 :
		TR_128 = RG_rl_187 ;
	7'h33 :
		TR_128 = RG_rl_187 ;
	7'h34 :
		TR_128 = RG_rl_187 ;
	7'h35 :
		TR_128 = RG_rl_187 ;
	7'h36 :
		TR_128 = RG_rl_187 ;
	7'h37 :
		TR_128 = RG_rl_187 ;
	7'h38 :
		TR_128 = RG_rl_187 ;
	7'h39 :
		TR_128 = RG_rl_187 ;
	7'h3a :
		TR_128 = RG_rl_187 ;
	7'h3b :
		TR_128 = RG_rl_187 ;
	7'h3c :
		TR_128 = RG_rl_187 ;
	7'h3d :
		TR_128 = RG_rl_187 ;
	7'h3e :
		TR_128 = RG_rl_187 ;
	7'h3f :
		TR_128 = RG_rl_187 ;
	7'h40 :
		TR_128 = RG_rl_187 ;
	7'h41 :
		TR_128 = RG_rl_187 ;
	7'h42 :
		TR_128 = RG_rl_187 ;
	7'h43 :
		TR_128 = RG_rl_187 ;
	7'h44 :
		TR_128 = RG_rl_187 ;
	7'h45 :
		TR_128 = RG_rl_187 ;
	7'h46 :
		TR_128 = RG_rl_187 ;
	7'h47 :
		TR_128 = RG_rl_187 ;
	7'h48 :
		TR_128 = RG_rl_187 ;
	7'h49 :
		TR_128 = RG_rl_187 ;
	7'h4a :
		TR_128 = RG_rl_187 ;
	7'h4b :
		TR_128 = RG_rl_187 ;
	7'h4c :
		TR_128 = RG_rl_187 ;
	7'h4d :
		TR_128 = RG_rl_187 ;
	7'h4e :
		TR_128 = RG_rl_187 ;
	7'h4f :
		TR_128 = RG_rl_187 ;
	7'h50 :
		TR_128 = RG_rl_187 ;
	7'h51 :
		TR_128 = RG_rl_187 ;
	7'h52 :
		TR_128 = RG_rl_187 ;
	7'h53 :
		TR_128 = RG_rl_187 ;
	7'h54 :
		TR_128 = RG_rl_187 ;
	7'h55 :
		TR_128 = RG_rl_187 ;
	7'h56 :
		TR_128 = RG_rl_187 ;
	7'h57 :
		TR_128 = RG_rl_187 ;
	7'h58 :
		TR_128 = RG_rl_187 ;
	7'h59 :
		TR_128 = RG_rl_187 ;
	7'h5a :
		TR_128 = RG_rl_187 ;
	7'h5b :
		TR_128 = RG_rl_187 ;
	7'h5c :
		TR_128 = RG_rl_187 ;
	7'h5d :
		TR_128 = RG_rl_187 ;
	7'h5e :
		TR_128 = RG_rl_187 ;
	7'h5f :
		TR_128 = RG_rl_187 ;
	7'h60 :
		TR_128 = RG_rl_187 ;
	7'h61 :
		TR_128 = RG_rl_187 ;
	7'h62 :
		TR_128 = RG_rl_187 ;
	7'h63 :
		TR_128 = RG_rl_187 ;
	7'h64 :
		TR_128 = RG_rl_187 ;
	7'h65 :
		TR_128 = RG_rl_187 ;
	7'h66 :
		TR_128 = RG_rl_187 ;
	7'h67 :
		TR_128 = RG_rl_187 ;
	7'h68 :
		TR_128 = RG_rl_187 ;
	7'h69 :
		TR_128 = RG_rl_187 ;
	7'h6a :
		TR_128 = RG_rl_187 ;
	7'h6b :
		TR_128 = RG_rl_187 ;
	7'h6c :
		TR_128 = RG_rl_187 ;
	7'h6d :
		TR_128 = RG_rl_187 ;
	7'h6e :
		TR_128 = RG_rl_187 ;
	7'h6f :
		TR_128 = RG_rl_187 ;
	7'h70 :
		TR_128 = RG_rl_187 ;
	7'h71 :
		TR_128 = RG_rl_187 ;
	7'h72 :
		TR_128 = RG_rl_187 ;
	7'h73 :
		TR_128 = RG_rl_187 ;
	7'h74 :
		TR_128 = 9'h000 ;	// line#=../rle.cpp:79
	7'h75 :
		TR_128 = RG_rl_187 ;
	7'h76 :
		TR_128 = RG_rl_187 ;
	7'h77 :
		TR_128 = RG_rl_187 ;
	7'h78 :
		TR_128 = RG_rl_187 ;
	7'h79 :
		TR_128 = RG_rl_187 ;
	7'h7a :
		TR_128 = RG_rl_187 ;
	7'h7b :
		TR_128 = RG_rl_187 ;
	7'h7c :
		TR_128 = RG_rl_187 ;
	7'h7d :
		TR_128 = RG_rl_187 ;
	7'h7e :
		TR_128 = RG_rl_187 ;
	7'h7f :
		TR_128 = RG_rl_187 ;
	default :
		TR_128 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_56 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h01 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h02 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h03 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h04 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h05 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h06 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h07 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h08 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h09 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h0a :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h0b :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h0c :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h0d :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h0e :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h0f :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h10 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h11 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h12 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h13 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h14 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h15 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h16 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h17 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h18 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h19 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h1a :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h1b :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h1c :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h1d :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h1e :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h1f :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h20 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h21 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h22 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h23 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h24 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h25 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h26 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h27 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h28 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h29 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h2a :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h2b :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h2c :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h2d :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h2e :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h2f :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h30 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h31 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h32 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h33 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h34 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h35 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h36 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h37 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h38 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h39 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h3a :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h3b :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h3c :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h3d :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h3e :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h3f :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h40 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h41 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h42 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h43 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h44 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h45 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h46 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h47 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h48 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h49 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h4a :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h4b :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h4c :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h4d :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h4e :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h4f :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h50 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h51 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h52 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h53 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h54 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h55 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h56 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h57 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h58 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h59 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h5a :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h5b :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h5c :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h5d :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h5e :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h5f :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h60 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h61 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h62 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h63 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h64 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h65 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h66 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h67 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h68 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h69 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h6a :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h6b :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h6c :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h6d :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h6e :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h6f :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h70 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h71 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h72 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h73 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h74 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h75 :
		TR_129 = 9'h000 ;	// line#=../rle.cpp:79
	7'h76 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h77 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h78 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h79 :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h7a :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h7b :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h7c :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h7d :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h7e :
		TR_129 = RG_quantized_block_rl_56 ;
	7'h7f :
		TR_129 = RG_quantized_block_rl_56 ;
	default :
		TR_129 = 9'hx ;
	endcase
always @ ( RG_rl_188 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_130 = RG_rl_188 ;
	7'h01 :
		TR_130 = RG_rl_188 ;
	7'h02 :
		TR_130 = RG_rl_188 ;
	7'h03 :
		TR_130 = RG_rl_188 ;
	7'h04 :
		TR_130 = RG_rl_188 ;
	7'h05 :
		TR_130 = RG_rl_188 ;
	7'h06 :
		TR_130 = RG_rl_188 ;
	7'h07 :
		TR_130 = RG_rl_188 ;
	7'h08 :
		TR_130 = RG_rl_188 ;
	7'h09 :
		TR_130 = RG_rl_188 ;
	7'h0a :
		TR_130 = RG_rl_188 ;
	7'h0b :
		TR_130 = RG_rl_188 ;
	7'h0c :
		TR_130 = RG_rl_188 ;
	7'h0d :
		TR_130 = RG_rl_188 ;
	7'h0e :
		TR_130 = RG_rl_188 ;
	7'h0f :
		TR_130 = RG_rl_188 ;
	7'h10 :
		TR_130 = RG_rl_188 ;
	7'h11 :
		TR_130 = RG_rl_188 ;
	7'h12 :
		TR_130 = RG_rl_188 ;
	7'h13 :
		TR_130 = RG_rl_188 ;
	7'h14 :
		TR_130 = RG_rl_188 ;
	7'h15 :
		TR_130 = RG_rl_188 ;
	7'h16 :
		TR_130 = RG_rl_188 ;
	7'h17 :
		TR_130 = RG_rl_188 ;
	7'h18 :
		TR_130 = RG_rl_188 ;
	7'h19 :
		TR_130 = RG_rl_188 ;
	7'h1a :
		TR_130 = RG_rl_188 ;
	7'h1b :
		TR_130 = RG_rl_188 ;
	7'h1c :
		TR_130 = RG_rl_188 ;
	7'h1d :
		TR_130 = RG_rl_188 ;
	7'h1e :
		TR_130 = RG_rl_188 ;
	7'h1f :
		TR_130 = RG_rl_188 ;
	7'h20 :
		TR_130 = RG_rl_188 ;
	7'h21 :
		TR_130 = RG_rl_188 ;
	7'h22 :
		TR_130 = RG_rl_188 ;
	7'h23 :
		TR_130 = RG_rl_188 ;
	7'h24 :
		TR_130 = RG_rl_188 ;
	7'h25 :
		TR_130 = RG_rl_188 ;
	7'h26 :
		TR_130 = RG_rl_188 ;
	7'h27 :
		TR_130 = RG_rl_188 ;
	7'h28 :
		TR_130 = RG_rl_188 ;
	7'h29 :
		TR_130 = RG_rl_188 ;
	7'h2a :
		TR_130 = RG_rl_188 ;
	7'h2b :
		TR_130 = RG_rl_188 ;
	7'h2c :
		TR_130 = RG_rl_188 ;
	7'h2d :
		TR_130 = RG_rl_188 ;
	7'h2e :
		TR_130 = RG_rl_188 ;
	7'h2f :
		TR_130 = RG_rl_188 ;
	7'h30 :
		TR_130 = RG_rl_188 ;
	7'h31 :
		TR_130 = RG_rl_188 ;
	7'h32 :
		TR_130 = RG_rl_188 ;
	7'h33 :
		TR_130 = RG_rl_188 ;
	7'h34 :
		TR_130 = RG_rl_188 ;
	7'h35 :
		TR_130 = RG_rl_188 ;
	7'h36 :
		TR_130 = RG_rl_188 ;
	7'h37 :
		TR_130 = RG_rl_188 ;
	7'h38 :
		TR_130 = RG_rl_188 ;
	7'h39 :
		TR_130 = RG_rl_188 ;
	7'h3a :
		TR_130 = RG_rl_188 ;
	7'h3b :
		TR_130 = RG_rl_188 ;
	7'h3c :
		TR_130 = RG_rl_188 ;
	7'h3d :
		TR_130 = RG_rl_188 ;
	7'h3e :
		TR_130 = RG_rl_188 ;
	7'h3f :
		TR_130 = RG_rl_188 ;
	7'h40 :
		TR_130 = RG_rl_188 ;
	7'h41 :
		TR_130 = RG_rl_188 ;
	7'h42 :
		TR_130 = RG_rl_188 ;
	7'h43 :
		TR_130 = RG_rl_188 ;
	7'h44 :
		TR_130 = RG_rl_188 ;
	7'h45 :
		TR_130 = RG_rl_188 ;
	7'h46 :
		TR_130 = RG_rl_188 ;
	7'h47 :
		TR_130 = RG_rl_188 ;
	7'h48 :
		TR_130 = RG_rl_188 ;
	7'h49 :
		TR_130 = RG_rl_188 ;
	7'h4a :
		TR_130 = RG_rl_188 ;
	7'h4b :
		TR_130 = RG_rl_188 ;
	7'h4c :
		TR_130 = RG_rl_188 ;
	7'h4d :
		TR_130 = RG_rl_188 ;
	7'h4e :
		TR_130 = RG_rl_188 ;
	7'h4f :
		TR_130 = RG_rl_188 ;
	7'h50 :
		TR_130 = RG_rl_188 ;
	7'h51 :
		TR_130 = RG_rl_188 ;
	7'h52 :
		TR_130 = RG_rl_188 ;
	7'h53 :
		TR_130 = RG_rl_188 ;
	7'h54 :
		TR_130 = RG_rl_188 ;
	7'h55 :
		TR_130 = RG_rl_188 ;
	7'h56 :
		TR_130 = RG_rl_188 ;
	7'h57 :
		TR_130 = RG_rl_188 ;
	7'h58 :
		TR_130 = RG_rl_188 ;
	7'h59 :
		TR_130 = RG_rl_188 ;
	7'h5a :
		TR_130 = RG_rl_188 ;
	7'h5b :
		TR_130 = RG_rl_188 ;
	7'h5c :
		TR_130 = RG_rl_188 ;
	7'h5d :
		TR_130 = RG_rl_188 ;
	7'h5e :
		TR_130 = RG_rl_188 ;
	7'h5f :
		TR_130 = RG_rl_188 ;
	7'h60 :
		TR_130 = RG_rl_188 ;
	7'h61 :
		TR_130 = RG_rl_188 ;
	7'h62 :
		TR_130 = RG_rl_188 ;
	7'h63 :
		TR_130 = RG_rl_188 ;
	7'h64 :
		TR_130 = RG_rl_188 ;
	7'h65 :
		TR_130 = RG_rl_188 ;
	7'h66 :
		TR_130 = RG_rl_188 ;
	7'h67 :
		TR_130 = RG_rl_188 ;
	7'h68 :
		TR_130 = RG_rl_188 ;
	7'h69 :
		TR_130 = RG_rl_188 ;
	7'h6a :
		TR_130 = RG_rl_188 ;
	7'h6b :
		TR_130 = RG_rl_188 ;
	7'h6c :
		TR_130 = RG_rl_188 ;
	7'h6d :
		TR_130 = RG_rl_188 ;
	7'h6e :
		TR_130 = RG_rl_188 ;
	7'h6f :
		TR_130 = RG_rl_188 ;
	7'h70 :
		TR_130 = RG_rl_188 ;
	7'h71 :
		TR_130 = RG_rl_188 ;
	7'h72 :
		TR_130 = RG_rl_188 ;
	7'h73 :
		TR_130 = RG_rl_188 ;
	7'h74 :
		TR_130 = RG_rl_188 ;
	7'h75 :
		TR_130 = RG_rl_188 ;
	7'h76 :
		TR_130 = 9'h000 ;	// line#=../rle.cpp:79
	7'h77 :
		TR_130 = RG_rl_188 ;
	7'h78 :
		TR_130 = RG_rl_188 ;
	7'h79 :
		TR_130 = RG_rl_188 ;
	7'h7a :
		TR_130 = RG_rl_188 ;
	7'h7b :
		TR_130 = RG_rl_188 ;
	7'h7c :
		TR_130 = RG_rl_188 ;
	7'h7d :
		TR_130 = RG_rl_188 ;
	7'h7e :
		TR_130 = RG_rl_188 ;
	7'h7f :
		TR_130 = RG_rl_188 ;
	default :
		TR_130 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_57 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h01 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h02 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h03 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h04 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h05 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h06 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h07 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h08 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h09 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h0a :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h0b :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h0c :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h0d :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h0e :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h0f :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h10 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h11 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h12 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h13 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h14 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h15 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h16 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h17 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h18 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h19 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h1a :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h1b :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h1c :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h1d :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h1e :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h1f :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h20 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h21 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h22 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h23 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h24 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h25 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h26 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h27 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h28 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h29 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h2a :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h2b :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h2c :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h2d :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h2e :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h2f :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h30 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h31 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h32 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h33 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h34 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h35 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h36 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h37 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h38 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h39 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h3a :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h3b :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h3c :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h3d :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h3e :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h3f :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h40 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h41 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h42 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h43 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h44 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h45 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h46 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h47 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h48 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h49 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h4a :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h4b :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h4c :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h4d :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h4e :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h4f :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h50 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h51 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h52 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h53 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h54 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h55 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h56 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h57 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h58 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h59 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h5a :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h5b :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h5c :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h5d :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h5e :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h5f :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h60 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h61 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h62 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h63 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h64 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h65 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h66 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h67 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h68 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h69 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h6a :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h6b :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h6c :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h6d :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h6e :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h6f :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h70 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h71 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h72 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h73 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h74 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h75 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h76 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h77 :
		TR_131 = 9'h000 ;	// line#=../rle.cpp:79
	7'h78 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h79 :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h7a :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h7b :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h7c :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h7d :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h7e :
		TR_131 = RG_quantized_block_rl_57 ;
	7'h7f :
		TR_131 = RG_quantized_block_rl_57 ;
	default :
		TR_131 = 9'hx ;
	endcase
always @ ( RG_rl_189 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_132 = RG_rl_189 ;
	7'h01 :
		TR_132 = RG_rl_189 ;
	7'h02 :
		TR_132 = RG_rl_189 ;
	7'h03 :
		TR_132 = RG_rl_189 ;
	7'h04 :
		TR_132 = RG_rl_189 ;
	7'h05 :
		TR_132 = RG_rl_189 ;
	7'h06 :
		TR_132 = RG_rl_189 ;
	7'h07 :
		TR_132 = RG_rl_189 ;
	7'h08 :
		TR_132 = RG_rl_189 ;
	7'h09 :
		TR_132 = RG_rl_189 ;
	7'h0a :
		TR_132 = RG_rl_189 ;
	7'h0b :
		TR_132 = RG_rl_189 ;
	7'h0c :
		TR_132 = RG_rl_189 ;
	7'h0d :
		TR_132 = RG_rl_189 ;
	7'h0e :
		TR_132 = RG_rl_189 ;
	7'h0f :
		TR_132 = RG_rl_189 ;
	7'h10 :
		TR_132 = RG_rl_189 ;
	7'h11 :
		TR_132 = RG_rl_189 ;
	7'h12 :
		TR_132 = RG_rl_189 ;
	7'h13 :
		TR_132 = RG_rl_189 ;
	7'h14 :
		TR_132 = RG_rl_189 ;
	7'h15 :
		TR_132 = RG_rl_189 ;
	7'h16 :
		TR_132 = RG_rl_189 ;
	7'h17 :
		TR_132 = RG_rl_189 ;
	7'h18 :
		TR_132 = RG_rl_189 ;
	7'h19 :
		TR_132 = RG_rl_189 ;
	7'h1a :
		TR_132 = RG_rl_189 ;
	7'h1b :
		TR_132 = RG_rl_189 ;
	7'h1c :
		TR_132 = RG_rl_189 ;
	7'h1d :
		TR_132 = RG_rl_189 ;
	7'h1e :
		TR_132 = RG_rl_189 ;
	7'h1f :
		TR_132 = RG_rl_189 ;
	7'h20 :
		TR_132 = RG_rl_189 ;
	7'h21 :
		TR_132 = RG_rl_189 ;
	7'h22 :
		TR_132 = RG_rl_189 ;
	7'h23 :
		TR_132 = RG_rl_189 ;
	7'h24 :
		TR_132 = RG_rl_189 ;
	7'h25 :
		TR_132 = RG_rl_189 ;
	7'h26 :
		TR_132 = RG_rl_189 ;
	7'h27 :
		TR_132 = RG_rl_189 ;
	7'h28 :
		TR_132 = RG_rl_189 ;
	7'h29 :
		TR_132 = RG_rl_189 ;
	7'h2a :
		TR_132 = RG_rl_189 ;
	7'h2b :
		TR_132 = RG_rl_189 ;
	7'h2c :
		TR_132 = RG_rl_189 ;
	7'h2d :
		TR_132 = RG_rl_189 ;
	7'h2e :
		TR_132 = RG_rl_189 ;
	7'h2f :
		TR_132 = RG_rl_189 ;
	7'h30 :
		TR_132 = RG_rl_189 ;
	7'h31 :
		TR_132 = RG_rl_189 ;
	7'h32 :
		TR_132 = RG_rl_189 ;
	7'h33 :
		TR_132 = RG_rl_189 ;
	7'h34 :
		TR_132 = RG_rl_189 ;
	7'h35 :
		TR_132 = RG_rl_189 ;
	7'h36 :
		TR_132 = RG_rl_189 ;
	7'h37 :
		TR_132 = RG_rl_189 ;
	7'h38 :
		TR_132 = RG_rl_189 ;
	7'h39 :
		TR_132 = RG_rl_189 ;
	7'h3a :
		TR_132 = RG_rl_189 ;
	7'h3b :
		TR_132 = RG_rl_189 ;
	7'h3c :
		TR_132 = RG_rl_189 ;
	7'h3d :
		TR_132 = RG_rl_189 ;
	7'h3e :
		TR_132 = RG_rl_189 ;
	7'h3f :
		TR_132 = RG_rl_189 ;
	7'h40 :
		TR_132 = RG_rl_189 ;
	7'h41 :
		TR_132 = RG_rl_189 ;
	7'h42 :
		TR_132 = RG_rl_189 ;
	7'h43 :
		TR_132 = RG_rl_189 ;
	7'h44 :
		TR_132 = RG_rl_189 ;
	7'h45 :
		TR_132 = RG_rl_189 ;
	7'h46 :
		TR_132 = RG_rl_189 ;
	7'h47 :
		TR_132 = RG_rl_189 ;
	7'h48 :
		TR_132 = RG_rl_189 ;
	7'h49 :
		TR_132 = RG_rl_189 ;
	7'h4a :
		TR_132 = RG_rl_189 ;
	7'h4b :
		TR_132 = RG_rl_189 ;
	7'h4c :
		TR_132 = RG_rl_189 ;
	7'h4d :
		TR_132 = RG_rl_189 ;
	7'h4e :
		TR_132 = RG_rl_189 ;
	7'h4f :
		TR_132 = RG_rl_189 ;
	7'h50 :
		TR_132 = RG_rl_189 ;
	7'h51 :
		TR_132 = RG_rl_189 ;
	7'h52 :
		TR_132 = RG_rl_189 ;
	7'h53 :
		TR_132 = RG_rl_189 ;
	7'h54 :
		TR_132 = RG_rl_189 ;
	7'h55 :
		TR_132 = RG_rl_189 ;
	7'h56 :
		TR_132 = RG_rl_189 ;
	7'h57 :
		TR_132 = RG_rl_189 ;
	7'h58 :
		TR_132 = RG_rl_189 ;
	7'h59 :
		TR_132 = RG_rl_189 ;
	7'h5a :
		TR_132 = RG_rl_189 ;
	7'h5b :
		TR_132 = RG_rl_189 ;
	7'h5c :
		TR_132 = RG_rl_189 ;
	7'h5d :
		TR_132 = RG_rl_189 ;
	7'h5e :
		TR_132 = RG_rl_189 ;
	7'h5f :
		TR_132 = RG_rl_189 ;
	7'h60 :
		TR_132 = RG_rl_189 ;
	7'h61 :
		TR_132 = RG_rl_189 ;
	7'h62 :
		TR_132 = RG_rl_189 ;
	7'h63 :
		TR_132 = RG_rl_189 ;
	7'h64 :
		TR_132 = RG_rl_189 ;
	7'h65 :
		TR_132 = RG_rl_189 ;
	7'h66 :
		TR_132 = RG_rl_189 ;
	7'h67 :
		TR_132 = RG_rl_189 ;
	7'h68 :
		TR_132 = RG_rl_189 ;
	7'h69 :
		TR_132 = RG_rl_189 ;
	7'h6a :
		TR_132 = RG_rl_189 ;
	7'h6b :
		TR_132 = RG_rl_189 ;
	7'h6c :
		TR_132 = RG_rl_189 ;
	7'h6d :
		TR_132 = RG_rl_189 ;
	7'h6e :
		TR_132 = RG_rl_189 ;
	7'h6f :
		TR_132 = RG_rl_189 ;
	7'h70 :
		TR_132 = RG_rl_189 ;
	7'h71 :
		TR_132 = RG_rl_189 ;
	7'h72 :
		TR_132 = RG_rl_189 ;
	7'h73 :
		TR_132 = RG_rl_189 ;
	7'h74 :
		TR_132 = RG_rl_189 ;
	7'h75 :
		TR_132 = RG_rl_189 ;
	7'h76 :
		TR_132 = RG_rl_189 ;
	7'h77 :
		TR_132 = RG_rl_189 ;
	7'h78 :
		TR_132 = 9'h000 ;	// line#=../rle.cpp:79
	7'h79 :
		TR_132 = RG_rl_189 ;
	7'h7a :
		TR_132 = RG_rl_189 ;
	7'h7b :
		TR_132 = RG_rl_189 ;
	7'h7c :
		TR_132 = RG_rl_189 ;
	7'h7d :
		TR_132 = RG_rl_189 ;
	7'h7e :
		TR_132 = RG_rl_189 ;
	7'h7f :
		TR_132 = RG_rl_189 ;
	default :
		TR_132 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_58 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h01 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h02 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h03 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h04 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h05 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h06 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h07 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h08 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h09 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h0a :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h0b :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h0c :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h0d :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h0e :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h0f :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h10 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h11 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h12 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h13 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h14 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h15 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h16 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h17 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h18 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h19 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h1a :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h1b :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h1c :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h1d :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h1e :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h1f :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h20 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h21 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h22 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h23 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h24 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h25 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h26 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h27 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h28 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h29 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h2a :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h2b :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h2c :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h2d :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h2e :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h2f :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h30 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h31 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h32 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h33 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h34 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h35 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h36 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h37 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h38 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h39 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h3a :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h3b :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h3c :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h3d :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h3e :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h3f :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h40 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h41 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h42 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h43 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h44 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h45 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h46 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h47 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h48 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h49 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h4a :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h4b :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h4c :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h4d :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h4e :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h4f :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h50 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h51 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h52 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h53 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h54 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h55 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h56 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h57 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h58 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h59 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h5a :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h5b :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h5c :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h5d :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h5e :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h5f :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h60 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h61 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h62 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h63 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h64 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h65 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h66 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h67 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h68 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h69 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h6a :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h6b :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h6c :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h6d :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h6e :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h6f :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h70 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h71 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h72 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h73 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h74 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h75 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h76 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h77 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h78 :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h79 :
		TR_133 = 9'h000 ;	// line#=../rle.cpp:79
	7'h7a :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h7b :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h7c :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h7d :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h7e :
		TR_133 = RG_quantized_block_rl_58 ;
	7'h7f :
		TR_133 = RG_quantized_block_rl_58 ;
	default :
		TR_133 = 9'hx ;
	endcase
always @ ( RG_rl_190 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_134 = RG_rl_190 ;
	7'h01 :
		TR_134 = RG_rl_190 ;
	7'h02 :
		TR_134 = RG_rl_190 ;
	7'h03 :
		TR_134 = RG_rl_190 ;
	7'h04 :
		TR_134 = RG_rl_190 ;
	7'h05 :
		TR_134 = RG_rl_190 ;
	7'h06 :
		TR_134 = RG_rl_190 ;
	7'h07 :
		TR_134 = RG_rl_190 ;
	7'h08 :
		TR_134 = RG_rl_190 ;
	7'h09 :
		TR_134 = RG_rl_190 ;
	7'h0a :
		TR_134 = RG_rl_190 ;
	7'h0b :
		TR_134 = RG_rl_190 ;
	7'h0c :
		TR_134 = RG_rl_190 ;
	7'h0d :
		TR_134 = RG_rl_190 ;
	7'h0e :
		TR_134 = RG_rl_190 ;
	7'h0f :
		TR_134 = RG_rl_190 ;
	7'h10 :
		TR_134 = RG_rl_190 ;
	7'h11 :
		TR_134 = RG_rl_190 ;
	7'h12 :
		TR_134 = RG_rl_190 ;
	7'h13 :
		TR_134 = RG_rl_190 ;
	7'h14 :
		TR_134 = RG_rl_190 ;
	7'h15 :
		TR_134 = RG_rl_190 ;
	7'h16 :
		TR_134 = RG_rl_190 ;
	7'h17 :
		TR_134 = RG_rl_190 ;
	7'h18 :
		TR_134 = RG_rl_190 ;
	7'h19 :
		TR_134 = RG_rl_190 ;
	7'h1a :
		TR_134 = RG_rl_190 ;
	7'h1b :
		TR_134 = RG_rl_190 ;
	7'h1c :
		TR_134 = RG_rl_190 ;
	7'h1d :
		TR_134 = RG_rl_190 ;
	7'h1e :
		TR_134 = RG_rl_190 ;
	7'h1f :
		TR_134 = RG_rl_190 ;
	7'h20 :
		TR_134 = RG_rl_190 ;
	7'h21 :
		TR_134 = RG_rl_190 ;
	7'h22 :
		TR_134 = RG_rl_190 ;
	7'h23 :
		TR_134 = RG_rl_190 ;
	7'h24 :
		TR_134 = RG_rl_190 ;
	7'h25 :
		TR_134 = RG_rl_190 ;
	7'h26 :
		TR_134 = RG_rl_190 ;
	7'h27 :
		TR_134 = RG_rl_190 ;
	7'h28 :
		TR_134 = RG_rl_190 ;
	7'h29 :
		TR_134 = RG_rl_190 ;
	7'h2a :
		TR_134 = RG_rl_190 ;
	7'h2b :
		TR_134 = RG_rl_190 ;
	7'h2c :
		TR_134 = RG_rl_190 ;
	7'h2d :
		TR_134 = RG_rl_190 ;
	7'h2e :
		TR_134 = RG_rl_190 ;
	7'h2f :
		TR_134 = RG_rl_190 ;
	7'h30 :
		TR_134 = RG_rl_190 ;
	7'h31 :
		TR_134 = RG_rl_190 ;
	7'h32 :
		TR_134 = RG_rl_190 ;
	7'h33 :
		TR_134 = RG_rl_190 ;
	7'h34 :
		TR_134 = RG_rl_190 ;
	7'h35 :
		TR_134 = RG_rl_190 ;
	7'h36 :
		TR_134 = RG_rl_190 ;
	7'h37 :
		TR_134 = RG_rl_190 ;
	7'h38 :
		TR_134 = RG_rl_190 ;
	7'h39 :
		TR_134 = RG_rl_190 ;
	7'h3a :
		TR_134 = RG_rl_190 ;
	7'h3b :
		TR_134 = RG_rl_190 ;
	7'h3c :
		TR_134 = RG_rl_190 ;
	7'h3d :
		TR_134 = RG_rl_190 ;
	7'h3e :
		TR_134 = RG_rl_190 ;
	7'h3f :
		TR_134 = RG_rl_190 ;
	7'h40 :
		TR_134 = RG_rl_190 ;
	7'h41 :
		TR_134 = RG_rl_190 ;
	7'h42 :
		TR_134 = RG_rl_190 ;
	7'h43 :
		TR_134 = RG_rl_190 ;
	7'h44 :
		TR_134 = RG_rl_190 ;
	7'h45 :
		TR_134 = RG_rl_190 ;
	7'h46 :
		TR_134 = RG_rl_190 ;
	7'h47 :
		TR_134 = RG_rl_190 ;
	7'h48 :
		TR_134 = RG_rl_190 ;
	7'h49 :
		TR_134 = RG_rl_190 ;
	7'h4a :
		TR_134 = RG_rl_190 ;
	7'h4b :
		TR_134 = RG_rl_190 ;
	7'h4c :
		TR_134 = RG_rl_190 ;
	7'h4d :
		TR_134 = RG_rl_190 ;
	7'h4e :
		TR_134 = RG_rl_190 ;
	7'h4f :
		TR_134 = RG_rl_190 ;
	7'h50 :
		TR_134 = RG_rl_190 ;
	7'h51 :
		TR_134 = RG_rl_190 ;
	7'h52 :
		TR_134 = RG_rl_190 ;
	7'h53 :
		TR_134 = RG_rl_190 ;
	7'h54 :
		TR_134 = RG_rl_190 ;
	7'h55 :
		TR_134 = RG_rl_190 ;
	7'h56 :
		TR_134 = RG_rl_190 ;
	7'h57 :
		TR_134 = RG_rl_190 ;
	7'h58 :
		TR_134 = RG_rl_190 ;
	7'h59 :
		TR_134 = RG_rl_190 ;
	7'h5a :
		TR_134 = RG_rl_190 ;
	7'h5b :
		TR_134 = RG_rl_190 ;
	7'h5c :
		TR_134 = RG_rl_190 ;
	7'h5d :
		TR_134 = RG_rl_190 ;
	7'h5e :
		TR_134 = RG_rl_190 ;
	7'h5f :
		TR_134 = RG_rl_190 ;
	7'h60 :
		TR_134 = RG_rl_190 ;
	7'h61 :
		TR_134 = RG_rl_190 ;
	7'h62 :
		TR_134 = RG_rl_190 ;
	7'h63 :
		TR_134 = RG_rl_190 ;
	7'h64 :
		TR_134 = RG_rl_190 ;
	7'h65 :
		TR_134 = RG_rl_190 ;
	7'h66 :
		TR_134 = RG_rl_190 ;
	7'h67 :
		TR_134 = RG_rl_190 ;
	7'h68 :
		TR_134 = RG_rl_190 ;
	7'h69 :
		TR_134 = RG_rl_190 ;
	7'h6a :
		TR_134 = RG_rl_190 ;
	7'h6b :
		TR_134 = RG_rl_190 ;
	7'h6c :
		TR_134 = RG_rl_190 ;
	7'h6d :
		TR_134 = RG_rl_190 ;
	7'h6e :
		TR_134 = RG_rl_190 ;
	7'h6f :
		TR_134 = RG_rl_190 ;
	7'h70 :
		TR_134 = RG_rl_190 ;
	7'h71 :
		TR_134 = RG_rl_190 ;
	7'h72 :
		TR_134 = RG_rl_190 ;
	7'h73 :
		TR_134 = RG_rl_190 ;
	7'h74 :
		TR_134 = RG_rl_190 ;
	7'h75 :
		TR_134 = RG_rl_190 ;
	7'h76 :
		TR_134 = RG_rl_190 ;
	7'h77 :
		TR_134 = RG_rl_190 ;
	7'h78 :
		TR_134 = RG_rl_190 ;
	7'h79 :
		TR_134 = RG_rl_190 ;
	7'h7a :
		TR_134 = 9'h000 ;	// line#=../rle.cpp:79
	7'h7b :
		TR_134 = RG_rl_190 ;
	7'h7c :
		TR_134 = RG_rl_190 ;
	7'h7d :
		TR_134 = RG_rl_190 ;
	7'h7e :
		TR_134 = RG_rl_190 ;
	7'h7f :
		TR_134 = RG_rl_190 ;
	default :
		TR_134 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_59 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h01 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h02 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h03 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h04 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h05 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h06 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h07 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h08 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h09 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h0a :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h0b :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h0c :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h0d :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h0e :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h0f :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h10 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h11 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h12 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h13 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h14 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h15 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h16 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h17 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h18 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h19 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h1a :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h1b :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h1c :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h1d :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h1e :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h1f :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h20 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h21 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h22 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h23 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h24 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h25 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h26 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h27 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h28 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h29 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h2a :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h2b :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h2c :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h2d :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h2e :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h2f :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h30 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h31 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h32 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h33 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h34 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h35 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h36 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h37 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h38 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h39 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h3a :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h3b :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h3c :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h3d :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h3e :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h3f :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h40 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h41 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h42 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h43 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h44 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h45 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h46 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h47 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h48 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h49 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h4a :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h4b :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h4c :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h4d :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h4e :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h4f :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h50 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h51 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h52 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h53 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h54 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h55 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h56 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h57 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h58 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h59 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h5a :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h5b :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h5c :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h5d :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h5e :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h5f :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h60 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h61 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h62 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h63 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h64 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h65 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h66 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h67 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h68 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h69 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h6a :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h6b :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h6c :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h6d :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h6e :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h6f :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h70 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h71 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h72 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h73 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h74 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h75 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h76 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h77 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h78 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h79 :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h7a :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h7b :
		TR_135 = 9'h000 ;	// line#=../rle.cpp:79
	7'h7c :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h7d :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h7e :
		TR_135 = RG_quantized_block_rl_59 ;
	7'h7f :
		TR_135 = RG_quantized_block_rl_59 ;
	default :
		TR_135 = 9'hx ;
	endcase
always @ ( RG_rl_191 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_136 = RG_rl_191 ;
	7'h01 :
		TR_136 = RG_rl_191 ;
	7'h02 :
		TR_136 = RG_rl_191 ;
	7'h03 :
		TR_136 = RG_rl_191 ;
	7'h04 :
		TR_136 = RG_rl_191 ;
	7'h05 :
		TR_136 = RG_rl_191 ;
	7'h06 :
		TR_136 = RG_rl_191 ;
	7'h07 :
		TR_136 = RG_rl_191 ;
	7'h08 :
		TR_136 = RG_rl_191 ;
	7'h09 :
		TR_136 = RG_rl_191 ;
	7'h0a :
		TR_136 = RG_rl_191 ;
	7'h0b :
		TR_136 = RG_rl_191 ;
	7'h0c :
		TR_136 = RG_rl_191 ;
	7'h0d :
		TR_136 = RG_rl_191 ;
	7'h0e :
		TR_136 = RG_rl_191 ;
	7'h0f :
		TR_136 = RG_rl_191 ;
	7'h10 :
		TR_136 = RG_rl_191 ;
	7'h11 :
		TR_136 = RG_rl_191 ;
	7'h12 :
		TR_136 = RG_rl_191 ;
	7'h13 :
		TR_136 = RG_rl_191 ;
	7'h14 :
		TR_136 = RG_rl_191 ;
	7'h15 :
		TR_136 = RG_rl_191 ;
	7'h16 :
		TR_136 = RG_rl_191 ;
	7'h17 :
		TR_136 = RG_rl_191 ;
	7'h18 :
		TR_136 = RG_rl_191 ;
	7'h19 :
		TR_136 = RG_rl_191 ;
	7'h1a :
		TR_136 = RG_rl_191 ;
	7'h1b :
		TR_136 = RG_rl_191 ;
	7'h1c :
		TR_136 = RG_rl_191 ;
	7'h1d :
		TR_136 = RG_rl_191 ;
	7'h1e :
		TR_136 = RG_rl_191 ;
	7'h1f :
		TR_136 = RG_rl_191 ;
	7'h20 :
		TR_136 = RG_rl_191 ;
	7'h21 :
		TR_136 = RG_rl_191 ;
	7'h22 :
		TR_136 = RG_rl_191 ;
	7'h23 :
		TR_136 = RG_rl_191 ;
	7'h24 :
		TR_136 = RG_rl_191 ;
	7'h25 :
		TR_136 = RG_rl_191 ;
	7'h26 :
		TR_136 = RG_rl_191 ;
	7'h27 :
		TR_136 = RG_rl_191 ;
	7'h28 :
		TR_136 = RG_rl_191 ;
	7'h29 :
		TR_136 = RG_rl_191 ;
	7'h2a :
		TR_136 = RG_rl_191 ;
	7'h2b :
		TR_136 = RG_rl_191 ;
	7'h2c :
		TR_136 = RG_rl_191 ;
	7'h2d :
		TR_136 = RG_rl_191 ;
	7'h2e :
		TR_136 = RG_rl_191 ;
	7'h2f :
		TR_136 = RG_rl_191 ;
	7'h30 :
		TR_136 = RG_rl_191 ;
	7'h31 :
		TR_136 = RG_rl_191 ;
	7'h32 :
		TR_136 = RG_rl_191 ;
	7'h33 :
		TR_136 = RG_rl_191 ;
	7'h34 :
		TR_136 = RG_rl_191 ;
	7'h35 :
		TR_136 = RG_rl_191 ;
	7'h36 :
		TR_136 = RG_rl_191 ;
	7'h37 :
		TR_136 = RG_rl_191 ;
	7'h38 :
		TR_136 = RG_rl_191 ;
	7'h39 :
		TR_136 = RG_rl_191 ;
	7'h3a :
		TR_136 = RG_rl_191 ;
	7'h3b :
		TR_136 = RG_rl_191 ;
	7'h3c :
		TR_136 = RG_rl_191 ;
	7'h3d :
		TR_136 = RG_rl_191 ;
	7'h3e :
		TR_136 = RG_rl_191 ;
	7'h3f :
		TR_136 = RG_rl_191 ;
	7'h40 :
		TR_136 = RG_rl_191 ;
	7'h41 :
		TR_136 = RG_rl_191 ;
	7'h42 :
		TR_136 = RG_rl_191 ;
	7'h43 :
		TR_136 = RG_rl_191 ;
	7'h44 :
		TR_136 = RG_rl_191 ;
	7'h45 :
		TR_136 = RG_rl_191 ;
	7'h46 :
		TR_136 = RG_rl_191 ;
	7'h47 :
		TR_136 = RG_rl_191 ;
	7'h48 :
		TR_136 = RG_rl_191 ;
	7'h49 :
		TR_136 = RG_rl_191 ;
	7'h4a :
		TR_136 = RG_rl_191 ;
	7'h4b :
		TR_136 = RG_rl_191 ;
	7'h4c :
		TR_136 = RG_rl_191 ;
	7'h4d :
		TR_136 = RG_rl_191 ;
	7'h4e :
		TR_136 = RG_rl_191 ;
	7'h4f :
		TR_136 = RG_rl_191 ;
	7'h50 :
		TR_136 = RG_rl_191 ;
	7'h51 :
		TR_136 = RG_rl_191 ;
	7'h52 :
		TR_136 = RG_rl_191 ;
	7'h53 :
		TR_136 = RG_rl_191 ;
	7'h54 :
		TR_136 = RG_rl_191 ;
	7'h55 :
		TR_136 = RG_rl_191 ;
	7'h56 :
		TR_136 = RG_rl_191 ;
	7'h57 :
		TR_136 = RG_rl_191 ;
	7'h58 :
		TR_136 = RG_rl_191 ;
	7'h59 :
		TR_136 = RG_rl_191 ;
	7'h5a :
		TR_136 = RG_rl_191 ;
	7'h5b :
		TR_136 = RG_rl_191 ;
	7'h5c :
		TR_136 = RG_rl_191 ;
	7'h5d :
		TR_136 = RG_rl_191 ;
	7'h5e :
		TR_136 = RG_rl_191 ;
	7'h5f :
		TR_136 = RG_rl_191 ;
	7'h60 :
		TR_136 = RG_rl_191 ;
	7'h61 :
		TR_136 = RG_rl_191 ;
	7'h62 :
		TR_136 = RG_rl_191 ;
	7'h63 :
		TR_136 = RG_rl_191 ;
	7'h64 :
		TR_136 = RG_rl_191 ;
	7'h65 :
		TR_136 = RG_rl_191 ;
	7'h66 :
		TR_136 = RG_rl_191 ;
	7'h67 :
		TR_136 = RG_rl_191 ;
	7'h68 :
		TR_136 = RG_rl_191 ;
	7'h69 :
		TR_136 = RG_rl_191 ;
	7'h6a :
		TR_136 = RG_rl_191 ;
	7'h6b :
		TR_136 = RG_rl_191 ;
	7'h6c :
		TR_136 = RG_rl_191 ;
	7'h6d :
		TR_136 = RG_rl_191 ;
	7'h6e :
		TR_136 = RG_rl_191 ;
	7'h6f :
		TR_136 = RG_rl_191 ;
	7'h70 :
		TR_136 = RG_rl_191 ;
	7'h71 :
		TR_136 = RG_rl_191 ;
	7'h72 :
		TR_136 = RG_rl_191 ;
	7'h73 :
		TR_136 = RG_rl_191 ;
	7'h74 :
		TR_136 = RG_rl_191 ;
	7'h75 :
		TR_136 = RG_rl_191 ;
	7'h76 :
		TR_136 = RG_rl_191 ;
	7'h77 :
		TR_136 = RG_rl_191 ;
	7'h78 :
		TR_136 = RG_rl_191 ;
	7'h79 :
		TR_136 = RG_rl_191 ;
	7'h7a :
		TR_136 = RG_rl_191 ;
	7'h7b :
		TR_136 = RG_rl_191 ;
	7'h7c :
		TR_136 = 9'h000 ;	// line#=../rle.cpp:79
	7'h7d :
		TR_136 = RG_rl_191 ;
	7'h7e :
		TR_136 = RG_rl_191 ;
	7'h7f :
		TR_136 = RG_rl_191 ;
	default :
		TR_136 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_60 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h01 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h02 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h03 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h04 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h05 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h06 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h07 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h08 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h09 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h0a :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h0b :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h0c :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h0d :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h0e :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h0f :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h10 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h11 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h12 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h13 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h14 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h15 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h16 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h17 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h18 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h19 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h1a :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h1b :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h1c :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h1d :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h1e :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h1f :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h20 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h21 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h22 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h23 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h24 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h25 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h26 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h27 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h28 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h29 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h2a :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h2b :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h2c :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h2d :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h2e :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h2f :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h30 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h31 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h32 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h33 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h34 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h35 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h36 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h37 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h38 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h39 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h3a :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h3b :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h3c :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h3d :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h3e :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h3f :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h40 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h41 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h42 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h43 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h44 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h45 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h46 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h47 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h48 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h49 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h4a :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h4b :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h4c :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h4d :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h4e :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h4f :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h50 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h51 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h52 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h53 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h54 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h55 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h56 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h57 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h58 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h59 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h5a :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h5b :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h5c :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h5d :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h5e :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h5f :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h60 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h61 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h62 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h63 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h64 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h65 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h66 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h67 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h68 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h69 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h6a :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h6b :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h6c :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h6d :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h6e :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h6f :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h70 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h71 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h72 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h73 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h74 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h75 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h76 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h77 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h78 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h79 :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h7a :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h7b :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h7c :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h7d :
		TR_137 = 9'h000 ;	// line#=../rle.cpp:79
	7'h7e :
		TR_137 = RG_quantized_block_rl_60 ;
	7'h7f :
		TR_137 = RG_quantized_block_rl_60 ;
	default :
		TR_137 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_61 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h01 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h02 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h03 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h04 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h05 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h06 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h07 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h08 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h09 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h0a :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h0b :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h0c :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h0d :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h0e :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h0f :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h10 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h11 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h12 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h13 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h14 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h15 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h16 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h17 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h18 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h19 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h1a :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h1b :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h1c :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h1d :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h1e :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h1f :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h20 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h21 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h22 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h23 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h24 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h25 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h26 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h27 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h28 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h29 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h2a :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h2b :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h2c :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h2d :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h2e :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h2f :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h30 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h31 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h32 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h33 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h34 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h35 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h36 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h37 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h38 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h39 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h3a :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h3b :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h3c :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h3d :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h3e :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h3f :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h40 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h41 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h42 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h43 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h44 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h45 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h46 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h47 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h48 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h49 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h4a :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h4b :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h4c :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h4d :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h4e :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h4f :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h50 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h51 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h52 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h53 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h54 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h55 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h56 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h57 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h58 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h59 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h5a :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h5b :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h5c :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h5d :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h5e :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h5f :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h60 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h61 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h62 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h63 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h64 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h65 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h66 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h67 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h68 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h69 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h6a :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h6b :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h6c :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h6d :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h6e :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h6f :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h70 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h71 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h72 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h73 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h74 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h75 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h76 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h77 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h78 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h79 :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h7a :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h7b :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h7c :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h7d :
		TR_138 = RG_quantized_block_rl_61 ;
	7'h7e :
		TR_138 = 9'h000 ;	// line#=../rle.cpp:79
	7'h7f :
		TR_138 = RG_quantized_block_rl_61 ;
	default :
		TR_138 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_len )	// line#=../rle.cpp:79
	case ( RG_len [6:0] )
	7'h00 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h01 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h02 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h03 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h04 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h05 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h06 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h07 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h08 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h09 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h0a :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h0b :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h0c :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h0d :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h0e :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h0f :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h10 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h11 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h12 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h13 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h14 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h15 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h16 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h17 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h18 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h19 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h1a :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h1b :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h1c :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h1d :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h1e :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h1f :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h20 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h21 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h22 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h23 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h24 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h25 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h26 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h27 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h28 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h29 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h2a :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h2b :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h2c :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h2d :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h2e :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h2f :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h30 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h31 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h32 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h33 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h34 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h35 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h36 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h37 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h38 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h39 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h3a :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h3b :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h3c :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h3d :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h3e :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h3f :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h40 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h41 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h42 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h43 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h44 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h45 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h46 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h47 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h48 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h49 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h4a :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h4b :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h4c :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h4d :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h4e :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h4f :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h50 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h51 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h52 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h53 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h54 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h55 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h56 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h57 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h58 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h59 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h5a :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h5b :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h5c :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h5d :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h5e :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h5f :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h60 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h61 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h62 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h63 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h64 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h65 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h66 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h67 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h68 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h69 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h6a :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h6b :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h6c :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h6d :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h6e :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h6f :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h70 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h71 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h72 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h73 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h74 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h75 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h76 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h77 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h78 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h79 :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h7a :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h7b :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h7c :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h7d :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h7e :
		rl_a127_t2 = RG_k_quantized_block_rl_01 ;
	7'h7f :
		rl_a127_t2 = 9'h000 ;	// line#=../rle.cpp:79
	default :
		rl_a127_t2 = 9'hx ;
	endcase
always @ ( RG_rl_127 or RG_rl_126 or RG_rl_125 or RG_rl_124 or RG_rl_123 or RG_rl_122 or 
	RG_rl_121 or RG_rl_120 or RG_rl_119 or RG_rl_118 or RG_rl_117 or RG_rl_116 or 
	RG_rl_115 or RG_rl_114 or RG_rl_113 or RG_rl_112 or RG_rl_111 or RG_rl_110 or 
	RG_rl_109 or RG_rl_108 or RG_rl_107 or RG_rl_106 or RG_rl_105 or RG_rl_104 or 
	RG_rl_103 or RG_rl_102 or RG_rl_101 or RG_rl_100 or RG_rl_99 or RG_rl_98 or 
	RG_rl_97 or RG_rl_96 or RG_rl_95 or RG_rl_94 or RG_rl_93 or RG_rl_92 or 
	RG_rl_91 or RG_rl_90 or RG_rl_89 or RG_rl_88 or RG_rl_87 or RG_rl_86 or 
	RG_rl_85 or RG_rl_84 or RG_rl_83 or RG_rl_82 or RG_rl_81 or RG_rl_80 or 
	RG_rl_79 or RG_rl_78 or RG_rl_77 or RG_rl_76 or RG_rl_75 or RG_rl_74 or 
	RG_rl_73 or RG_rl_72 or RG_rl_71 or RG_rl_70 or RG_rl_69 or RG_rl_68 or 
	RG_rl_67 or RG_rl_66 or RG_rl_65 or RG_rl_64 or RG_rl_63 or RG_rl_62 or 
	RG_rl_61 or RG_rl_60 or RG_rl_59 or RG_rl_58 or RG_rl_57 or RG_rl_56 or 
	RG_rl_55 or RG_rl_54 or RG_rl_53 or RG_rl_52 or RG_rl_51 or RG_rl_50 or 
	RG_rl_49 or RG_rl_48 or RG_rl_47 or RG_rl_46 or RG_rl_45 or RG_rl_44 or 
	RG_rl_43 or RG_rl_42 or RG_rl_41 or RG_rl_40 or RG_rl_39 or RG_rl_38 or 
	RG_rl_37 or RG_rl_36 or RG_rl_35 or RG_rl_34 or RG_rl_33 or RG_rl_32 or 
	RG_rl_31 or RG_rl_30 or RG_rl_29 or RG_rl_28 or RG_rl_27 or RG_rl_26 or 
	RG_rl_25 or RG_rl_24 or RG_rl_23 or RG_rl_22 or RG_rl_21 or RG_rl_20 or 
	RG_rl_19 or RG_rl_18 or RG_rl_17 or RG_rl_16 or RG_rl_15 or RG_rl_14 or 
	RG_rl_13 or RG_rl_12 or RG_rl_11 or RG_rl_10 or RG_rl_9 or RG_rl_8 or RG_rl_7 or 
	RG_rl_6 or RG_rl_5 or RG_rl_4 or RG_rl_3 or RG_rl_2 or RG_rl_1 or RG_rl or 
	sub8u_71ot )	// line#=../rle.cpp:83,84
	case ( sub8u_71ot )
	7'h00 :
		M_15_t128 = ~|{ RG_rl [8:4] , ~RG_rl [3:0] } ;	// line#=../rle.cpp:83,84
	7'h01 :
		M_15_t128 = ~|{ RG_rl_1 [8:4] , ~RG_rl_1 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h02 :
		M_15_t128 = ~|{ RG_rl_2 [8:4] , ~RG_rl_2 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h03 :
		M_15_t128 = ~|{ RG_rl_3 [8:4] , ~RG_rl_3 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h04 :
		M_15_t128 = ~|{ RG_rl_4 [8:4] , ~RG_rl_4 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h05 :
		M_15_t128 = ~|{ RG_rl_5 [8:4] , ~RG_rl_5 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h06 :
		M_15_t128 = ~|{ RG_rl_6 [8:4] , ~RG_rl_6 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h07 :
		M_15_t128 = ~|{ RG_rl_7 [8:4] , ~RG_rl_7 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h08 :
		M_15_t128 = ~|{ RG_rl_8 [8:4] , ~RG_rl_8 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h09 :
		M_15_t128 = ~|{ RG_rl_9 [8:4] , ~RG_rl_9 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0a :
		M_15_t128 = ~|{ RG_rl_10 [8:4] , ~RG_rl_10 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0b :
		M_15_t128 = ~|{ RG_rl_11 [8:4] , ~RG_rl_11 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0c :
		M_15_t128 = ~|{ RG_rl_12 [8:4] , ~RG_rl_12 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0d :
		M_15_t128 = ~|{ RG_rl_13 [8:4] , ~RG_rl_13 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0e :
		M_15_t128 = ~|{ RG_rl_14 [8:4] , ~RG_rl_14 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0f :
		M_15_t128 = ~|{ RG_rl_15 [8:4] , ~RG_rl_15 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h10 :
		M_15_t128 = ~|{ RG_rl_16 [8:4] , ~RG_rl_16 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h11 :
		M_15_t128 = ~|{ RG_rl_17 [8:4] , ~RG_rl_17 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h12 :
		M_15_t128 = ~|{ RG_rl_18 [8:4] , ~RG_rl_18 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h13 :
		M_15_t128 = ~|{ RG_rl_19 [8:4] , ~RG_rl_19 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h14 :
		M_15_t128 = ~|{ RG_rl_20 [8:4] , ~RG_rl_20 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h15 :
		M_15_t128 = ~|{ RG_rl_21 [8:4] , ~RG_rl_21 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h16 :
		M_15_t128 = ~|{ RG_rl_22 [8:4] , ~RG_rl_22 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h17 :
		M_15_t128 = ~|{ RG_rl_23 [8:4] , ~RG_rl_23 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h18 :
		M_15_t128 = ~|{ RG_rl_24 [8:4] , ~RG_rl_24 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h19 :
		M_15_t128 = ~|{ RG_rl_25 [8:4] , ~RG_rl_25 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1a :
		M_15_t128 = ~|{ RG_rl_26 [8:4] , ~RG_rl_26 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1b :
		M_15_t128 = ~|{ RG_rl_27 [8:4] , ~RG_rl_27 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1c :
		M_15_t128 = ~|{ RG_rl_28 [8:4] , ~RG_rl_28 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1d :
		M_15_t128 = ~|{ RG_rl_29 [8:4] , ~RG_rl_29 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1e :
		M_15_t128 = ~|{ RG_rl_30 [8:4] , ~RG_rl_30 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1f :
		M_15_t128 = ~|{ RG_rl_31 [8:4] , ~RG_rl_31 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h20 :
		M_15_t128 = ~|{ RG_rl_32 [8:4] , ~RG_rl_32 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h21 :
		M_15_t128 = ~|{ RG_rl_33 [8:4] , ~RG_rl_33 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h22 :
		M_15_t128 = ~|{ RG_rl_34 [8:4] , ~RG_rl_34 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h23 :
		M_15_t128 = ~|{ RG_rl_35 [8:4] , ~RG_rl_35 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h24 :
		M_15_t128 = ~|{ RG_rl_36 [8:4] , ~RG_rl_36 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h25 :
		M_15_t128 = ~|{ RG_rl_37 [8:4] , ~RG_rl_37 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h26 :
		M_15_t128 = ~|{ RG_rl_38 [8:4] , ~RG_rl_38 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h27 :
		M_15_t128 = ~|{ RG_rl_39 [8:4] , ~RG_rl_39 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h28 :
		M_15_t128 = ~|{ RG_rl_40 [8:4] , ~RG_rl_40 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h29 :
		M_15_t128 = ~|{ RG_rl_41 [8:4] , ~RG_rl_41 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2a :
		M_15_t128 = ~|{ RG_rl_42 [8:4] , ~RG_rl_42 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2b :
		M_15_t128 = ~|{ RG_rl_43 [8:4] , ~RG_rl_43 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2c :
		M_15_t128 = ~|{ RG_rl_44 [8:4] , ~RG_rl_44 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2d :
		M_15_t128 = ~|{ RG_rl_45 [8:4] , ~RG_rl_45 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2e :
		M_15_t128 = ~|{ RG_rl_46 [8:4] , ~RG_rl_46 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2f :
		M_15_t128 = ~|{ RG_rl_47 [8:4] , ~RG_rl_47 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h30 :
		M_15_t128 = ~|{ RG_rl_48 [8:4] , ~RG_rl_48 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h31 :
		M_15_t128 = ~|{ RG_rl_49 [8:4] , ~RG_rl_49 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h32 :
		M_15_t128 = ~|{ RG_rl_50 [8:4] , ~RG_rl_50 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h33 :
		M_15_t128 = ~|{ RG_rl_51 [8:4] , ~RG_rl_51 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h34 :
		M_15_t128 = ~|{ RG_rl_52 [8:4] , ~RG_rl_52 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h35 :
		M_15_t128 = ~|{ RG_rl_53 [8:4] , ~RG_rl_53 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h36 :
		M_15_t128 = ~|{ RG_rl_54 [8:4] , ~RG_rl_54 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h37 :
		M_15_t128 = ~|{ RG_rl_55 [8:4] , ~RG_rl_55 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h38 :
		M_15_t128 = ~|{ RG_rl_56 [8:4] , ~RG_rl_56 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h39 :
		M_15_t128 = ~|{ RG_rl_57 [8:4] , ~RG_rl_57 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3a :
		M_15_t128 = ~|{ RG_rl_58 [8:4] , ~RG_rl_58 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3b :
		M_15_t128 = ~|{ RG_rl_59 [8:4] , ~RG_rl_59 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3c :
		M_15_t128 = ~|{ RG_rl_60 [8:4] , ~RG_rl_60 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3d :
		M_15_t128 = ~|{ RG_rl_61 [8:4] , ~RG_rl_61 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3e :
		M_15_t128 = ~|{ RG_rl_62 [8:4] , ~RG_rl_62 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3f :
		M_15_t128 = ~|{ RG_rl_63 [8:4] , ~RG_rl_63 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h40 :
		M_15_t128 = ~|{ RG_rl_64 [8:4] , ~RG_rl_64 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h41 :
		M_15_t128 = ~|{ RG_rl_65 [8:4] , ~RG_rl_65 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h42 :
		M_15_t128 = ~|{ RG_rl_66 [8:4] , ~RG_rl_66 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h43 :
		M_15_t128 = ~|{ RG_rl_67 [8:4] , ~RG_rl_67 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h44 :
		M_15_t128 = ~|{ RG_rl_68 [8:4] , ~RG_rl_68 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h45 :
		M_15_t128 = ~|{ RG_rl_69 [8:4] , ~RG_rl_69 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h46 :
		M_15_t128 = ~|{ RG_rl_70 [8:4] , ~RG_rl_70 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h47 :
		M_15_t128 = ~|{ RG_rl_71 [8:4] , ~RG_rl_71 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h48 :
		M_15_t128 = ~|{ RG_rl_72 [8:4] , ~RG_rl_72 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h49 :
		M_15_t128 = ~|{ RG_rl_73 [8:4] , ~RG_rl_73 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4a :
		M_15_t128 = ~|{ RG_rl_74 [8:4] , ~RG_rl_74 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4b :
		M_15_t128 = ~|{ RG_rl_75 [8:4] , ~RG_rl_75 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4c :
		M_15_t128 = ~|{ RG_rl_76 [8:4] , ~RG_rl_76 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4d :
		M_15_t128 = ~|{ RG_rl_77 [8:4] , ~RG_rl_77 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4e :
		M_15_t128 = ~|{ RG_rl_78 [8:4] , ~RG_rl_78 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4f :
		M_15_t128 = ~|{ RG_rl_79 [8:4] , ~RG_rl_79 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h50 :
		M_15_t128 = ~|{ RG_rl_80 [8:4] , ~RG_rl_80 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h51 :
		M_15_t128 = ~|{ RG_rl_81 [8:4] , ~RG_rl_81 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h52 :
		M_15_t128 = ~|{ RG_rl_82 [8:4] , ~RG_rl_82 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h53 :
		M_15_t128 = ~|{ RG_rl_83 [8:4] , ~RG_rl_83 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h54 :
		M_15_t128 = ~|{ RG_rl_84 [8:4] , ~RG_rl_84 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h55 :
		M_15_t128 = ~|{ RG_rl_85 [8:4] , ~RG_rl_85 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h56 :
		M_15_t128 = ~|{ RG_rl_86 [8:4] , ~RG_rl_86 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h57 :
		M_15_t128 = ~|{ RG_rl_87 [8:4] , ~RG_rl_87 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h58 :
		M_15_t128 = ~|{ RG_rl_88 [8:4] , ~RG_rl_88 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h59 :
		M_15_t128 = ~|{ RG_rl_89 [8:4] , ~RG_rl_89 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5a :
		M_15_t128 = ~|{ RG_rl_90 [8:4] , ~RG_rl_90 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5b :
		M_15_t128 = ~|{ RG_rl_91 [8:4] , ~RG_rl_91 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5c :
		M_15_t128 = ~|{ RG_rl_92 [8:4] , ~RG_rl_92 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5d :
		M_15_t128 = ~|{ RG_rl_93 [8:4] , ~RG_rl_93 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5e :
		M_15_t128 = ~|{ RG_rl_94 [8:4] , ~RG_rl_94 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5f :
		M_15_t128 = ~|{ RG_rl_95 [8:4] , ~RG_rl_95 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h60 :
		M_15_t128 = ~|{ RG_rl_96 [8:4] , ~RG_rl_96 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h61 :
		M_15_t128 = ~|{ RG_rl_97 [8:4] , ~RG_rl_97 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h62 :
		M_15_t128 = ~|{ RG_rl_98 [8:4] , ~RG_rl_98 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h63 :
		M_15_t128 = ~|{ RG_rl_99 [8:4] , ~RG_rl_99 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h64 :
		M_15_t128 = ~|{ RG_rl_100 [8:4] , ~RG_rl_100 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h65 :
		M_15_t128 = ~|{ RG_rl_101 [8:4] , ~RG_rl_101 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h66 :
		M_15_t128 = ~|{ RG_rl_102 [8:4] , ~RG_rl_102 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h67 :
		M_15_t128 = ~|{ RG_rl_103 [8:4] , ~RG_rl_103 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h68 :
		M_15_t128 = ~|{ RG_rl_104 [8:4] , ~RG_rl_104 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h69 :
		M_15_t128 = ~|{ RG_rl_105 [8:4] , ~RG_rl_105 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6a :
		M_15_t128 = ~|{ RG_rl_106 [8:4] , ~RG_rl_106 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6b :
		M_15_t128 = ~|{ RG_rl_107 [8:4] , ~RG_rl_107 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6c :
		M_15_t128 = ~|{ RG_rl_108 [8:4] , ~RG_rl_108 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6d :
		M_15_t128 = ~|{ RG_rl_109 [8:4] , ~RG_rl_109 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6e :
		M_15_t128 = ~|{ RG_rl_110 [8:4] , ~RG_rl_110 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6f :
		M_15_t128 = ~|{ RG_rl_111 [8:4] , ~RG_rl_111 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h70 :
		M_15_t128 = ~|{ RG_rl_112 [8:4] , ~RG_rl_112 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h71 :
		M_15_t128 = ~|{ RG_rl_113 [8:4] , ~RG_rl_113 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h72 :
		M_15_t128 = ~|{ RG_rl_114 [8:4] , ~RG_rl_114 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h73 :
		M_15_t128 = ~|{ RG_rl_115 [8:4] , ~RG_rl_115 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h74 :
		M_15_t128 = ~|{ RG_rl_116 [8:4] , ~RG_rl_116 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h75 :
		M_15_t128 = ~|{ RG_rl_117 [8:4] , ~RG_rl_117 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h76 :
		M_15_t128 = ~|{ RG_rl_118 [8:4] , ~RG_rl_118 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h77 :
		M_15_t128 = ~|{ RG_rl_119 [8:4] , ~RG_rl_119 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h78 :
		M_15_t128 = ~|{ RG_rl_120 [8:4] , ~RG_rl_120 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h79 :
		M_15_t128 = ~|{ RG_rl_121 [8:4] , ~RG_rl_121 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7a :
		M_15_t128 = ~|{ RG_rl_122 [8:4] , ~RG_rl_122 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7b :
		M_15_t128 = ~|{ RG_rl_123 [8:4] , ~RG_rl_123 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7c :
		M_15_t128 = ~|{ RG_rl_124 [8:4] , ~RG_rl_124 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7d :
		M_15_t128 = ~|{ RG_rl_125 [8:4] , ~RG_rl_125 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7e :
		M_15_t128 = ~|{ RG_rl_126 [8:4] , ~RG_rl_126 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7f :
		M_15_t128 = ~|{ RG_rl_127 [8:4] , ~RG_rl_127 [3:0] } ;	// line#=../rle.cpp:83,84
	default :
		M_15_t128 = 1'hx ;
	endcase
always @ ( RG_zz_62 or RG_zz_61 or RG_zz_60 or RG_zz_59 or RG_zz_58 or RG_zz_57 or 
	RG_zz_56 or RG_zz_55 or RG_zz_54 or RG_zz_53 or RG_zz_52 or RG_zz_51 or 
	RG_zz_50 or RG_zz_49 or RG_zz_48 or RG_zz_47 or RG_zz_46 or RG_zz_45 or 
	RG_zz_44 or RG_zz_43 or RG_zz_42 or RG_zz_41 or RG_zz_40 or RG_zz_39 or 
	RG_zz_38 or RG_zz_37 or RG_zz_36 or RG_zz_35 or RG_zz_34 or RG_zz_33 or 
	RG_zz_32 or RG_zz_31 or RG_zz_30 or RG_zz_29 or RG_zz_28 or RG_zz_27 or 
	RG_zz_26 or RG_zz_25 or RG_zz_24 or RG_zz_23 or RG_zz_22 or RG_zz_21 or 
	RG_zz_20 or RG_zz_19 or RG_zz_18 or RG_zz_17 or RG_zz_16 or RG_zz_15 or 
	RG_zz_14 or RG_zz_13 or RG_zz_12 or RG_zz_11 or RG_zz_10 or RG_zz_9 or RG_zz_8 or 
	RG_zz_7 or RG_zz_6 or RG_zz_5 or RG_zz_4 or RG_zz_3 or RG_zz_2 or RG_zz_1 or 
	RG_zz or RG_quantized_block_rl_zz or RG_i_j_01 )	// line#=../rle.cpp:74
	case ( RG_i_j_01 [5:0] )
	6'h00 :
		M_16_t = RG_quantized_block_rl_zz ;	// line#=../rle.cpp:74
	6'h01 :
		M_16_t = RG_zz ;	// line#=../rle.cpp:74
	6'h02 :
		M_16_t = RG_zz_1 ;	// line#=../rle.cpp:74
	6'h03 :
		M_16_t = RG_zz_2 ;	// line#=../rle.cpp:74
	6'h04 :
		M_16_t = RG_zz_3 ;	// line#=../rle.cpp:74
	6'h05 :
		M_16_t = RG_zz_4 ;	// line#=../rle.cpp:74
	6'h06 :
		M_16_t = RG_zz_5 ;	// line#=../rle.cpp:74
	6'h07 :
		M_16_t = RG_zz_6 ;	// line#=../rle.cpp:74
	6'h08 :
		M_16_t = RG_zz_7 ;	// line#=../rle.cpp:74
	6'h09 :
		M_16_t = RG_zz_8 ;	// line#=../rle.cpp:74
	6'h0a :
		M_16_t = RG_zz_9 ;	// line#=../rle.cpp:74
	6'h0b :
		M_16_t = RG_zz_10 ;	// line#=../rle.cpp:74
	6'h0c :
		M_16_t = RG_zz_11 ;	// line#=../rle.cpp:74
	6'h0d :
		M_16_t = RG_zz_12 ;	// line#=../rle.cpp:74
	6'h0e :
		M_16_t = RG_zz_13 ;	// line#=../rle.cpp:74
	6'h0f :
		M_16_t = RG_zz_14 ;	// line#=../rle.cpp:74
	6'h10 :
		M_16_t = RG_zz_15 ;	// line#=../rle.cpp:74
	6'h11 :
		M_16_t = RG_zz_16 ;	// line#=../rle.cpp:74
	6'h12 :
		M_16_t = RG_zz_17 ;	// line#=../rle.cpp:74
	6'h13 :
		M_16_t = RG_zz_18 ;	// line#=../rle.cpp:74
	6'h14 :
		M_16_t = RG_zz_19 ;	// line#=../rle.cpp:74
	6'h15 :
		M_16_t = RG_zz_20 ;	// line#=../rle.cpp:74
	6'h16 :
		M_16_t = RG_zz_21 ;	// line#=../rle.cpp:74
	6'h17 :
		M_16_t = RG_zz_22 ;	// line#=../rle.cpp:74
	6'h18 :
		M_16_t = RG_zz_23 ;	// line#=../rle.cpp:74
	6'h19 :
		M_16_t = RG_zz_24 ;	// line#=../rle.cpp:74
	6'h1a :
		M_16_t = RG_zz_25 ;	// line#=../rle.cpp:74
	6'h1b :
		M_16_t = RG_zz_26 ;	// line#=../rle.cpp:74
	6'h1c :
		M_16_t = RG_zz_27 ;	// line#=../rle.cpp:74
	6'h1d :
		M_16_t = RG_zz_28 ;	// line#=../rle.cpp:74
	6'h1e :
		M_16_t = RG_zz_29 ;	// line#=../rle.cpp:74
	6'h1f :
		M_16_t = RG_zz_30 ;	// line#=../rle.cpp:74
	6'h20 :
		M_16_t = RG_zz_31 ;	// line#=../rle.cpp:74
	6'h21 :
		M_16_t = RG_zz_32 ;	// line#=../rle.cpp:74
	6'h22 :
		M_16_t = RG_zz_33 ;	// line#=../rle.cpp:74
	6'h23 :
		M_16_t = RG_zz_34 ;	// line#=../rle.cpp:74
	6'h24 :
		M_16_t = RG_zz_35 ;	// line#=../rle.cpp:74
	6'h25 :
		M_16_t = RG_zz_36 ;	// line#=../rle.cpp:74
	6'h26 :
		M_16_t = RG_zz_37 ;	// line#=../rle.cpp:74
	6'h27 :
		M_16_t = RG_zz_38 ;	// line#=../rle.cpp:74
	6'h28 :
		M_16_t = RG_zz_39 ;	// line#=../rle.cpp:74
	6'h29 :
		M_16_t = RG_zz_40 ;	// line#=../rle.cpp:74
	6'h2a :
		M_16_t = RG_zz_41 ;	// line#=../rle.cpp:74
	6'h2b :
		M_16_t = RG_zz_42 ;	// line#=../rle.cpp:74
	6'h2c :
		M_16_t = RG_zz_43 ;	// line#=../rle.cpp:74
	6'h2d :
		M_16_t = RG_zz_44 ;	// line#=../rle.cpp:74
	6'h2e :
		M_16_t = RG_zz_45 ;	// line#=../rle.cpp:74
	6'h2f :
		M_16_t = RG_zz_46 ;	// line#=../rle.cpp:74
	6'h30 :
		M_16_t = RG_zz_47 ;	// line#=../rle.cpp:74
	6'h31 :
		M_16_t = RG_zz_48 ;	// line#=../rle.cpp:74
	6'h32 :
		M_16_t = RG_zz_49 ;	// line#=../rle.cpp:74
	6'h33 :
		M_16_t = RG_zz_50 ;	// line#=../rle.cpp:74
	6'h34 :
		M_16_t = RG_zz_51 ;	// line#=../rle.cpp:74
	6'h35 :
		M_16_t = RG_zz_52 ;	// line#=../rle.cpp:74
	6'h36 :
		M_16_t = RG_zz_53 ;	// line#=../rle.cpp:74
	6'h37 :
		M_16_t = RG_zz_54 ;	// line#=../rle.cpp:74
	6'h38 :
		M_16_t = RG_zz_55 ;	// line#=../rle.cpp:74
	6'h39 :
		M_16_t = RG_zz_56 ;	// line#=../rle.cpp:74
	6'h3a :
		M_16_t = RG_zz_57 ;	// line#=../rle.cpp:74
	6'h3b :
		M_16_t = RG_zz_58 ;	// line#=../rle.cpp:74
	6'h3c :
		M_16_t = RG_zz_59 ;	// line#=../rle.cpp:74
	6'h3d :
		M_16_t = RG_zz_60 ;	// line#=../rle.cpp:74
	6'h3e :
		M_16_t = RG_zz_61 ;	// line#=../rle.cpp:74
	6'h3f :
		M_16_t = RG_zz_62 ;	// line#=../rle.cpp:74
	default :
		M_16_t = 9'hx ;
	endcase
always @ ( RG_previous_dc_rl or RG_k_quantized_block_rl_01 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a00_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h01 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h02 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h03 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h04 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h05 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h06 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h07 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h08 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h09 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h0a :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h0b :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h0c :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h0d :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h0e :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h0f :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h10 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h11 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h12 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h13 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h14 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h15 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h16 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h17 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h18 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h19 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h1a :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h1b :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h1c :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h1d :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h1e :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h1f :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h20 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h21 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h22 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h23 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h24 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h25 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h26 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h27 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h28 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h29 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h2a :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h2b :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h2c :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h2d :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h2e :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h2f :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h30 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h31 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h32 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h33 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h34 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h35 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h36 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h37 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h38 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h39 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h3a :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h3b :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h3c :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h3d :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h3e :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h3f :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h40 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h41 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h42 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h43 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h44 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h45 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h46 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h47 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h48 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h49 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h4a :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h4b :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h4c :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h4d :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h4e :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h4f :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h50 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h51 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h52 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h53 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h54 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h55 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h56 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h57 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h58 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h59 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h5a :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h5b :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h5c :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h5d :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h5e :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h5f :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h60 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h61 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h62 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h63 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h64 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h65 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h66 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h67 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h68 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h69 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h6a :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h6b :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h6c :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h6d :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h6e :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h6f :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h70 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h71 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h72 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h73 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h74 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h75 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h76 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h77 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h78 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h79 :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h7a :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h7b :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h7c :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h7d :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h7e :
		rl_a00_t8 = RG_previous_dc_rl ;
	7'h7f :
		rl_a00_t8 = RG_previous_dc_rl ;
	default :
		rl_a00_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_128 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a01_t8 = RG_rl_128 ;
	7'h01 :
		rl_a01_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h02 :
		rl_a01_t8 = RG_rl_128 ;
	7'h03 :
		rl_a01_t8 = RG_rl_128 ;
	7'h04 :
		rl_a01_t8 = RG_rl_128 ;
	7'h05 :
		rl_a01_t8 = RG_rl_128 ;
	7'h06 :
		rl_a01_t8 = RG_rl_128 ;
	7'h07 :
		rl_a01_t8 = RG_rl_128 ;
	7'h08 :
		rl_a01_t8 = RG_rl_128 ;
	7'h09 :
		rl_a01_t8 = RG_rl_128 ;
	7'h0a :
		rl_a01_t8 = RG_rl_128 ;
	7'h0b :
		rl_a01_t8 = RG_rl_128 ;
	7'h0c :
		rl_a01_t8 = RG_rl_128 ;
	7'h0d :
		rl_a01_t8 = RG_rl_128 ;
	7'h0e :
		rl_a01_t8 = RG_rl_128 ;
	7'h0f :
		rl_a01_t8 = RG_rl_128 ;
	7'h10 :
		rl_a01_t8 = RG_rl_128 ;
	7'h11 :
		rl_a01_t8 = RG_rl_128 ;
	7'h12 :
		rl_a01_t8 = RG_rl_128 ;
	7'h13 :
		rl_a01_t8 = RG_rl_128 ;
	7'h14 :
		rl_a01_t8 = RG_rl_128 ;
	7'h15 :
		rl_a01_t8 = RG_rl_128 ;
	7'h16 :
		rl_a01_t8 = RG_rl_128 ;
	7'h17 :
		rl_a01_t8 = RG_rl_128 ;
	7'h18 :
		rl_a01_t8 = RG_rl_128 ;
	7'h19 :
		rl_a01_t8 = RG_rl_128 ;
	7'h1a :
		rl_a01_t8 = RG_rl_128 ;
	7'h1b :
		rl_a01_t8 = RG_rl_128 ;
	7'h1c :
		rl_a01_t8 = RG_rl_128 ;
	7'h1d :
		rl_a01_t8 = RG_rl_128 ;
	7'h1e :
		rl_a01_t8 = RG_rl_128 ;
	7'h1f :
		rl_a01_t8 = RG_rl_128 ;
	7'h20 :
		rl_a01_t8 = RG_rl_128 ;
	7'h21 :
		rl_a01_t8 = RG_rl_128 ;
	7'h22 :
		rl_a01_t8 = RG_rl_128 ;
	7'h23 :
		rl_a01_t8 = RG_rl_128 ;
	7'h24 :
		rl_a01_t8 = RG_rl_128 ;
	7'h25 :
		rl_a01_t8 = RG_rl_128 ;
	7'h26 :
		rl_a01_t8 = RG_rl_128 ;
	7'h27 :
		rl_a01_t8 = RG_rl_128 ;
	7'h28 :
		rl_a01_t8 = RG_rl_128 ;
	7'h29 :
		rl_a01_t8 = RG_rl_128 ;
	7'h2a :
		rl_a01_t8 = RG_rl_128 ;
	7'h2b :
		rl_a01_t8 = RG_rl_128 ;
	7'h2c :
		rl_a01_t8 = RG_rl_128 ;
	7'h2d :
		rl_a01_t8 = RG_rl_128 ;
	7'h2e :
		rl_a01_t8 = RG_rl_128 ;
	7'h2f :
		rl_a01_t8 = RG_rl_128 ;
	7'h30 :
		rl_a01_t8 = RG_rl_128 ;
	7'h31 :
		rl_a01_t8 = RG_rl_128 ;
	7'h32 :
		rl_a01_t8 = RG_rl_128 ;
	7'h33 :
		rl_a01_t8 = RG_rl_128 ;
	7'h34 :
		rl_a01_t8 = RG_rl_128 ;
	7'h35 :
		rl_a01_t8 = RG_rl_128 ;
	7'h36 :
		rl_a01_t8 = RG_rl_128 ;
	7'h37 :
		rl_a01_t8 = RG_rl_128 ;
	7'h38 :
		rl_a01_t8 = RG_rl_128 ;
	7'h39 :
		rl_a01_t8 = RG_rl_128 ;
	7'h3a :
		rl_a01_t8 = RG_rl_128 ;
	7'h3b :
		rl_a01_t8 = RG_rl_128 ;
	7'h3c :
		rl_a01_t8 = RG_rl_128 ;
	7'h3d :
		rl_a01_t8 = RG_rl_128 ;
	7'h3e :
		rl_a01_t8 = RG_rl_128 ;
	7'h3f :
		rl_a01_t8 = RG_rl_128 ;
	7'h40 :
		rl_a01_t8 = RG_rl_128 ;
	7'h41 :
		rl_a01_t8 = RG_rl_128 ;
	7'h42 :
		rl_a01_t8 = RG_rl_128 ;
	7'h43 :
		rl_a01_t8 = RG_rl_128 ;
	7'h44 :
		rl_a01_t8 = RG_rl_128 ;
	7'h45 :
		rl_a01_t8 = RG_rl_128 ;
	7'h46 :
		rl_a01_t8 = RG_rl_128 ;
	7'h47 :
		rl_a01_t8 = RG_rl_128 ;
	7'h48 :
		rl_a01_t8 = RG_rl_128 ;
	7'h49 :
		rl_a01_t8 = RG_rl_128 ;
	7'h4a :
		rl_a01_t8 = RG_rl_128 ;
	7'h4b :
		rl_a01_t8 = RG_rl_128 ;
	7'h4c :
		rl_a01_t8 = RG_rl_128 ;
	7'h4d :
		rl_a01_t8 = RG_rl_128 ;
	7'h4e :
		rl_a01_t8 = RG_rl_128 ;
	7'h4f :
		rl_a01_t8 = RG_rl_128 ;
	7'h50 :
		rl_a01_t8 = RG_rl_128 ;
	7'h51 :
		rl_a01_t8 = RG_rl_128 ;
	7'h52 :
		rl_a01_t8 = RG_rl_128 ;
	7'h53 :
		rl_a01_t8 = RG_rl_128 ;
	7'h54 :
		rl_a01_t8 = RG_rl_128 ;
	7'h55 :
		rl_a01_t8 = RG_rl_128 ;
	7'h56 :
		rl_a01_t8 = RG_rl_128 ;
	7'h57 :
		rl_a01_t8 = RG_rl_128 ;
	7'h58 :
		rl_a01_t8 = RG_rl_128 ;
	7'h59 :
		rl_a01_t8 = RG_rl_128 ;
	7'h5a :
		rl_a01_t8 = RG_rl_128 ;
	7'h5b :
		rl_a01_t8 = RG_rl_128 ;
	7'h5c :
		rl_a01_t8 = RG_rl_128 ;
	7'h5d :
		rl_a01_t8 = RG_rl_128 ;
	7'h5e :
		rl_a01_t8 = RG_rl_128 ;
	7'h5f :
		rl_a01_t8 = RG_rl_128 ;
	7'h60 :
		rl_a01_t8 = RG_rl_128 ;
	7'h61 :
		rl_a01_t8 = RG_rl_128 ;
	7'h62 :
		rl_a01_t8 = RG_rl_128 ;
	7'h63 :
		rl_a01_t8 = RG_rl_128 ;
	7'h64 :
		rl_a01_t8 = RG_rl_128 ;
	7'h65 :
		rl_a01_t8 = RG_rl_128 ;
	7'h66 :
		rl_a01_t8 = RG_rl_128 ;
	7'h67 :
		rl_a01_t8 = RG_rl_128 ;
	7'h68 :
		rl_a01_t8 = RG_rl_128 ;
	7'h69 :
		rl_a01_t8 = RG_rl_128 ;
	7'h6a :
		rl_a01_t8 = RG_rl_128 ;
	7'h6b :
		rl_a01_t8 = RG_rl_128 ;
	7'h6c :
		rl_a01_t8 = RG_rl_128 ;
	7'h6d :
		rl_a01_t8 = RG_rl_128 ;
	7'h6e :
		rl_a01_t8 = RG_rl_128 ;
	7'h6f :
		rl_a01_t8 = RG_rl_128 ;
	7'h70 :
		rl_a01_t8 = RG_rl_128 ;
	7'h71 :
		rl_a01_t8 = RG_rl_128 ;
	7'h72 :
		rl_a01_t8 = RG_rl_128 ;
	7'h73 :
		rl_a01_t8 = RG_rl_128 ;
	7'h74 :
		rl_a01_t8 = RG_rl_128 ;
	7'h75 :
		rl_a01_t8 = RG_rl_128 ;
	7'h76 :
		rl_a01_t8 = RG_rl_128 ;
	7'h77 :
		rl_a01_t8 = RG_rl_128 ;
	7'h78 :
		rl_a01_t8 = RG_rl_128 ;
	7'h79 :
		rl_a01_t8 = RG_rl_128 ;
	7'h7a :
		rl_a01_t8 = RG_rl_128 ;
	7'h7b :
		rl_a01_t8 = RG_rl_128 ;
	7'h7c :
		rl_a01_t8 = RG_rl_128 ;
	7'h7d :
		rl_a01_t8 = RG_rl_128 ;
	7'h7e :
		rl_a01_t8 = RG_rl_128 ;
	7'h7f :
		rl_a01_t8 = RG_rl_128 ;
	default :
		rl_a01_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_129 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a02_t8 = RG_rl_129 ;
	7'h01 :
		rl_a02_t8 = RG_rl_129 ;
	7'h02 :
		rl_a02_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h03 :
		rl_a02_t8 = RG_rl_129 ;
	7'h04 :
		rl_a02_t8 = RG_rl_129 ;
	7'h05 :
		rl_a02_t8 = RG_rl_129 ;
	7'h06 :
		rl_a02_t8 = RG_rl_129 ;
	7'h07 :
		rl_a02_t8 = RG_rl_129 ;
	7'h08 :
		rl_a02_t8 = RG_rl_129 ;
	7'h09 :
		rl_a02_t8 = RG_rl_129 ;
	7'h0a :
		rl_a02_t8 = RG_rl_129 ;
	7'h0b :
		rl_a02_t8 = RG_rl_129 ;
	7'h0c :
		rl_a02_t8 = RG_rl_129 ;
	7'h0d :
		rl_a02_t8 = RG_rl_129 ;
	7'h0e :
		rl_a02_t8 = RG_rl_129 ;
	7'h0f :
		rl_a02_t8 = RG_rl_129 ;
	7'h10 :
		rl_a02_t8 = RG_rl_129 ;
	7'h11 :
		rl_a02_t8 = RG_rl_129 ;
	7'h12 :
		rl_a02_t8 = RG_rl_129 ;
	7'h13 :
		rl_a02_t8 = RG_rl_129 ;
	7'h14 :
		rl_a02_t8 = RG_rl_129 ;
	7'h15 :
		rl_a02_t8 = RG_rl_129 ;
	7'h16 :
		rl_a02_t8 = RG_rl_129 ;
	7'h17 :
		rl_a02_t8 = RG_rl_129 ;
	7'h18 :
		rl_a02_t8 = RG_rl_129 ;
	7'h19 :
		rl_a02_t8 = RG_rl_129 ;
	7'h1a :
		rl_a02_t8 = RG_rl_129 ;
	7'h1b :
		rl_a02_t8 = RG_rl_129 ;
	7'h1c :
		rl_a02_t8 = RG_rl_129 ;
	7'h1d :
		rl_a02_t8 = RG_rl_129 ;
	7'h1e :
		rl_a02_t8 = RG_rl_129 ;
	7'h1f :
		rl_a02_t8 = RG_rl_129 ;
	7'h20 :
		rl_a02_t8 = RG_rl_129 ;
	7'h21 :
		rl_a02_t8 = RG_rl_129 ;
	7'h22 :
		rl_a02_t8 = RG_rl_129 ;
	7'h23 :
		rl_a02_t8 = RG_rl_129 ;
	7'h24 :
		rl_a02_t8 = RG_rl_129 ;
	7'h25 :
		rl_a02_t8 = RG_rl_129 ;
	7'h26 :
		rl_a02_t8 = RG_rl_129 ;
	7'h27 :
		rl_a02_t8 = RG_rl_129 ;
	7'h28 :
		rl_a02_t8 = RG_rl_129 ;
	7'h29 :
		rl_a02_t8 = RG_rl_129 ;
	7'h2a :
		rl_a02_t8 = RG_rl_129 ;
	7'h2b :
		rl_a02_t8 = RG_rl_129 ;
	7'h2c :
		rl_a02_t8 = RG_rl_129 ;
	7'h2d :
		rl_a02_t8 = RG_rl_129 ;
	7'h2e :
		rl_a02_t8 = RG_rl_129 ;
	7'h2f :
		rl_a02_t8 = RG_rl_129 ;
	7'h30 :
		rl_a02_t8 = RG_rl_129 ;
	7'h31 :
		rl_a02_t8 = RG_rl_129 ;
	7'h32 :
		rl_a02_t8 = RG_rl_129 ;
	7'h33 :
		rl_a02_t8 = RG_rl_129 ;
	7'h34 :
		rl_a02_t8 = RG_rl_129 ;
	7'h35 :
		rl_a02_t8 = RG_rl_129 ;
	7'h36 :
		rl_a02_t8 = RG_rl_129 ;
	7'h37 :
		rl_a02_t8 = RG_rl_129 ;
	7'h38 :
		rl_a02_t8 = RG_rl_129 ;
	7'h39 :
		rl_a02_t8 = RG_rl_129 ;
	7'h3a :
		rl_a02_t8 = RG_rl_129 ;
	7'h3b :
		rl_a02_t8 = RG_rl_129 ;
	7'h3c :
		rl_a02_t8 = RG_rl_129 ;
	7'h3d :
		rl_a02_t8 = RG_rl_129 ;
	7'h3e :
		rl_a02_t8 = RG_rl_129 ;
	7'h3f :
		rl_a02_t8 = RG_rl_129 ;
	7'h40 :
		rl_a02_t8 = RG_rl_129 ;
	7'h41 :
		rl_a02_t8 = RG_rl_129 ;
	7'h42 :
		rl_a02_t8 = RG_rl_129 ;
	7'h43 :
		rl_a02_t8 = RG_rl_129 ;
	7'h44 :
		rl_a02_t8 = RG_rl_129 ;
	7'h45 :
		rl_a02_t8 = RG_rl_129 ;
	7'h46 :
		rl_a02_t8 = RG_rl_129 ;
	7'h47 :
		rl_a02_t8 = RG_rl_129 ;
	7'h48 :
		rl_a02_t8 = RG_rl_129 ;
	7'h49 :
		rl_a02_t8 = RG_rl_129 ;
	7'h4a :
		rl_a02_t8 = RG_rl_129 ;
	7'h4b :
		rl_a02_t8 = RG_rl_129 ;
	7'h4c :
		rl_a02_t8 = RG_rl_129 ;
	7'h4d :
		rl_a02_t8 = RG_rl_129 ;
	7'h4e :
		rl_a02_t8 = RG_rl_129 ;
	7'h4f :
		rl_a02_t8 = RG_rl_129 ;
	7'h50 :
		rl_a02_t8 = RG_rl_129 ;
	7'h51 :
		rl_a02_t8 = RG_rl_129 ;
	7'h52 :
		rl_a02_t8 = RG_rl_129 ;
	7'h53 :
		rl_a02_t8 = RG_rl_129 ;
	7'h54 :
		rl_a02_t8 = RG_rl_129 ;
	7'h55 :
		rl_a02_t8 = RG_rl_129 ;
	7'h56 :
		rl_a02_t8 = RG_rl_129 ;
	7'h57 :
		rl_a02_t8 = RG_rl_129 ;
	7'h58 :
		rl_a02_t8 = RG_rl_129 ;
	7'h59 :
		rl_a02_t8 = RG_rl_129 ;
	7'h5a :
		rl_a02_t8 = RG_rl_129 ;
	7'h5b :
		rl_a02_t8 = RG_rl_129 ;
	7'h5c :
		rl_a02_t8 = RG_rl_129 ;
	7'h5d :
		rl_a02_t8 = RG_rl_129 ;
	7'h5e :
		rl_a02_t8 = RG_rl_129 ;
	7'h5f :
		rl_a02_t8 = RG_rl_129 ;
	7'h60 :
		rl_a02_t8 = RG_rl_129 ;
	7'h61 :
		rl_a02_t8 = RG_rl_129 ;
	7'h62 :
		rl_a02_t8 = RG_rl_129 ;
	7'h63 :
		rl_a02_t8 = RG_rl_129 ;
	7'h64 :
		rl_a02_t8 = RG_rl_129 ;
	7'h65 :
		rl_a02_t8 = RG_rl_129 ;
	7'h66 :
		rl_a02_t8 = RG_rl_129 ;
	7'h67 :
		rl_a02_t8 = RG_rl_129 ;
	7'h68 :
		rl_a02_t8 = RG_rl_129 ;
	7'h69 :
		rl_a02_t8 = RG_rl_129 ;
	7'h6a :
		rl_a02_t8 = RG_rl_129 ;
	7'h6b :
		rl_a02_t8 = RG_rl_129 ;
	7'h6c :
		rl_a02_t8 = RG_rl_129 ;
	7'h6d :
		rl_a02_t8 = RG_rl_129 ;
	7'h6e :
		rl_a02_t8 = RG_rl_129 ;
	7'h6f :
		rl_a02_t8 = RG_rl_129 ;
	7'h70 :
		rl_a02_t8 = RG_rl_129 ;
	7'h71 :
		rl_a02_t8 = RG_rl_129 ;
	7'h72 :
		rl_a02_t8 = RG_rl_129 ;
	7'h73 :
		rl_a02_t8 = RG_rl_129 ;
	7'h74 :
		rl_a02_t8 = RG_rl_129 ;
	7'h75 :
		rl_a02_t8 = RG_rl_129 ;
	7'h76 :
		rl_a02_t8 = RG_rl_129 ;
	7'h77 :
		rl_a02_t8 = RG_rl_129 ;
	7'h78 :
		rl_a02_t8 = RG_rl_129 ;
	7'h79 :
		rl_a02_t8 = RG_rl_129 ;
	7'h7a :
		rl_a02_t8 = RG_rl_129 ;
	7'h7b :
		rl_a02_t8 = RG_rl_129 ;
	7'h7c :
		rl_a02_t8 = RG_rl_129 ;
	7'h7d :
		rl_a02_t8 = RG_rl_129 ;
	7'h7e :
		rl_a02_t8 = RG_rl_129 ;
	7'h7f :
		rl_a02_t8 = RG_rl_129 ;
	default :
		rl_a02_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_130 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a03_t8 = RG_rl_130 ;
	7'h01 :
		rl_a03_t8 = RG_rl_130 ;
	7'h02 :
		rl_a03_t8 = RG_rl_130 ;
	7'h03 :
		rl_a03_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h04 :
		rl_a03_t8 = RG_rl_130 ;
	7'h05 :
		rl_a03_t8 = RG_rl_130 ;
	7'h06 :
		rl_a03_t8 = RG_rl_130 ;
	7'h07 :
		rl_a03_t8 = RG_rl_130 ;
	7'h08 :
		rl_a03_t8 = RG_rl_130 ;
	7'h09 :
		rl_a03_t8 = RG_rl_130 ;
	7'h0a :
		rl_a03_t8 = RG_rl_130 ;
	7'h0b :
		rl_a03_t8 = RG_rl_130 ;
	7'h0c :
		rl_a03_t8 = RG_rl_130 ;
	7'h0d :
		rl_a03_t8 = RG_rl_130 ;
	7'h0e :
		rl_a03_t8 = RG_rl_130 ;
	7'h0f :
		rl_a03_t8 = RG_rl_130 ;
	7'h10 :
		rl_a03_t8 = RG_rl_130 ;
	7'h11 :
		rl_a03_t8 = RG_rl_130 ;
	7'h12 :
		rl_a03_t8 = RG_rl_130 ;
	7'h13 :
		rl_a03_t8 = RG_rl_130 ;
	7'h14 :
		rl_a03_t8 = RG_rl_130 ;
	7'h15 :
		rl_a03_t8 = RG_rl_130 ;
	7'h16 :
		rl_a03_t8 = RG_rl_130 ;
	7'h17 :
		rl_a03_t8 = RG_rl_130 ;
	7'h18 :
		rl_a03_t8 = RG_rl_130 ;
	7'h19 :
		rl_a03_t8 = RG_rl_130 ;
	7'h1a :
		rl_a03_t8 = RG_rl_130 ;
	7'h1b :
		rl_a03_t8 = RG_rl_130 ;
	7'h1c :
		rl_a03_t8 = RG_rl_130 ;
	7'h1d :
		rl_a03_t8 = RG_rl_130 ;
	7'h1e :
		rl_a03_t8 = RG_rl_130 ;
	7'h1f :
		rl_a03_t8 = RG_rl_130 ;
	7'h20 :
		rl_a03_t8 = RG_rl_130 ;
	7'h21 :
		rl_a03_t8 = RG_rl_130 ;
	7'h22 :
		rl_a03_t8 = RG_rl_130 ;
	7'h23 :
		rl_a03_t8 = RG_rl_130 ;
	7'h24 :
		rl_a03_t8 = RG_rl_130 ;
	7'h25 :
		rl_a03_t8 = RG_rl_130 ;
	7'h26 :
		rl_a03_t8 = RG_rl_130 ;
	7'h27 :
		rl_a03_t8 = RG_rl_130 ;
	7'h28 :
		rl_a03_t8 = RG_rl_130 ;
	7'h29 :
		rl_a03_t8 = RG_rl_130 ;
	7'h2a :
		rl_a03_t8 = RG_rl_130 ;
	7'h2b :
		rl_a03_t8 = RG_rl_130 ;
	7'h2c :
		rl_a03_t8 = RG_rl_130 ;
	7'h2d :
		rl_a03_t8 = RG_rl_130 ;
	7'h2e :
		rl_a03_t8 = RG_rl_130 ;
	7'h2f :
		rl_a03_t8 = RG_rl_130 ;
	7'h30 :
		rl_a03_t8 = RG_rl_130 ;
	7'h31 :
		rl_a03_t8 = RG_rl_130 ;
	7'h32 :
		rl_a03_t8 = RG_rl_130 ;
	7'h33 :
		rl_a03_t8 = RG_rl_130 ;
	7'h34 :
		rl_a03_t8 = RG_rl_130 ;
	7'h35 :
		rl_a03_t8 = RG_rl_130 ;
	7'h36 :
		rl_a03_t8 = RG_rl_130 ;
	7'h37 :
		rl_a03_t8 = RG_rl_130 ;
	7'h38 :
		rl_a03_t8 = RG_rl_130 ;
	7'h39 :
		rl_a03_t8 = RG_rl_130 ;
	7'h3a :
		rl_a03_t8 = RG_rl_130 ;
	7'h3b :
		rl_a03_t8 = RG_rl_130 ;
	7'h3c :
		rl_a03_t8 = RG_rl_130 ;
	7'h3d :
		rl_a03_t8 = RG_rl_130 ;
	7'h3e :
		rl_a03_t8 = RG_rl_130 ;
	7'h3f :
		rl_a03_t8 = RG_rl_130 ;
	7'h40 :
		rl_a03_t8 = RG_rl_130 ;
	7'h41 :
		rl_a03_t8 = RG_rl_130 ;
	7'h42 :
		rl_a03_t8 = RG_rl_130 ;
	7'h43 :
		rl_a03_t8 = RG_rl_130 ;
	7'h44 :
		rl_a03_t8 = RG_rl_130 ;
	7'h45 :
		rl_a03_t8 = RG_rl_130 ;
	7'h46 :
		rl_a03_t8 = RG_rl_130 ;
	7'h47 :
		rl_a03_t8 = RG_rl_130 ;
	7'h48 :
		rl_a03_t8 = RG_rl_130 ;
	7'h49 :
		rl_a03_t8 = RG_rl_130 ;
	7'h4a :
		rl_a03_t8 = RG_rl_130 ;
	7'h4b :
		rl_a03_t8 = RG_rl_130 ;
	7'h4c :
		rl_a03_t8 = RG_rl_130 ;
	7'h4d :
		rl_a03_t8 = RG_rl_130 ;
	7'h4e :
		rl_a03_t8 = RG_rl_130 ;
	7'h4f :
		rl_a03_t8 = RG_rl_130 ;
	7'h50 :
		rl_a03_t8 = RG_rl_130 ;
	7'h51 :
		rl_a03_t8 = RG_rl_130 ;
	7'h52 :
		rl_a03_t8 = RG_rl_130 ;
	7'h53 :
		rl_a03_t8 = RG_rl_130 ;
	7'h54 :
		rl_a03_t8 = RG_rl_130 ;
	7'h55 :
		rl_a03_t8 = RG_rl_130 ;
	7'h56 :
		rl_a03_t8 = RG_rl_130 ;
	7'h57 :
		rl_a03_t8 = RG_rl_130 ;
	7'h58 :
		rl_a03_t8 = RG_rl_130 ;
	7'h59 :
		rl_a03_t8 = RG_rl_130 ;
	7'h5a :
		rl_a03_t8 = RG_rl_130 ;
	7'h5b :
		rl_a03_t8 = RG_rl_130 ;
	7'h5c :
		rl_a03_t8 = RG_rl_130 ;
	7'h5d :
		rl_a03_t8 = RG_rl_130 ;
	7'h5e :
		rl_a03_t8 = RG_rl_130 ;
	7'h5f :
		rl_a03_t8 = RG_rl_130 ;
	7'h60 :
		rl_a03_t8 = RG_rl_130 ;
	7'h61 :
		rl_a03_t8 = RG_rl_130 ;
	7'h62 :
		rl_a03_t8 = RG_rl_130 ;
	7'h63 :
		rl_a03_t8 = RG_rl_130 ;
	7'h64 :
		rl_a03_t8 = RG_rl_130 ;
	7'h65 :
		rl_a03_t8 = RG_rl_130 ;
	7'h66 :
		rl_a03_t8 = RG_rl_130 ;
	7'h67 :
		rl_a03_t8 = RG_rl_130 ;
	7'h68 :
		rl_a03_t8 = RG_rl_130 ;
	7'h69 :
		rl_a03_t8 = RG_rl_130 ;
	7'h6a :
		rl_a03_t8 = RG_rl_130 ;
	7'h6b :
		rl_a03_t8 = RG_rl_130 ;
	7'h6c :
		rl_a03_t8 = RG_rl_130 ;
	7'h6d :
		rl_a03_t8 = RG_rl_130 ;
	7'h6e :
		rl_a03_t8 = RG_rl_130 ;
	7'h6f :
		rl_a03_t8 = RG_rl_130 ;
	7'h70 :
		rl_a03_t8 = RG_rl_130 ;
	7'h71 :
		rl_a03_t8 = RG_rl_130 ;
	7'h72 :
		rl_a03_t8 = RG_rl_130 ;
	7'h73 :
		rl_a03_t8 = RG_rl_130 ;
	7'h74 :
		rl_a03_t8 = RG_rl_130 ;
	7'h75 :
		rl_a03_t8 = RG_rl_130 ;
	7'h76 :
		rl_a03_t8 = RG_rl_130 ;
	7'h77 :
		rl_a03_t8 = RG_rl_130 ;
	7'h78 :
		rl_a03_t8 = RG_rl_130 ;
	7'h79 :
		rl_a03_t8 = RG_rl_130 ;
	7'h7a :
		rl_a03_t8 = RG_rl_130 ;
	7'h7b :
		rl_a03_t8 = RG_rl_130 ;
	7'h7c :
		rl_a03_t8 = RG_rl_130 ;
	7'h7d :
		rl_a03_t8 = RG_rl_130 ;
	7'h7e :
		rl_a03_t8 = RG_rl_130 ;
	7'h7f :
		rl_a03_t8 = RG_rl_130 ;
	default :
		rl_a03_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_131 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a04_t8 = RG_rl_131 ;
	7'h01 :
		rl_a04_t8 = RG_rl_131 ;
	7'h02 :
		rl_a04_t8 = RG_rl_131 ;
	7'h03 :
		rl_a04_t8 = RG_rl_131 ;
	7'h04 :
		rl_a04_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h05 :
		rl_a04_t8 = RG_rl_131 ;
	7'h06 :
		rl_a04_t8 = RG_rl_131 ;
	7'h07 :
		rl_a04_t8 = RG_rl_131 ;
	7'h08 :
		rl_a04_t8 = RG_rl_131 ;
	7'h09 :
		rl_a04_t8 = RG_rl_131 ;
	7'h0a :
		rl_a04_t8 = RG_rl_131 ;
	7'h0b :
		rl_a04_t8 = RG_rl_131 ;
	7'h0c :
		rl_a04_t8 = RG_rl_131 ;
	7'h0d :
		rl_a04_t8 = RG_rl_131 ;
	7'h0e :
		rl_a04_t8 = RG_rl_131 ;
	7'h0f :
		rl_a04_t8 = RG_rl_131 ;
	7'h10 :
		rl_a04_t8 = RG_rl_131 ;
	7'h11 :
		rl_a04_t8 = RG_rl_131 ;
	7'h12 :
		rl_a04_t8 = RG_rl_131 ;
	7'h13 :
		rl_a04_t8 = RG_rl_131 ;
	7'h14 :
		rl_a04_t8 = RG_rl_131 ;
	7'h15 :
		rl_a04_t8 = RG_rl_131 ;
	7'h16 :
		rl_a04_t8 = RG_rl_131 ;
	7'h17 :
		rl_a04_t8 = RG_rl_131 ;
	7'h18 :
		rl_a04_t8 = RG_rl_131 ;
	7'h19 :
		rl_a04_t8 = RG_rl_131 ;
	7'h1a :
		rl_a04_t8 = RG_rl_131 ;
	7'h1b :
		rl_a04_t8 = RG_rl_131 ;
	7'h1c :
		rl_a04_t8 = RG_rl_131 ;
	7'h1d :
		rl_a04_t8 = RG_rl_131 ;
	7'h1e :
		rl_a04_t8 = RG_rl_131 ;
	7'h1f :
		rl_a04_t8 = RG_rl_131 ;
	7'h20 :
		rl_a04_t8 = RG_rl_131 ;
	7'h21 :
		rl_a04_t8 = RG_rl_131 ;
	7'h22 :
		rl_a04_t8 = RG_rl_131 ;
	7'h23 :
		rl_a04_t8 = RG_rl_131 ;
	7'h24 :
		rl_a04_t8 = RG_rl_131 ;
	7'h25 :
		rl_a04_t8 = RG_rl_131 ;
	7'h26 :
		rl_a04_t8 = RG_rl_131 ;
	7'h27 :
		rl_a04_t8 = RG_rl_131 ;
	7'h28 :
		rl_a04_t8 = RG_rl_131 ;
	7'h29 :
		rl_a04_t8 = RG_rl_131 ;
	7'h2a :
		rl_a04_t8 = RG_rl_131 ;
	7'h2b :
		rl_a04_t8 = RG_rl_131 ;
	7'h2c :
		rl_a04_t8 = RG_rl_131 ;
	7'h2d :
		rl_a04_t8 = RG_rl_131 ;
	7'h2e :
		rl_a04_t8 = RG_rl_131 ;
	7'h2f :
		rl_a04_t8 = RG_rl_131 ;
	7'h30 :
		rl_a04_t8 = RG_rl_131 ;
	7'h31 :
		rl_a04_t8 = RG_rl_131 ;
	7'h32 :
		rl_a04_t8 = RG_rl_131 ;
	7'h33 :
		rl_a04_t8 = RG_rl_131 ;
	7'h34 :
		rl_a04_t8 = RG_rl_131 ;
	7'h35 :
		rl_a04_t8 = RG_rl_131 ;
	7'h36 :
		rl_a04_t8 = RG_rl_131 ;
	7'h37 :
		rl_a04_t8 = RG_rl_131 ;
	7'h38 :
		rl_a04_t8 = RG_rl_131 ;
	7'h39 :
		rl_a04_t8 = RG_rl_131 ;
	7'h3a :
		rl_a04_t8 = RG_rl_131 ;
	7'h3b :
		rl_a04_t8 = RG_rl_131 ;
	7'h3c :
		rl_a04_t8 = RG_rl_131 ;
	7'h3d :
		rl_a04_t8 = RG_rl_131 ;
	7'h3e :
		rl_a04_t8 = RG_rl_131 ;
	7'h3f :
		rl_a04_t8 = RG_rl_131 ;
	7'h40 :
		rl_a04_t8 = RG_rl_131 ;
	7'h41 :
		rl_a04_t8 = RG_rl_131 ;
	7'h42 :
		rl_a04_t8 = RG_rl_131 ;
	7'h43 :
		rl_a04_t8 = RG_rl_131 ;
	7'h44 :
		rl_a04_t8 = RG_rl_131 ;
	7'h45 :
		rl_a04_t8 = RG_rl_131 ;
	7'h46 :
		rl_a04_t8 = RG_rl_131 ;
	7'h47 :
		rl_a04_t8 = RG_rl_131 ;
	7'h48 :
		rl_a04_t8 = RG_rl_131 ;
	7'h49 :
		rl_a04_t8 = RG_rl_131 ;
	7'h4a :
		rl_a04_t8 = RG_rl_131 ;
	7'h4b :
		rl_a04_t8 = RG_rl_131 ;
	7'h4c :
		rl_a04_t8 = RG_rl_131 ;
	7'h4d :
		rl_a04_t8 = RG_rl_131 ;
	7'h4e :
		rl_a04_t8 = RG_rl_131 ;
	7'h4f :
		rl_a04_t8 = RG_rl_131 ;
	7'h50 :
		rl_a04_t8 = RG_rl_131 ;
	7'h51 :
		rl_a04_t8 = RG_rl_131 ;
	7'h52 :
		rl_a04_t8 = RG_rl_131 ;
	7'h53 :
		rl_a04_t8 = RG_rl_131 ;
	7'h54 :
		rl_a04_t8 = RG_rl_131 ;
	7'h55 :
		rl_a04_t8 = RG_rl_131 ;
	7'h56 :
		rl_a04_t8 = RG_rl_131 ;
	7'h57 :
		rl_a04_t8 = RG_rl_131 ;
	7'h58 :
		rl_a04_t8 = RG_rl_131 ;
	7'h59 :
		rl_a04_t8 = RG_rl_131 ;
	7'h5a :
		rl_a04_t8 = RG_rl_131 ;
	7'h5b :
		rl_a04_t8 = RG_rl_131 ;
	7'h5c :
		rl_a04_t8 = RG_rl_131 ;
	7'h5d :
		rl_a04_t8 = RG_rl_131 ;
	7'h5e :
		rl_a04_t8 = RG_rl_131 ;
	7'h5f :
		rl_a04_t8 = RG_rl_131 ;
	7'h60 :
		rl_a04_t8 = RG_rl_131 ;
	7'h61 :
		rl_a04_t8 = RG_rl_131 ;
	7'h62 :
		rl_a04_t8 = RG_rl_131 ;
	7'h63 :
		rl_a04_t8 = RG_rl_131 ;
	7'h64 :
		rl_a04_t8 = RG_rl_131 ;
	7'h65 :
		rl_a04_t8 = RG_rl_131 ;
	7'h66 :
		rl_a04_t8 = RG_rl_131 ;
	7'h67 :
		rl_a04_t8 = RG_rl_131 ;
	7'h68 :
		rl_a04_t8 = RG_rl_131 ;
	7'h69 :
		rl_a04_t8 = RG_rl_131 ;
	7'h6a :
		rl_a04_t8 = RG_rl_131 ;
	7'h6b :
		rl_a04_t8 = RG_rl_131 ;
	7'h6c :
		rl_a04_t8 = RG_rl_131 ;
	7'h6d :
		rl_a04_t8 = RG_rl_131 ;
	7'h6e :
		rl_a04_t8 = RG_rl_131 ;
	7'h6f :
		rl_a04_t8 = RG_rl_131 ;
	7'h70 :
		rl_a04_t8 = RG_rl_131 ;
	7'h71 :
		rl_a04_t8 = RG_rl_131 ;
	7'h72 :
		rl_a04_t8 = RG_rl_131 ;
	7'h73 :
		rl_a04_t8 = RG_rl_131 ;
	7'h74 :
		rl_a04_t8 = RG_rl_131 ;
	7'h75 :
		rl_a04_t8 = RG_rl_131 ;
	7'h76 :
		rl_a04_t8 = RG_rl_131 ;
	7'h77 :
		rl_a04_t8 = RG_rl_131 ;
	7'h78 :
		rl_a04_t8 = RG_rl_131 ;
	7'h79 :
		rl_a04_t8 = RG_rl_131 ;
	7'h7a :
		rl_a04_t8 = RG_rl_131 ;
	7'h7b :
		rl_a04_t8 = RG_rl_131 ;
	7'h7c :
		rl_a04_t8 = RG_rl_131 ;
	7'h7d :
		rl_a04_t8 = RG_rl_131 ;
	7'h7e :
		rl_a04_t8 = RG_rl_131 ;
	7'h7f :
		rl_a04_t8 = RG_rl_131 ;
	default :
		rl_a04_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h01 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h02 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h03 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h04 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h05 :
		rl_a05_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h06 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h07 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h08 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h09 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h0a :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h0b :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h0c :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h0d :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h0e :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h0f :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h10 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h11 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h12 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h13 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h14 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h15 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h16 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h17 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h18 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h19 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h1a :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h1b :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h1c :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h1d :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h1e :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h1f :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h20 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h21 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h22 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h23 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h24 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h25 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h26 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h27 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h28 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h29 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h2a :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h2b :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h2c :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h2d :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h2e :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h2f :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h30 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h31 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h32 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h33 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h34 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h35 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h36 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h37 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h38 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h39 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h3a :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h3b :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h3c :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h3d :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h3e :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h3f :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h40 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h41 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h42 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h43 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h44 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h45 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h46 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h47 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h48 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h49 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h4a :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h4b :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h4c :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h4d :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h4e :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h4f :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h50 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h51 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h52 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h53 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h54 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h55 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h56 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h57 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h58 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h59 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h5a :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h5b :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h5c :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h5d :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h5e :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h5f :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h60 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h61 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h62 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h63 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h64 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h65 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h66 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h67 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h68 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h69 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h6a :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h6b :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h6c :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h6d :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h6e :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h6f :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h70 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h71 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h72 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h73 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h74 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h75 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h76 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h77 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h78 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h79 :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h7a :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h7b :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h7c :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h7d :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h7e :
		rl_a05_t8 = RG_quantized_block_rl ;
	7'h7f :
		rl_a05_t8 = RG_quantized_block_rl ;
	default :
		rl_a05_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_132 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a06_t8 = RG_rl_132 ;
	7'h01 :
		rl_a06_t8 = RG_rl_132 ;
	7'h02 :
		rl_a06_t8 = RG_rl_132 ;
	7'h03 :
		rl_a06_t8 = RG_rl_132 ;
	7'h04 :
		rl_a06_t8 = RG_rl_132 ;
	7'h05 :
		rl_a06_t8 = RG_rl_132 ;
	7'h06 :
		rl_a06_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h07 :
		rl_a06_t8 = RG_rl_132 ;
	7'h08 :
		rl_a06_t8 = RG_rl_132 ;
	7'h09 :
		rl_a06_t8 = RG_rl_132 ;
	7'h0a :
		rl_a06_t8 = RG_rl_132 ;
	7'h0b :
		rl_a06_t8 = RG_rl_132 ;
	7'h0c :
		rl_a06_t8 = RG_rl_132 ;
	7'h0d :
		rl_a06_t8 = RG_rl_132 ;
	7'h0e :
		rl_a06_t8 = RG_rl_132 ;
	7'h0f :
		rl_a06_t8 = RG_rl_132 ;
	7'h10 :
		rl_a06_t8 = RG_rl_132 ;
	7'h11 :
		rl_a06_t8 = RG_rl_132 ;
	7'h12 :
		rl_a06_t8 = RG_rl_132 ;
	7'h13 :
		rl_a06_t8 = RG_rl_132 ;
	7'h14 :
		rl_a06_t8 = RG_rl_132 ;
	7'h15 :
		rl_a06_t8 = RG_rl_132 ;
	7'h16 :
		rl_a06_t8 = RG_rl_132 ;
	7'h17 :
		rl_a06_t8 = RG_rl_132 ;
	7'h18 :
		rl_a06_t8 = RG_rl_132 ;
	7'h19 :
		rl_a06_t8 = RG_rl_132 ;
	7'h1a :
		rl_a06_t8 = RG_rl_132 ;
	7'h1b :
		rl_a06_t8 = RG_rl_132 ;
	7'h1c :
		rl_a06_t8 = RG_rl_132 ;
	7'h1d :
		rl_a06_t8 = RG_rl_132 ;
	7'h1e :
		rl_a06_t8 = RG_rl_132 ;
	7'h1f :
		rl_a06_t8 = RG_rl_132 ;
	7'h20 :
		rl_a06_t8 = RG_rl_132 ;
	7'h21 :
		rl_a06_t8 = RG_rl_132 ;
	7'h22 :
		rl_a06_t8 = RG_rl_132 ;
	7'h23 :
		rl_a06_t8 = RG_rl_132 ;
	7'h24 :
		rl_a06_t8 = RG_rl_132 ;
	7'h25 :
		rl_a06_t8 = RG_rl_132 ;
	7'h26 :
		rl_a06_t8 = RG_rl_132 ;
	7'h27 :
		rl_a06_t8 = RG_rl_132 ;
	7'h28 :
		rl_a06_t8 = RG_rl_132 ;
	7'h29 :
		rl_a06_t8 = RG_rl_132 ;
	7'h2a :
		rl_a06_t8 = RG_rl_132 ;
	7'h2b :
		rl_a06_t8 = RG_rl_132 ;
	7'h2c :
		rl_a06_t8 = RG_rl_132 ;
	7'h2d :
		rl_a06_t8 = RG_rl_132 ;
	7'h2e :
		rl_a06_t8 = RG_rl_132 ;
	7'h2f :
		rl_a06_t8 = RG_rl_132 ;
	7'h30 :
		rl_a06_t8 = RG_rl_132 ;
	7'h31 :
		rl_a06_t8 = RG_rl_132 ;
	7'h32 :
		rl_a06_t8 = RG_rl_132 ;
	7'h33 :
		rl_a06_t8 = RG_rl_132 ;
	7'h34 :
		rl_a06_t8 = RG_rl_132 ;
	7'h35 :
		rl_a06_t8 = RG_rl_132 ;
	7'h36 :
		rl_a06_t8 = RG_rl_132 ;
	7'h37 :
		rl_a06_t8 = RG_rl_132 ;
	7'h38 :
		rl_a06_t8 = RG_rl_132 ;
	7'h39 :
		rl_a06_t8 = RG_rl_132 ;
	7'h3a :
		rl_a06_t8 = RG_rl_132 ;
	7'h3b :
		rl_a06_t8 = RG_rl_132 ;
	7'h3c :
		rl_a06_t8 = RG_rl_132 ;
	7'h3d :
		rl_a06_t8 = RG_rl_132 ;
	7'h3e :
		rl_a06_t8 = RG_rl_132 ;
	7'h3f :
		rl_a06_t8 = RG_rl_132 ;
	7'h40 :
		rl_a06_t8 = RG_rl_132 ;
	7'h41 :
		rl_a06_t8 = RG_rl_132 ;
	7'h42 :
		rl_a06_t8 = RG_rl_132 ;
	7'h43 :
		rl_a06_t8 = RG_rl_132 ;
	7'h44 :
		rl_a06_t8 = RG_rl_132 ;
	7'h45 :
		rl_a06_t8 = RG_rl_132 ;
	7'h46 :
		rl_a06_t8 = RG_rl_132 ;
	7'h47 :
		rl_a06_t8 = RG_rl_132 ;
	7'h48 :
		rl_a06_t8 = RG_rl_132 ;
	7'h49 :
		rl_a06_t8 = RG_rl_132 ;
	7'h4a :
		rl_a06_t8 = RG_rl_132 ;
	7'h4b :
		rl_a06_t8 = RG_rl_132 ;
	7'h4c :
		rl_a06_t8 = RG_rl_132 ;
	7'h4d :
		rl_a06_t8 = RG_rl_132 ;
	7'h4e :
		rl_a06_t8 = RG_rl_132 ;
	7'h4f :
		rl_a06_t8 = RG_rl_132 ;
	7'h50 :
		rl_a06_t8 = RG_rl_132 ;
	7'h51 :
		rl_a06_t8 = RG_rl_132 ;
	7'h52 :
		rl_a06_t8 = RG_rl_132 ;
	7'h53 :
		rl_a06_t8 = RG_rl_132 ;
	7'h54 :
		rl_a06_t8 = RG_rl_132 ;
	7'h55 :
		rl_a06_t8 = RG_rl_132 ;
	7'h56 :
		rl_a06_t8 = RG_rl_132 ;
	7'h57 :
		rl_a06_t8 = RG_rl_132 ;
	7'h58 :
		rl_a06_t8 = RG_rl_132 ;
	7'h59 :
		rl_a06_t8 = RG_rl_132 ;
	7'h5a :
		rl_a06_t8 = RG_rl_132 ;
	7'h5b :
		rl_a06_t8 = RG_rl_132 ;
	7'h5c :
		rl_a06_t8 = RG_rl_132 ;
	7'h5d :
		rl_a06_t8 = RG_rl_132 ;
	7'h5e :
		rl_a06_t8 = RG_rl_132 ;
	7'h5f :
		rl_a06_t8 = RG_rl_132 ;
	7'h60 :
		rl_a06_t8 = RG_rl_132 ;
	7'h61 :
		rl_a06_t8 = RG_rl_132 ;
	7'h62 :
		rl_a06_t8 = RG_rl_132 ;
	7'h63 :
		rl_a06_t8 = RG_rl_132 ;
	7'h64 :
		rl_a06_t8 = RG_rl_132 ;
	7'h65 :
		rl_a06_t8 = RG_rl_132 ;
	7'h66 :
		rl_a06_t8 = RG_rl_132 ;
	7'h67 :
		rl_a06_t8 = RG_rl_132 ;
	7'h68 :
		rl_a06_t8 = RG_rl_132 ;
	7'h69 :
		rl_a06_t8 = RG_rl_132 ;
	7'h6a :
		rl_a06_t8 = RG_rl_132 ;
	7'h6b :
		rl_a06_t8 = RG_rl_132 ;
	7'h6c :
		rl_a06_t8 = RG_rl_132 ;
	7'h6d :
		rl_a06_t8 = RG_rl_132 ;
	7'h6e :
		rl_a06_t8 = RG_rl_132 ;
	7'h6f :
		rl_a06_t8 = RG_rl_132 ;
	7'h70 :
		rl_a06_t8 = RG_rl_132 ;
	7'h71 :
		rl_a06_t8 = RG_rl_132 ;
	7'h72 :
		rl_a06_t8 = RG_rl_132 ;
	7'h73 :
		rl_a06_t8 = RG_rl_132 ;
	7'h74 :
		rl_a06_t8 = RG_rl_132 ;
	7'h75 :
		rl_a06_t8 = RG_rl_132 ;
	7'h76 :
		rl_a06_t8 = RG_rl_132 ;
	7'h77 :
		rl_a06_t8 = RG_rl_132 ;
	7'h78 :
		rl_a06_t8 = RG_rl_132 ;
	7'h79 :
		rl_a06_t8 = RG_rl_132 ;
	7'h7a :
		rl_a06_t8 = RG_rl_132 ;
	7'h7b :
		rl_a06_t8 = RG_rl_132 ;
	7'h7c :
		rl_a06_t8 = RG_rl_132 ;
	7'h7d :
		rl_a06_t8 = RG_rl_132 ;
	7'h7e :
		rl_a06_t8 = RG_rl_132 ;
	7'h7f :
		rl_a06_t8 = RG_rl_132 ;
	default :
		rl_a06_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_1 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h01 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h02 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h03 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h04 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h05 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h06 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h07 :
		rl_a07_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h08 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h09 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h0a :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h0b :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h0c :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h0d :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h0e :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h0f :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h10 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h11 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h12 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h13 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h14 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h15 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h16 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h17 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h18 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h19 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h1a :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h1b :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h1c :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h1d :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h1e :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h1f :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h20 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h21 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h22 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h23 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h24 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h25 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h26 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h27 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h28 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h29 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h2a :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h2b :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h2c :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h2d :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h2e :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h2f :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h30 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h31 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h32 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h33 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h34 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h35 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h36 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h37 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h38 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h39 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h3a :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h3b :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h3c :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h3d :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h3e :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h3f :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h40 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h41 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h42 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h43 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h44 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h45 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h46 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h47 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h48 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h49 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h4a :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h4b :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h4c :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h4d :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h4e :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h4f :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h50 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h51 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h52 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h53 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h54 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h55 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h56 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h57 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h58 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h59 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h5a :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h5b :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h5c :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h5d :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h5e :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h5f :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h60 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h61 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h62 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h63 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h64 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h65 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h66 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h67 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h68 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h69 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h6a :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h6b :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h6c :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h6d :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h6e :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h6f :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h70 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h71 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h72 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h73 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h74 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h75 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h76 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h77 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h78 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h79 :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h7a :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h7b :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h7c :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h7d :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h7e :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	7'h7f :
		rl_a07_t8 = RG_quantized_block_rl_1 ;
	default :
		rl_a07_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_133 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a08_t8 = RG_rl_133 ;
	7'h01 :
		rl_a08_t8 = RG_rl_133 ;
	7'h02 :
		rl_a08_t8 = RG_rl_133 ;
	7'h03 :
		rl_a08_t8 = RG_rl_133 ;
	7'h04 :
		rl_a08_t8 = RG_rl_133 ;
	7'h05 :
		rl_a08_t8 = RG_rl_133 ;
	7'h06 :
		rl_a08_t8 = RG_rl_133 ;
	7'h07 :
		rl_a08_t8 = RG_rl_133 ;
	7'h08 :
		rl_a08_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h09 :
		rl_a08_t8 = RG_rl_133 ;
	7'h0a :
		rl_a08_t8 = RG_rl_133 ;
	7'h0b :
		rl_a08_t8 = RG_rl_133 ;
	7'h0c :
		rl_a08_t8 = RG_rl_133 ;
	7'h0d :
		rl_a08_t8 = RG_rl_133 ;
	7'h0e :
		rl_a08_t8 = RG_rl_133 ;
	7'h0f :
		rl_a08_t8 = RG_rl_133 ;
	7'h10 :
		rl_a08_t8 = RG_rl_133 ;
	7'h11 :
		rl_a08_t8 = RG_rl_133 ;
	7'h12 :
		rl_a08_t8 = RG_rl_133 ;
	7'h13 :
		rl_a08_t8 = RG_rl_133 ;
	7'h14 :
		rl_a08_t8 = RG_rl_133 ;
	7'h15 :
		rl_a08_t8 = RG_rl_133 ;
	7'h16 :
		rl_a08_t8 = RG_rl_133 ;
	7'h17 :
		rl_a08_t8 = RG_rl_133 ;
	7'h18 :
		rl_a08_t8 = RG_rl_133 ;
	7'h19 :
		rl_a08_t8 = RG_rl_133 ;
	7'h1a :
		rl_a08_t8 = RG_rl_133 ;
	7'h1b :
		rl_a08_t8 = RG_rl_133 ;
	7'h1c :
		rl_a08_t8 = RG_rl_133 ;
	7'h1d :
		rl_a08_t8 = RG_rl_133 ;
	7'h1e :
		rl_a08_t8 = RG_rl_133 ;
	7'h1f :
		rl_a08_t8 = RG_rl_133 ;
	7'h20 :
		rl_a08_t8 = RG_rl_133 ;
	7'h21 :
		rl_a08_t8 = RG_rl_133 ;
	7'h22 :
		rl_a08_t8 = RG_rl_133 ;
	7'h23 :
		rl_a08_t8 = RG_rl_133 ;
	7'h24 :
		rl_a08_t8 = RG_rl_133 ;
	7'h25 :
		rl_a08_t8 = RG_rl_133 ;
	7'h26 :
		rl_a08_t8 = RG_rl_133 ;
	7'h27 :
		rl_a08_t8 = RG_rl_133 ;
	7'h28 :
		rl_a08_t8 = RG_rl_133 ;
	7'h29 :
		rl_a08_t8 = RG_rl_133 ;
	7'h2a :
		rl_a08_t8 = RG_rl_133 ;
	7'h2b :
		rl_a08_t8 = RG_rl_133 ;
	7'h2c :
		rl_a08_t8 = RG_rl_133 ;
	7'h2d :
		rl_a08_t8 = RG_rl_133 ;
	7'h2e :
		rl_a08_t8 = RG_rl_133 ;
	7'h2f :
		rl_a08_t8 = RG_rl_133 ;
	7'h30 :
		rl_a08_t8 = RG_rl_133 ;
	7'h31 :
		rl_a08_t8 = RG_rl_133 ;
	7'h32 :
		rl_a08_t8 = RG_rl_133 ;
	7'h33 :
		rl_a08_t8 = RG_rl_133 ;
	7'h34 :
		rl_a08_t8 = RG_rl_133 ;
	7'h35 :
		rl_a08_t8 = RG_rl_133 ;
	7'h36 :
		rl_a08_t8 = RG_rl_133 ;
	7'h37 :
		rl_a08_t8 = RG_rl_133 ;
	7'h38 :
		rl_a08_t8 = RG_rl_133 ;
	7'h39 :
		rl_a08_t8 = RG_rl_133 ;
	7'h3a :
		rl_a08_t8 = RG_rl_133 ;
	7'h3b :
		rl_a08_t8 = RG_rl_133 ;
	7'h3c :
		rl_a08_t8 = RG_rl_133 ;
	7'h3d :
		rl_a08_t8 = RG_rl_133 ;
	7'h3e :
		rl_a08_t8 = RG_rl_133 ;
	7'h3f :
		rl_a08_t8 = RG_rl_133 ;
	7'h40 :
		rl_a08_t8 = RG_rl_133 ;
	7'h41 :
		rl_a08_t8 = RG_rl_133 ;
	7'h42 :
		rl_a08_t8 = RG_rl_133 ;
	7'h43 :
		rl_a08_t8 = RG_rl_133 ;
	7'h44 :
		rl_a08_t8 = RG_rl_133 ;
	7'h45 :
		rl_a08_t8 = RG_rl_133 ;
	7'h46 :
		rl_a08_t8 = RG_rl_133 ;
	7'h47 :
		rl_a08_t8 = RG_rl_133 ;
	7'h48 :
		rl_a08_t8 = RG_rl_133 ;
	7'h49 :
		rl_a08_t8 = RG_rl_133 ;
	7'h4a :
		rl_a08_t8 = RG_rl_133 ;
	7'h4b :
		rl_a08_t8 = RG_rl_133 ;
	7'h4c :
		rl_a08_t8 = RG_rl_133 ;
	7'h4d :
		rl_a08_t8 = RG_rl_133 ;
	7'h4e :
		rl_a08_t8 = RG_rl_133 ;
	7'h4f :
		rl_a08_t8 = RG_rl_133 ;
	7'h50 :
		rl_a08_t8 = RG_rl_133 ;
	7'h51 :
		rl_a08_t8 = RG_rl_133 ;
	7'h52 :
		rl_a08_t8 = RG_rl_133 ;
	7'h53 :
		rl_a08_t8 = RG_rl_133 ;
	7'h54 :
		rl_a08_t8 = RG_rl_133 ;
	7'h55 :
		rl_a08_t8 = RG_rl_133 ;
	7'h56 :
		rl_a08_t8 = RG_rl_133 ;
	7'h57 :
		rl_a08_t8 = RG_rl_133 ;
	7'h58 :
		rl_a08_t8 = RG_rl_133 ;
	7'h59 :
		rl_a08_t8 = RG_rl_133 ;
	7'h5a :
		rl_a08_t8 = RG_rl_133 ;
	7'h5b :
		rl_a08_t8 = RG_rl_133 ;
	7'h5c :
		rl_a08_t8 = RG_rl_133 ;
	7'h5d :
		rl_a08_t8 = RG_rl_133 ;
	7'h5e :
		rl_a08_t8 = RG_rl_133 ;
	7'h5f :
		rl_a08_t8 = RG_rl_133 ;
	7'h60 :
		rl_a08_t8 = RG_rl_133 ;
	7'h61 :
		rl_a08_t8 = RG_rl_133 ;
	7'h62 :
		rl_a08_t8 = RG_rl_133 ;
	7'h63 :
		rl_a08_t8 = RG_rl_133 ;
	7'h64 :
		rl_a08_t8 = RG_rl_133 ;
	7'h65 :
		rl_a08_t8 = RG_rl_133 ;
	7'h66 :
		rl_a08_t8 = RG_rl_133 ;
	7'h67 :
		rl_a08_t8 = RG_rl_133 ;
	7'h68 :
		rl_a08_t8 = RG_rl_133 ;
	7'h69 :
		rl_a08_t8 = RG_rl_133 ;
	7'h6a :
		rl_a08_t8 = RG_rl_133 ;
	7'h6b :
		rl_a08_t8 = RG_rl_133 ;
	7'h6c :
		rl_a08_t8 = RG_rl_133 ;
	7'h6d :
		rl_a08_t8 = RG_rl_133 ;
	7'h6e :
		rl_a08_t8 = RG_rl_133 ;
	7'h6f :
		rl_a08_t8 = RG_rl_133 ;
	7'h70 :
		rl_a08_t8 = RG_rl_133 ;
	7'h71 :
		rl_a08_t8 = RG_rl_133 ;
	7'h72 :
		rl_a08_t8 = RG_rl_133 ;
	7'h73 :
		rl_a08_t8 = RG_rl_133 ;
	7'h74 :
		rl_a08_t8 = RG_rl_133 ;
	7'h75 :
		rl_a08_t8 = RG_rl_133 ;
	7'h76 :
		rl_a08_t8 = RG_rl_133 ;
	7'h77 :
		rl_a08_t8 = RG_rl_133 ;
	7'h78 :
		rl_a08_t8 = RG_rl_133 ;
	7'h79 :
		rl_a08_t8 = RG_rl_133 ;
	7'h7a :
		rl_a08_t8 = RG_rl_133 ;
	7'h7b :
		rl_a08_t8 = RG_rl_133 ;
	7'h7c :
		rl_a08_t8 = RG_rl_133 ;
	7'h7d :
		rl_a08_t8 = RG_rl_133 ;
	7'h7e :
		rl_a08_t8 = RG_rl_133 ;
	7'h7f :
		rl_a08_t8 = RG_rl_133 ;
	default :
		rl_a08_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_2 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h01 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h02 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h03 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h04 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h05 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h06 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h07 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h08 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h09 :
		rl_a09_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h0a :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h0b :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h0c :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h0d :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h0e :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h0f :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h10 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h11 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h12 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h13 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h14 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h15 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h16 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h17 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h18 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h19 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h1a :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h1b :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h1c :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h1d :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h1e :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h1f :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h20 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h21 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h22 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h23 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h24 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h25 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h26 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h27 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h28 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h29 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h2a :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h2b :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h2c :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h2d :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h2e :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h2f :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h30 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h31 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h32 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h33 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h34 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h35 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h36 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h37 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h38 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h39 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h3a :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h3b :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h3c :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h3d :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h3e :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h3f :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h40 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h41 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h42 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h43 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h44 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h45 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h46 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h47 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h48 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h49 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h4a :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h4b :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h4c :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h4d :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h4e :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h4f :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h50 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h51 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h52 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h53 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h54 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h55 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h56 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h57 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h58 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h59 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h5a :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h5b :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h5c :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h5d :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h5e :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h5f :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h60 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h61 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h62 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h63 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h64 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h65 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h66 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h67 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h68 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h69 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h6a :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h6b :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h6c :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h6d :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h6e :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h6f :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h70 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h71 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h72 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h73 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h74 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h75 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h76 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h77 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h78 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h79 :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h7a :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h7b :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h7c :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h7d :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h7e :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	7'h7f :
		rl_a09_t8 = RG_quantized_block_rl_2 ;
	default :
		rl_a09_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_134 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a10_t8 = RG_rl_134 ;
	7'h01 :
		rl_a10_t8 = RG_rl_134 ;
	7'h02 :
		rl_a10_t8 = RG_rl_134 ;
	7'h03 :
		rl_a10_t8 = RG_rl_134 ;
	7'h04 :
		rl_a10_t8 = RG_rl_134 ;
	7'h05 :
		rl_a10_t8 = RG_rl_134 ;
	7'h06 :
		rl_a10_t8 = RG_rl_134 ;
	7'h07 :
		rl_a10_t8 = RG_rl_134 ;
	7'h08 :
		rl_a10_t8 = RG_rl_134 ;
	7'h09 :
		rl_a10_t8 = RG_rl_134 ;
	7'h0a :
		rl_a10_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h0b :
		rl_a10_t8 = RG_rl_134 ;
	7'h0c :
		rl_a10_t8 = RG_rl_134 ;
	7'h0d :
		rl_a10_t8 = RG_rl_134 ;
	7'h0e :
		rl_a10_t8 = RG_rl_134 ;
	7'h0f :
		rl_a10_t8 = RG_rl_134 ;
	7'h10 :
		rl_a10_t8 = RG_rl_134 ;
	7'h11 :
		rl_a10_t8 = RG_rl_134 ;
	7'h12 :
		rl_a10_t8 = RG_rl_134 ;
	7'h13 :
		rl_a10_t8 = RG_rl_134 ;
	7'h14 :
		rl_a10_t8 = RG_rl_134 ;
	7'h15 :
		rl_a10_t8 = RG_rl_134 ;
	7'h16 :
		rl_a10_t8 = RG_rl_134 ;
	7'h17 :
		rl_a10_t8 = RG_rl_134 ;
	7'h18 :
		rl_a10_t8 = RG_rl_134 ;
	7'h19 :
		rl_a10_t8 = RG_rl_134 ;
	7'h1a :
		rl_a10_t8 = RG_rl_134 ;
	7'h1b :
		rl_a10_t8 = RG_rl_134 ;
	7'h1c :
		rl_a10_t8 = RG_rl_134 ;
	7'h1d :
		rl_a10_t8 = RG_rl_134 ;
	7'h1e :
		rl_a10_t8 = RG_rl_134 ;
	7'h1f :
		rl_a10_t8 = RG_rl_134 ;
	7'h20 :
		rl_a10_t8 = RG_rl_134 ;
	7'h21 :
		rl_a10_t8 = RG_rl_134 ;
	7'h22 :
		rl_a10_t8 = RG_rl_134 ;
	7'h23 :
		rl_a10_t8 = RG_rl_134 ;
	7'h24 :
		rl_a10_t8 = RG_rl_134 ;
	7'h25 :
		rl_a10_t8 = RG_rl_134 ;
	7'h26 :
		rl_a10_t8 = RG_rl_134 ;
	7'h27 :
		rl_a10_t8 = RG_rl_134 ;
	7'h28 :
		rl_a10_t8 = RG_rl_134 ;
	7'h29 :
		rl_a10_t8 = RG_rl_134 ;
	7'h2a :
		rl_a10_t8 = RG_rl_134 ;
	7'h2b :
		rl_a10_t8 = RG_rl_134 ;
	7'h2c :
		rl_a10_t8 = RG_rl_134 ;
	7'h2d :
		rl_a10_t8 = RG_rl_134 ;
	7'h2e :
		rl_a10_t8 = RG_rl_134 ;
	7'h2f :
		rl_a10_t8 = RG_rl_134 ;
	7'h30 :
		rl_a10_t8 = RG_rl_134 ;
	7'h31 :
		rl_a10_t8 = RG_rl_134 ;
	7'h32 :
		rl_a10_t8 = RG_rl_134 ;
	7'h33 :
		rl_a10_t8 = RG_rl_134 ;
	7'h34 :
		rl_a10_t8 = RG_rl_134 ;
	7'h35 :
		rl_a10_t8 = RG_rl_134 ;
	7'h36 :
		rl_a10_t8 = RG_rl_134 ;
	7'h37 :
		rl_a10_t8 = RG_rl_134 ;
	7'h38 :
		rl_a10_t8 = RG_rl_134 ;
	7'h39 :
		rl_a10_t8 = RG_rl_134 ;
	7'h3a :
		rl_a10_t8 = RG_rl_134 ;
	7'h3b :
		rl_a10_t8 = RG_rl_134 ;
	7'h3c :
		rl_a10_t8 = RG_rl_134 ;
	7'h3d :
		rl_a10_t8 = RG_rl_134 ;
	7'h3e :
		rl_a10_t8 = RG_rl_134 ;
	7'h3f :
		rl_a10_t8 = RG_rl_134 ;
	7'h40 :
		rl_a10_t8 = RG_rl_134 ;
	7'h41 :
		rl_a10_t8 = RG_rl_134 ;
	7'h42 :
		rl_a10_t8 = RG_rl_134 ;
	7'h43 :
		rl_a10_t8 = RG_rl_134 ;
	7'h44 :
		rl_a10_t8 = RG_rl_134 ;
	7'h45 :
		rl_a10_t8 = RG_rl_134 ;
	7'h46 :
		rl_a10_t8 = RG_rl_134 ;
	7'h47 :
		rl_a10_t8 = RG_rl_134 ;
	7'h48 :
		rl_a10_t8 = RG_rl_134 ;
	7'h49 :
		rl_a10_t8 = RG_rl_134 ;
	7'h4a :
		rl_a10_t8 = RG_rl_134 ;
	7'h4b :
		rl_a10_t8 = RG_rl_134 ;
	7'h4c :
		rl_a10_t8 = RG_rl_134 ;
	7'h4d :
		rl_a10_t8 = RG_rl_134 ;
	7'h4e :
		rl_a10_t8 = RG_rl_134 ;
	7'h4f :
		rl_a10_t8 = RG_rl_134 ;
	7'h50 :
		rl_a10_t8 = RG_rl_134 ;
	7'h51 :
		rl_a10_t8 = RG_rl_134 ;
	7'h52 :
		rl_a10_t8 = RG_rl_134 ;
	7'h53 :
		rl_a10_t8 = RG_rl_134 ;
	7'h54 :
		rl_a10_t8 = RG_rl_134 ;
	7'h55 :
		rl_a10_t8 = RG_rl_134 ;
	7'h56 :
		rl_a10_t8 = RG_rl_134 ;
	7'h57 :
		rl_a10_t8 = RG_rl_134 ;
	7'h58 :
		rl_a10_t8 = RG_rl_134 ;
	7'h59 :
		rl_a10_t8 = RG_rl_134 ;
	7'h5a :
		rl_a10_t8 = RG_rl_134 ;
	7'h5b :
		rl_a10_t8 = RG_rl_134 ;
	7'h5c :
		rl_a10_t8 = RG_rl_134 ;
	7'h5d :
		rl_a10_t8 = RG_rl_134 ;
	7'h5e :
		rl_a10_t8 = RG_rl_134 ;
	7'h5f :
		rl_a10_t8 = RG_rl_134 ;
	7'h60 :
		rl_a10_t8 = RG_rl_134 ;
	7'h61 :
		rl_a10_t8 = RG_rl_134 ;
	7'h62 :
		rl_a10_t8 = RG_rl_134 ;
	7'h63 :
		rl_a10_t8 = RG_rl_134 ;
	7'h64 :
		rl_a10_t8 = RG_rl_134 ;
	7'h65 :
		rl_a10_t8 = RG_rl_134 ;
	7'h66 :
		rl_a10_t8 = RG_rl_134 ;
	7'h67 :
		rl_a10_t8 = RG_rl_134 ;
	7'h68 :
		rl_a10_t8 = RG_rl_134 ;
	7'h69 :
		rl_a10_t8 = RG_rl_134 ;
	7'h6a :
		rl_a10_t8 = RG_rl_134 ;
	7'h6b :
		rl_a10_t8 = RG_rl_134 ;
	7'h6c :
		rl_a10_t8 = RG_rl_134 ;
	7'h6d :
		rl_a10_t8 = RG_rl_134 ;
	7'h6e :
		rl_a10_t8 = RG_rl_134 ;
	7'h6f :
		rl_a10_t8 = RG_rl_134 ;
	7'h70 :
		rl_a10_t8 = RG_rl_134 ;
	7'h71 :
		rl_a10_t8 = RG_rl_134 ;
	7'h72 :
		rl_a10_t8 = RG_rl_134 ;
	7'h73 :
		rl_a10_t8 = RG_rl_134 ;
	7'h74 :
		rl_a10_t8 = RG_rl_134 ;
	7'h75 :
		rl_a10_t8 = RG_rl_134 ;
	7'h76 :
		rl_a10_t8 = RG_rl_134 ;
	7'h77 :
		rl_a10_t8 = RG_rl_134 ;
	7'h78 :
		rl_a10_t8 = RG_rl_134 ;
	7'h79 :
		rl_a10_t8 = RG_rl_134 ;
	7'h7a :
		rl_a10_t8 = RG_rl_134 ;
	7'h7b :
		rl_a10_t8 = RG_rl_134 ;
	7'h7c :
		rl_a10_t8 = RG_rl_134 ;
	7'h7d :
		rl_a10_t8 = RG_rl_134 ;
	7'h7e :
		rl_a10_t8 = RG_rl_134 ;
	7'h7f :
		rl_a10_t8 = RG_rl_134 ;
	default :
		rl_a10_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_3 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h01 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h02 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h03 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h04 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h05 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h06 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h07 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h08 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h09 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h0a :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h0b :
		rl_a11_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h0c :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h0d :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h0e :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h0f :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h10 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h11 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h12 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h13 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h14 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h15 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h16 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h17 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h18 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h19 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h1a :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h1b :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h1c :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h1d :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h1e :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h1f :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h20 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h21 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h22 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h23 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h24 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h25 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h26 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h27 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h28 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h29 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h2a :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h2b :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h2c :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h2d :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h2e :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h2f :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h30 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h31 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h32 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h33 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h34 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h35 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h36 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h37 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h38 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h39 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h3a :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h3b :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h3c :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h3d :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h3e :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h3f :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h40 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h41 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h42 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h43 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h44 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h45 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h46 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h47 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h48 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h49 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h4a :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h4b :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h4c :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h4d :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h4e :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h4f :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h50 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h51 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h52 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h53 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h54 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h55 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h56 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h57 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h58 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h59 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h5a :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h5b :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h5c :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h5d :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h5e :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h5f :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h60 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h61 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h62 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h63 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h64 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h65 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h66 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h67 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h68 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h69 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h6a :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h6b :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h6c :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h6d :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h6e :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h6f :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h70 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h71 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h72 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h73 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h74 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h75 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h76 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h77 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h78 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h79 :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h7a :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h7b :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h7c :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h7d :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h7e :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	7'h7f :
		rl_a11_t8 = RG_quantized_block_rl_3 ;
	default :
		rl_a11_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_135 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a12_t8 = RG_rl_135 ;
	7'h01 :
		rl_a12_t8 = RG_rl_135 ;
	7'h02 :
		rl_a12_t8 = RG_rl_135 ;
	7'h03 :
		rl_a12_t8 = RG_rl_135 ;
	7'h04 :
		rl_a12_t8 = RG_rl_135 ;
	7'h05 :
		rl_a12_t8 = RG_rl_135 ;
	7'h06 :
		rl_a12_t8 = RG_rl_135 ;
	7'h07 :
		rl_a12_t8 = RG_rl_135 ;
	7'h08 :
		rl_a12_t8 = RG_rl_135 ;
	7'h09 :
		rl_a12_t8 = RG_rl_135 ;
	7'h0a :
		rl_a12_t8 = RG_rl_135 ;
	7'h0b :
		rl_a12_t8 = RG_rl_135 ;
	7'h0c :
		rl_a12_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h0d :
		rl_a12_t8 = RG_rl_135 ;
	7'h0e :
		rl_a12_t8 = RG_rl_135 ;
	7'h0f :
		rl_a12_t8 = RG_rl_135 ;
	7'h10 :
		rl_a12_t8 = RG_rl_135 ;
	7'h11 :
		rl_a12_t8 = RG_rl_135 ;
	7'h12 :
		rl_a12_t8 = RG_rl_135 ;
	7'h13 :
		rl_a12_t8 = RG_rl_135 ;
	7'h14 :
		rl_a12_t8 = RG_rl_135 ;
	7'h15 :
		rl_a12_t8 = RG_rl_135 ;
	7'h16 :
		rl_a12_t8 = RG_rl_135 ;
	7'h17 :
		rl_a12_t8 = RG_rl_135 ;
	7'h18 :
		rl_a12_t8 = RG_rl_135 ;
	7'h19 :
		rl_a12_t8 = RG_rl_135 ;
	7'h1a :
		rl_a12_t8 = RG_rl_135 ;
	7'h1b :
		rl_a12_t8 = RG_rl_135 ;
	7'h1c :
		rl_a12_t8 = RG_rl_135 ;
	7'h1d :
		rl_a12_t8 = RG_rl_135 ;
	7'h1e :
		rl_a12_t8 = RG_rl_135 ;
	7'h1f :
		rl_a12_t8 = RG_rl_135 ;
	7'h20 :
		rl_a12_t8 = RG_rl_135 ;
	7'h21 :
		rl_a12_t8 = RG_rl_135 ;
	7'h22 :
		rl_a12_t8 = RG_rl_135 ;
	7'h23 :
		rl_a12_t8 = RG_rl_135 ;
	7'h24 :
		rl_a12_t8 = RG_rl_135 ;
	7'h25 :
		rl_a12_t8 = RG_rl_135 ;
	7'h26 :
		rl_a12_t8 = RG_rl_135 ;
	7'h27 :
		rl_a12_t8 = RG_rl_135 ;
	7'h28 :
		rl_a12_t8 = RG_rl_135 ;
	7'h29 :
		rl_a12_t8 = RG_rl_135 ;
	7'h2a :
		rl_a12_t8 = RG_rl_135 ;
	7'h2b :
		rl_a12_t8 = RG_rl_135 ;
	7'h2c :
		rl_a12_t8 = RG_rl_135 ;
	7'h2d :
		rl_a12_t8 = RG_rl_135 ;
	7'h2e :
		rl_a12_t8 = RG_rl_135 ;
	7'h2f :
		rl_a12_t8 = RG_rl_135 ;
	7'h30 :
		rl_a12_t8 = RG_rl_135 ;
	7'h31 :
		rl_a12_t8 = RG_rl_135 ;
	7'h32 :
		rl_a12_t8 = RG_rl_135 ;
	7'h33 :
		rl_a12_t8 = RG_rl_135 ;
	7'h34 :
		rl_a12_t8 = RG_rl_135 ;
	7'h35 :
		rl_a12_t8 = RG_rl_135 ;
	7'h36 :
		rl_a12_t8 = RG_rl_135 ;
	7'h37 :
		rl_a12_t8 = RG_rl_135 ;
	7'h38 :
		rl_a12_t8 = RG_rl_135 ;
	7'h39 :
		rl_a12_t8 = RG_rl_135 ;
	7'h3a :
		rl_a12_t8 = RG_rl_135 ;
	7'h3b :
		rl_a12_t8 = RG_rl_135 ;
	7'h3c :
		rl_a12_t8 = RG_rl_135 ;
	7'h3d :
		rl_a12_t8 = RG_rl_135 ;
	7'h3e :
		rl_a12_t8 = RG_rl_135 ;
	7'h3f :
		rl_a12_t8 = RG_rl_135 ;
	7'h40 :
		rl_a12_t8 = RG_rl_135 ;
	7'h41 :
		rl_a12_t8 = RG_rl_135 ;
	7'h42 :
		rl_a12_t8 = RG_rl_135 ;
	7'h43 :
		rl_a12_t8 = RG_rl_135 ;
	7'h44 :
		rl_a12_t8 = RG_rl_135 ;
	7'h45 :
		rl_a12_t8 = RG_rl_135 ;
	7'h46 :
		rl_a12_t8 = RG_rl_135 ;
	7'h47 :
		rl_a12_t8 = RG_rl_135 ;
	7'h48 :
		rl_a12_t8 = RG_rl_135 ;
	7'h49 :
		rl_a12_t8 = RG_rl_135 ;
	7'h4a :
		rl_a12_t8 = RG_rl_135 ;
	7'h4b :
		rl_a12_t8 = RG_rl_135 ;
	7'h4c :
		rl_a12_t8 = RG_rl_135 ;
	7'h4d :
		rl_a12_t8 = RG_rl_135 ;
	7'h4e :
		rl_a12_t8 = RG_rl_135 ;
	7'h4f :
		rl_a12_t8 = RG_rl_135 ;
	7'h50 :
		rl_a12_t8 = RG_rl_135 ;
	7'h51 :
		rl_a12_t8 = RG_rl_135 ;
	7'h52 :
		rl_a12_t8 = RG_rl_135 ;
	7'h53 :
		rl_a12_t8 = RG_rl_135 ;
	7'h54 :
		rl_a12_t8 = RG_rl_135 ;
	7'h55 :
		rl_a12_t8 = RG_rl_135 ;
	7'h56 :
		rl_a12_t8 = RG_rl_135 ;
	7'h57 :
		rl_a12_t8 = RG_rl_135 ;
	7'h58 :
		rl_a12_t8 = RG_rl_135 ;
	7'h59 :
		rl_a12_t8 = RG_rl_135 ;
	7'h5a :
		rl_a12_t8 = RG_rl_135 ;
	7'h5b :
		rl_a12_t8 = RG_rl_135 ;
	7'h5c :
		rl_a12_t8 = RG_rl_135 ;
	7'h5d :
		rl_a12_t8 = RG_rl_135 ;
	7'h5e :
		rl_a12_t8 = RG_rl_135 ;
	7'h5f :
		rl_a12_t8 = RG_rl_135 ;
	7'h60 :
		rl_a12_t8 = RG_rl_135 ;
	7'h61 :
		rl_a12_t8 = RG_rl_135 ;
	7'h62 :
		rl_a12_t8 = RG_rl_135 ;
	7'h63 :
		rl_a12_t8 = RG_rl_135 ;
	7'h64 :
		rl_a12_t8 = RG_rl_135 ;
	7'h65 :
		rl_a12_t8 = RG_rl_135 ;
	7'h66 :
		rl_a12_t8 = RG_rl_135 ;
	7'h67 :
		rl_a12_t8 = RG_rl_135 ;
	7'h68 :
		rl_a12_t8 = RG_rl_135 ;
	7'h69 :
		rl_a12_t8 = RG_rl_135 ;
	7'h6a :
		rl_a12_t8 = RG_rl_135 ;
	7'h6b :
		rl_a12_t8 = RG_rl_135 ;
	7'h6c :
		rl_a12_t8 = RG_rl_135 ;
	7'h6d :
		rl_a12_t8 = RG_rl_135 ;
	7'h6e :
		rl_a12_t8 = RG_rl_135 ;
	7'h6f :
		rl_a12_t8 = RG_rl_135 ;
	7'h70 :
		rl_a12_t8 = RG_rl_135 ;
	7'h71 :
		rl_a12_t8 = RG_rl_135 ;
	7'h72 :
		rl_a12_t8 = RG_rl_135 ;
	7'h73 :
		rl_a12_t8 = RG_rl_135 ;
	7'h74 :
		rl_a12_t8 = RG_rl_135 ;
	7'h75 :
		rl_a12_t8 = RG_rl_135 ;
	7'h76 :
		rl_a12_t8 = RG_rl_135 ;
	7'h77 :
		rl_a12_t8 = RG_rl_135 ;
	7'h78 :
		rl_a12_t8 = RG_rl_135 ;
	7'h79 :
		rl_a12_t8 = RG_rl_135 ;
	7'h7a :
		rl_a12_t8 = RG_rl_135 ;
	7'h7b :
		rl_a12_t8 = RG_rl_135 ;
	7'h7c :
		rl_a12_t8 = RG_rl_135 ;
	7'h7d :
		rl_a12_t8 = RG_rl_135 ;
	7'h7e :
		rl_a12_t8 = RG_rl_135 ;
	7'h7f :
		rl_a12_t8 = RG_rl_135 ;
	default :
		rl_a12_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_4 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h01 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h02 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h03 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h04 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h05 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h06 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h07 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h08 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h09 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h0a :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h0b :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h0c :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h0d :
		rl_a13_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h0e :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h0f :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h10 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h11 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h12 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h13 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h14 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h15 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h16 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h17 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h18 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h19 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h1a :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h1b :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h1c :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h1d :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h1e :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h1f :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h20 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h21 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h22 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h23 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h24 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h25 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h26 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h27 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h28 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h29 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h2a :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h2b :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h2c :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h2d :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h2e :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h2f :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h30 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h31 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h32 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h33 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h34 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h35 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h36 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h37 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h38 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h39 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h3a :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h3b :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h3c :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h3d :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h3e :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h3f :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h40 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h41 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h42 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h43 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h44 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h45 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h46 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h47 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h48 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h49 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h4a :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h4b :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h4c :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h4d :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h4e :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h4f :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h50 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h51 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h52 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h53 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h54 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h55 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h56 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h57 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h58 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h59 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h5a :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h5b :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h5c :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h5d :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h5e :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h5f :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h60 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h61 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h62 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h63 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h64 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h65 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h66 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h67 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h68 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h69 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h6a :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h6b :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h6c :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h6d :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h6e :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h6f :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h70 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h71 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h72 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h73 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h74 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h75 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h76 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h77 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h78 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h79 :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h7a :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h7b :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h7c :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h7d :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h7e :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	7'h7f :
		rl_a13_t8 = RG_quantized_block_rl_4 ;
	default :
		rl_a13_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_136 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a14_t8 = RG_rl_136 ;
	7'h01 :
		rl_a14_t8 = RG_rl_136 ;
	7'h02 :
		rl_a14_t8 = RG_rl_136 ;
	7'h03 :
		rl_a14_t8 = RG_rl_136 ;
	7'h04 :
		rl_a14_t8 = RG_rl_136 ;
	7'h05 :
		rl_a14_t8 = RG_rl_136 ;
	7'h06 :
		rl_a14_t8 = RG_rl_136 ;
	7'h07 :
		rl_a14_t8 = RG_rl_136 ;
	7'h08 :
		rl_a14_t8 = RG_rl_136 ;
	7'h09 :
		rl_a14_t8 = RG_rl_136 ;
	7'h0a :
		rl_a14_t8 = RG_rl_136 ;
	7'h0b :
		rl_a14_t8 = RG_rl_136 ;
	7'h0c :
		rl_a14_t8 = RG_rl_136 ;
	7'h0d :
		rl_a14_t8 = RG_rl_136 ;
	7'h0e :
		rl_a14_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h0f :
		rl_a14_t8 = RG_rl_136 ;
	7'h10 :
		rl_a14_t8 = RG_rl_136 ;
	7'h11 :
		rl_a14_t8 = RG_rl_136 ;
	7'h12 :
		rl_a14_t8 = RG_rl_136 ;
	7'h13 :
		rl_a14_t8 = RG_rl_136 ;
	7'h14 :
		rl_a14_t8 = RG_rl_136 ;
	7'h15 :
		rl_a14_t8 = RG_rl_136 ;
	7'h16 :
		rl_a14_t8 = RG_rl_136 ;
	7'h17 :
		rl_a14_t8 = RG_rl_136 ;
	7'h18 :
		rl_a14_t8 = RG_rl_136 ;
	7'h19 :
		rl_a14_t8 = RG_rl_136 ;
	7'h1a :
		rl_a14_t8 = RG_rl_136 ;
	7'h1b :
		rl_a14_t8 = RG_rl_136 ;
	7'h1c :
		rl_a14_t8 = RG_rl_136 ;
	7'h1d :
		rl_a14_t8 = RG_rl_136 ;
	7'h1e :
		rl_a14_t8 = RG_rl_136 ;
	7'h1f :
		rl_a14_t8 = RG_rl_136 ;
	7'h20 :
		rl_a14_t8 = RG_rl_136 ;
	7'h21 :
		rl_a14_t8 = RG_rl_136 ;
	7'h22 :
		rl_a14_t8 = RG_rl_136 ;
	7'h23 :
		rl_a14_t8 = RG_rl_136 ;
	7'h24 :
		rl_a14_t8 = RG_rl_136 ;
	7'h25 :
		rl_a14_t8 = RG_rl_136 ;
	7'h26 :
		rl_a14_t8 = RG_rl_136 ;
	7'h27 :
		rl_a14_t8 = RG_rl_136 ;
	7'h28 :
		rl_a14_t8 = RG_rl_136 ;
	7'h29 :
		rl_a14_t8 = RG_rl_136 ;
	7'h2a :
		rl_a14_t8 = RG_rl_136 ;
	7'h2b :
		rl_a14_t8 = RG_rl_136 ;
	7'h2c :
		rl_a14_t8 = RG_rl_136 ;
	7'h2d :
		rl_a14_t8 = RG_rl_136 ;
	7'h2e :
		rl_a14_t8 = RG_rl_136 ;
	7'h2f :
		rl_a14_t8 = RG_rl_136 ;
	7'h30 :
		rl_a14_t8 = RG_rl_136 ;
	7'h31 :
		rl_a14_t8 = RG_rl_136 ;
	7'h32 :
		rl_a14_t8 = RG_rl_136 ;
	7'h33 :
		rl_a14_t8 = RG_rl_136 ;
	7'h34 :
		rl_a14_t8 = RG_rl_136 ;
	7'h35 :
		rl_a14_t8 = RG_rl_136 ;
	7'h36 :
		rl_a14_t8 = RG_rl_136 ;
	7'h37 :
		rl_a14_t8 = RG_rl_136 ;
	7'h38 :
		rl_a14_t8 = RG_rl_136 ;
	7'h39 :
		rl_a14_t8 = RG_rl_136 ;
	7'h3a :
		rl_a14_t8 = RG_rl_136 ;
	7'h3b :
		rl_a14_t8 = RG_rl_136 ;
	7'h3c :
		rl_a14_t8 = RG_rl_136 ;
	7'h3d :
		rl_a14_t8 = RG_rl_136 ;
	7'h3e :
		rl_a14_t8 = RG_rl_136 ;
	7'h3f :
		rl_a14_t8 = RG_rl_136 ;
	7'h40 :
		rl_a14_t8 = RG_rl_136 ;
	7'h41 :
		rl_a14_t8 = RG_rl_136 ;
	7'h42 :
		rl_a14_t8 = RG_rl_136 ;
	7'h43 :
		rl_a14_t8 = RG_rl_136 ;
	7'h44 :
		rl_a14_t8 = RG_rl_136 ;
	7'h45 :
		rl_a14_t8 = RG_rl_136 ;
	7'h46 :
		rl_a14_t8 = RG_rl_136 ;
	7'h47 :
		rl_a14_t8 = RG_rl_136 ;
	7'h48 :
		rl_a14_t8 = RG_rl_136 ;
	7'h49 :
		rl_a14_t8 = RG_rl_136 ;
	7'h4a :
		rl_a14_t8 = RG_rl_136 ;
	7'h4b :
		rl_a14_t8 = RG_rl_136 ;
	7'h4c :
		rl_a14_t8 = RG_rl_136 ;
	7'h4d :
		rl_a14_t8 = RG_rl_136 ;
	7'h4e :
		rl_a14_t8 = RG_rl_136 ;
	7'h4f :
		rl_a14_t8 = RG_rl_136 ;
	7'h50 :
		rl_a14_t8 = RG_rl_136 ;
	7'h51 :
		rl_a14_t8 = RG_rl_136 ;
	7'h52 :
		rl_a14_t8 = RG_rl_136 ;
	7'h53 :
		rl_a14_t8 = RG_rl_136 ;
	7'h54 :
		rl_a14_t8 = RG_rl_136 ;
	7'h55 :
		rl_a14_t8 = RG_rl_136 ;
	7'h56 :
		rl_a14_t8 = RG_rl_136 ;
	7'h57 :
		rl_a14_t8 = RG_rl_136 ;
	7'h58 :
		rl_a14_t8 = RG_rl_136 ;
	7'h59 :
		rl_a14_t8 = RG_rl_136 ;
	7'h5a :
		rl_a14_t8 = RG_rl_136 ;
	7'h5b :
		rl_a14_t8 = RG_rl_136 ;
	7'h5c :
		rl_a14_t8 = RG_rl_136 ;
	7'h5d :
		rl_a14_t8 = RG_rl_136 ;
	7'h5e :
		rl_a14_t8 = RG_rl_136 ;
	7'h5f :
		rl_a14_t8 = RG_rl_136 ;
	7'h60 :
		rl_a14_t8 = RG_rl_136 ;
	7'h61 :
		rl_a14_t8 = RG_rl_136 ;
	7'h62 :
		rl_a14_t8 = RG_rl_136 ;
	7'h63 :
		rl_a14_t8 = RG_rl_136 ;
	7'h64 :
		rl_a14_t8 = RG_rl_136 ;
	7'h65 :
		rl_a14_t8 = RG_rl_136 ;
	7'h66 :
		rl_a14_t8 = RG_rl_136 ;
	7'h67 :
		rl_a14_t8 = RG_rl_136 ;
	7'h68 :
		rl_a14_t8 = RG_rl_136 ;
	7'h69 :
		rl_a14_t8 = RG_rl_136 ;
	7'h6a :
		rl_a14_t8 = RG_rl_136 ;
	7'h6b :
		rl_a14_t8 = RG_rl_136 ;
	7'h6c :
		rl_a14_t8 = RG_rl_136 ;
	7'h6d :
		rl_a14_t8 = RG_rl_136 ;
	7'h6e :
		rl_a14_t8 = RG_rl_136 ;
	7'h6f :
		rl_a14_t8 = RG_rl_136 ;
	7'h70 :
		rl_a14_t8 = RG_rl_136 ;
	7'h71 :
		rl_a14_t8 = RG_rl_136 ;
	7'h72 :
		rl_a14_t8 = RG_rl_136 ;
	7'h73 :
		rl_a14_t8 = RG_rl_136 ;
	7'h74 :
		rl_a14_t8 = RG_rl_136 ;
	7'h75 :
		rl_a14_t8 = RG_rl_136 ;
	7'h76 :
		rl_a14_t8 = RG_rl_136 ;
	7'h77 :
		rl_a14_t8 = RG_rl_136 ;
	7'h78 :
		rl_a14_t8 = RG_rl_136 ;
	7'h79 :
		rl_a14_t8 = RG_rl_136 ;
	7'h7a :
		rl_a14_t8 = RG_rl_136 ;
	7'h7b :
		rl_a14_t8 = RG_rl_136 ;
	7'h7c :
		rl_a14_t8 = RG_rl_136 ;
	7'h7d :
		rl_a14_t8 = RG_rl_136 ;
	7'h7e :
		rl_a14_t8 = RG_rl_136 ;
	7'h7f :
		rl_a14_t8 = RG_rl_136 ;
	default :
		rl_a14_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_5 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h01 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h02 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h03 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h04 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h05 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h06 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h07 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h08 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h09 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h0a :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h0b :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h0c :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h0d :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h0e :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h0f :
		rl_a15_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h10 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h11 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h12 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h13 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h14 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h15 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h16 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h17 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h18 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h19 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h1a :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h1b :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h1c :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h1d :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h1e :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h1f :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h20 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h21 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h22 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h23 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h24 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h25 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h26 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h27 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h28 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h29 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h2a :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h2b :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h2c :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h2d :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h2e :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h2f :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h30 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h31 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h32 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h33 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h34 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h35 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h36 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h37 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h38 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h39 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h3a :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h3b :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h3c :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h3d :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h3e :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h3f :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h40 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h41 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h42 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h43 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h44 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h45 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h46 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h47 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h48 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h49 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h4a :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h4b :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h4c :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h4d :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h4e :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h4f :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h50 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h51 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h52 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h53 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h54 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h55 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h56 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h57 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h58 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h59 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h5a :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h5b :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h5c :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h5d :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h5e :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h5f :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h60 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h61 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h62 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h63 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h64 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h65 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h66 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h67 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h68 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h69 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h6a :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h6b :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h6c :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h6d :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h6e :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h6f :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h70 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h71 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h72 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h73 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h74 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h75 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h76 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h77 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h78 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h79 :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h7a :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h7b :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h7c :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h7d :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h7e :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	7'h7f :
		rl_a15_t8 = RG_quantized_block_rl_5 ;
	default :
		rl_a15_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_137 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a16_t8 = RG_rl_137 ;
	7'h01 :
		rl_a16_t8 = RG_rl_137 ;
	7'h02 :
		rl_a16_t8 = RG_rl_137 ;
	7'h03 :
		rl_a16_t8 = RG_rl_137 ;
	7'h04 :
		rl_a16_t8 = RG_rl_137 ;
	7'h05 :
		rl_a16_t8 = RG_rl_137 ;
	7'h06 :
		rl_a16_t8 = RG_rl_137 ;
	7'h07 :
		rl_a16_t8 = RG_rl_137 ;
	7'h08 :
		rl_a16_t8 = RG_rl_137 ;
	7'h09 :
		rl_a16_t8 = RG_rl_137 ;
	7'h0a :
		rl_a16_t8 = RG_rl_137 ;
	7'h0b :
		rl_a16_t8 = RG_rl_137 ;
	7'h0c :
		rl_a16_t8 = RG_rl_137 ;
	7'h0d :
		rl_a16_t8 = RG_rl_137 ;
	7'h0e :
		rl_a16_t8 = RG_rl_137 ;
	7'h0f :
		rl_a16_t8 = RG_rl_137 ;
	7'h10 :
		rl_a16_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h11 :
		rl_a16_t8 = RG_rl_137 ;
	7'h12 :
		rl_a16_t8 = RG_rl_137 ;
	7'h13 :
		rl_a16_t8 = RG_rl_137 ;
	7'h14 :
		rl_a16_t8 = RG_rl_137 ;
	7'h15 :
		rl_a16_t8 = RG_rl_137 ;
	7'h16 :
		rl_a16_t8 = RG_rl_137 ;
	7'h17 :
		rl_a16_t8 = RG_rl_137 ;
	7'h18 :
		rl_a16_t8 = RG_rl_137 ;
	7'h19 :
		rl_a16_t8 = RG_rl_137 ;
	7'h1a :
		rl_a16_t8 = RG_rl_137 ;
	7'h1b :
		rl_a16_t8 = RG_rl_137 ;
	7'h1c :
		rl_a16_t8 = RG_rl_137 ;
	7'h1d :
		rl_a16_t8 = RG_rl_137 ;
	7'h1e :
		rl_a16_t8 = RG_rl_137 ;
	7'h1f :
		rl_a16_t8 = RG_rl_137 ;
	7'h20 :
		rl_a16_t8 = RG_rl_137 ;
	7'h21 :
		rl_a16_t8 = RG_rl_137 ;
	7'h22 :
		rl_a16_t8 = RG_rl_137 ;
	7'h23 :
		rl_a16_t8 = RG_rl_137 ;
	7'h24 :
		rl_a16_t8 = RG_rl_137 ;
	7'h25 :
		rl_a16_t8 = RG_rl_137 ;
	7'h26 :
		rl_a16_t8 = RG_rl_137 ;
	7'h27 :
		rl_a16_t8 = RG_rl_137 ;
	7'h28 :
		rl_a16_t8 = RG_rl_137 ;
	7'h29 :
		rl_a16_t8 = RG_rl_137 ;
	7'h2a :
		rl_a16_t8 = RG_rl_137 ;
	7'h2b :
		rl_a16_t8 = RG_rl_137 ;
	7'h2c :
		rl_a16_t8 = RG_rl_137 ;
	7'h2d :
		rl_a16_t8 = RG_rl_137 ;
	7'h2e :
		rl_a16_t8 = RG_rl_137 ;
	7'h2f :
		rl_a16_t8 = RG_rl_137 ;
	7'h30 :
		rl_a16_t8 = RG_rl_137 ;
	7'h31 :
		rl_a16_t8 = RG_rl_137 ;
	7'h32 :
		rl_a16_t8 = RG_rl_137 ;
	7'h33 :
		rl_a16_t8 = RG_rl_137 ;
	7'h34 :
		rl_a16_t8 = RG_rl_137 ;
	7'h35 :
		rl_a16_t8 = RG_rl_137 ;
	7'h36 :
		rl_a16_t8 = RG_rl_137 ;
	7'h37 :
		rl_a16_t8 = RG_rl_137 ;
	7'h38 :
		rl_a16_t8 = RG_rl_137 ;
	7'h39 :
		rl_a16_t8 = RG_rl_137 ;
	7'h3a :
		rl_a16_t8 = RG_rl_137 ;
	7'h3b :
		rl_a16_t8 = RG_rl_137 ;
	7'h3c :
		rl_a16_t8 = RG_rl_137 ;
	7'h3d :
		rl_a16_t8 = RG_rl_137 ;
	7'h3e :
		rl_a16_t8 = RG_rl_137 ;
	7'h3f :
		rl_a16_t8 = RG_rl_137 ;
	7'h40 :
		rl_a16_t8 = RG_rl_137 ;
	7'h41 :
		rl_a16_t8 = RG_rl_137 ;
	7'h42 :
		rl_a16_t8 = RG_rl_137 ;
	7'h43 :
		rl_a16_t8 = RG_rl_137 ;
	7'h44 :
		rl_a16_t8 = RG_rl_137 ;
	7'h45 :
		rl_a16_t8 = RG_rl_137 ;
	7'h46 :
		rl_a16_t8 = RG_rl_137 ;
	7'h47 :
		rl_a16_t8 = RG_rl_137 ;
	7'h48 :
		rl_a16_t8 = RG_rl_137 ;
	7'h49 :
		rl_a16_t8 = RG_rl_137 ;
	7'h4a :
		rl_a16_t8 = RG_rl_137 ;
	7'h4b :
		rl_a16_t8 = RG_rl_137 ;
	7'h4c :
		rl_a16_t8 = RG_rl_137 ;
	7'h4d :
		rl_a16_t8 = RG_rl_137 ;
	7'h4e :
		rl_a16_t8 = RG_rl_137 ;
	7'h4f :
		rl_a16_t8 = RG_rl_137 ;
	7'h50 :
		rl_a16_t8 = RG_rl_137 ;
	7'h51 :
		rl_a16_t8 = RG_rl_137 ;
	7'h52 :
		rl_a16_t8 = RG_rl_137 ;
	7'h53 :
		rl_a16_t8 = RG_rl_137 ;
	7'h54 :
		rl_a16_t8 = RG_rl_137 ;
	7'h55 :
		rl_a16_t8 = RG_rl_137 ;
	7'h56 :
		rl_a16_t8 = RG_rl_137 ;
	7'h57 :
		rl_a16_t8 = RG_rl_137 ;
	7'h58 :
		rl_a16_t8 = RG_rl_137 ;
	7'h59 :
		rl_a16_t8 = RG_rl_137 ;
	7'h5a :
		rl_a16_t8 = RG_rl_137 ;
	7'h5b :
		rl_a16_t8 = RG_rl_137 ;
	7'h5c :
		rl_a16_t8 = RG_rl_137 ;
	7'h5d :
		rl_a16_t8 = RG_rl_137 ;
	7'h5e :
		rl_a16_t8 = RG_rl_137 ;
	7'h5f :
		rl_a16_t8 = RG_rl_137 ;
	7'h60 :
		rl_a16_t8 = RG_rl_137 ;
	7'h61 :
		rl_a16_t8 = RG_rl_137 ;
	7'h62 :
		rl_a16_t8 = RG_rl_137 ;
	7'h63 :
		rl_a16_t8 = RG_rl_137 ;
	7'h64 :
		rl_a16_t8 = RG_rl_137 ;
	7'h65 :
		rl_a16_t8 = RG_rl_137 ;
	7'h66 :
		rl_a16_t8 = RG_rl_137 ;
	7'h67 :
		rl_a16_t8 = RG_rl_137 ;
	7'h68 :
		rl_a16_t8 = RG_rl_137 ;
	7'h69 :
		rl_a16_t8 = RG_rl_137 ;
	7'h6a :
		rl_a16_t8 = RG_rl_137 ;
	7'h6b :
		rl_a16_t8 = RG_rl_137 ;
	7'h6c :
		rl_a16_t8 = RG_rl_137 ;
	7'h6d :
		rl_a16_t8 = RG_rl_137 ;
	7'h6e :
		rl_a16_t8 = RG_rl_137 ;
	7'h6f :
		rl_a16_t8 = RG_rl_137 ;
	7'h70 :
		rl_a16_t8 = RG_rl_137 ;
	7'h71 :
		rl_a16_t8 = RG_rl_137 ;
	7'h72 :
		rl_a16_t8 = RG_rl_137 ;
	7'h73 :
		rl_a16_t8 = RG_rl_137 ;
	7'h74 :
		rl_a16_t8 = RG_rl_137 ;
	7'h75 :
		rl_a16_t8 = RG_rl_137 ;
	7'h76 :
		rl_a16_t8 = RG_rl_137 ;
	7'h77 :
		rl_a16_t8 = RG_rl_137 ;
	7'h78 :
		rl_a16_t8 = RG_rl_137 ;
	7'h79 :
		rl_a16_t8 = RG_rl_137 ;
	7'h7a :
		rl_a16_t8 = RG_rl_137 ;
	7'h7b :
		rl_a16_t8 = RG_rl_137 ;
	7'h7c :
		rl_a16_t8 = RG_rl_137 ;
	7'h7d :
		rl_a16_t8 = RG_rl_137 ;
	7'h7e :
		rl_a16_t8 = RG_rl_137 ;
	7'h7f :
		rl_a16_t8 = RG_rl_137 ;
	default :
		rl_a16_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_6 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h01 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h02 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h03 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h04 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h05 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h06 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h07 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h08 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h09 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h0a :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h0b :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h0c :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h0d :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h0e :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h0f :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h10 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h11 :
		rl_a17_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h12 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h13 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h14 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h15 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h16 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h17 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h18 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h19 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h1a :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h1b :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h1c :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h1d :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h1e :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h1f :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h20 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h21 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h22 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h23 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h24 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h25 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h26 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h27 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h28 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h29 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h2a :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h2b :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h2c :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h2d :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h2e :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h2f :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h30 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h31 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h32 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h33 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h34 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h35 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h36 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h37 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h38 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h39 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h3a :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h3b :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h3c :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h3d :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h3e :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h3f :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h40 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h41 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h42 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h43 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h44 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h45 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h46 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h47 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h48 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h49 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h4a :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h4b :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h4c :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h4d :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h4e :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h4f :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h50 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h51 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h52 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h53 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h54 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h55 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h56 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h57 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h58 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h59 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h5a :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h5b :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h5c :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h5d :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h5e :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h5f :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h60 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h61 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h62 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h63 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h64 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h65 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h66 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h67 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h68 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h69 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h6a :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h6b :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h6c :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h6d :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h6e :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h6f :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h70 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h71 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h72 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h73 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h74 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h75 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h76 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h77 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h78 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h79 :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h7a :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h7b :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h7c :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h7d :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h7e :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	7'h7f :
		rl_a17_t8 = RG_quantized_block_rl_6 ;
	default :
		rl_a17_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_138 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a18_t8 = RG_rl_138 ;
	7'h01 :
		rl_a18_t8 = RG_rl_138 ;
	7'h02 :
		rl_a18_t8 = RG_rl_138 ;
	7'h03 :
		rl_a18_t8 = RG_rl_138 ;
	7'h04 :
		rl_a18_t8 = RG_rl_138 ;
	7'h05 :
		rl_a18_t8 = RG_rl_138 ;
	7'h06 :
		rl_a18_t8 = RG_rl_138 ;
	7'h07 :
		rl_a18_t8 = RG_rl_138 ;
	7'h08 :
		rl_a18_t8 = RG_rl_138 ;
	7'h09 :
		rl_a18_t8 = RG_rl_138 ;
	7'h0a :
		rl_a18_t8 = RG_rl_138 ;
	7'h0b :
		rl_a18_t8 = RG_rl_138 ;
	7'h0c :
		rl_a18_t8 = RG_rl_138 ;
	7'h0d :
		rl_a18_t8 = RG_rl_138 ;
	7'h0e :
		rl_a18_t8 = RG_rl_138 ;
	7'h0f :
		rl_a18_t8 = RG_rl_138 ;
	7'h10 :
		rl_a18_t8 = RG_rl_138 ;
	7'h11 :
		rl_a18_t8 = RG_rl_138 ;
	7'h12 :
		rl_a18_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h13 :
		rl_a18_t8 = RG_rl_138 ;
	7'h14 :
		rl_a18_t8 = RG_rl_138 ;
	7'h15 :
		rl_a18_t8 = RG_rl_138 ;
	7'h16 :
		rl_a18_t8 = RG_rl_138 ;
	7'h17 :
		rl_a18_t8 = RG_rl_138 ;
	7'h18 :
		rl_a18_t8 = RG_rl_138 ;
	7'h19 :
		rl_a18_t8 = RG_rl_138 ;
	7'h1a :
		rl_a18_t8 = RG_rl_138 ;
	7'h1b :
		rl_a18_t8 = RG_rl_138 ;
	7'h1c :
		rl_a18_t8 = RG_rl_138 ;
	7'h1d :
		rl_a18_t8 = RG_rl_138 ;
	7'h1e :
		rl_a18_t8 = RG_rl_138 ;
	7'h1f :
		rl_a18_t8 = RG_rl_138 ;
	7'h20 :
		rl_a18_t8 = RG_rl_138 ;
	7'h21 :
		rl_a18_t8 = RG_rl_138 ;
	7'h22 :
		rl_a18_t8 = RG_rl_138 ;
	7'h23 :
		rl_a18_t8 = RG_rl_138 ;
	7'h24 :
		rl_a18_t8 = RG_rl_138 ;
	7'h25 :
		rl_a18_t8 = RG_rl_138 ;
	7'h26 :
		rl_a18_t8 = RG_rl_138 ;
	7'h27 :
		rl_a18_t8 = RG_rl_138 ;
	7'h28 :
		rl_a18_t8 = RG_rl_138 ;
	7'h29 :
		rl_a18_t8 = RG_rl_138 ;
	7'h2a :
		rl_a18_t8 = RG_rl_138 ;
	7'h2b :
		rl_a18_t8 = RG_rl_138 ;
	7'h2c :
		rl_a18_t8 = RG_rl_138 ;
	7'h2d :
		rl_a18_t8 = RG_rl_138 ;
	7'h2e :
		rl_a18_t8 = RG_rl_138 ;
	7'h2f :
		rl_a18_t8 = RG_rl_138 ;
	7'h30 :
		rl_a18_t8 = RG_rl_138 ;
	7'h31 :
		rl_a18_t8 = RG_rl_138 ;
	7'h32 :
		rl_a18_t8 = RG_rl_138 ;
	7'h33 :
		rl_a18_t8 = RG_rl_138 ;
	7'h34 :
		rl_a18_t8 = RG_rl_138 ;
	7'h35 :
		rl_a18_t8 = RG_rl_138 ;
	7'h36 :
		rl_a18_t8 = RG_rl_138 ;
	7'h37 :
		rl_a18_t8 = RG_rl_138 ;
	7'h38 :
		rl_a18_t8 = RG_rl_138 ;
	7'h39 :
		rl_a18_t8 = RG_rl_138 ;
	7'h3a :
		rl_a18_t8 = RG_rl_138 ;
	7'h3b :
		rl_a18_t8 = RG_rl_138 ;
	7'h3c :
		rl_a18_t8 = RG_rl_138 ;
	7'h3d :
		rl_a18_t8 = RG_rl_138 ;
	7'h3e :
		rl_a18_t8 = RG_rl_138 ;
	7'h3f :
		rl_a18_t8 = RG_rl_138 ;
	7'h40 :
		rl_a18_t8 = RG_rl_138 ;
	7'h41 :
		rl_a18_t8 = RG_rl_138 ;
	7'h42 :
		rl_a18_t8 = RG_rl_138 ;
	7'h43 :
		rl_a18_t8 = RG_rl_138 ;
	7'h44 :
		rl_a18_t8 = RG_rl_138 ;
	7'h45 :
		rl_a18_t8 = RG_rl_138 ;
	7'h46 :
		rl_a18_t8 = RG_rl_138 ;
	7'h47 :
		rl_a18_t8 = RG_rl_138 ;
	7'h48 :
		rl_a18_t8 = RG_rl_138 ;
	7'h49 :
		rl_a18_t8 = RG_rl_138 ;
	7'h4a :
		rl_a18_t8 = RG_rl_138 ;
	7'h4b :
		rl_a18_t8 = RG_rl_138 ;
	7'h4c :
		rl_a18_t8 = RG_rl_138 ;
	7'h4d :
		rl_a18_t8 = RG_rl_138 ;
	7'h4e :
		rl_a18_t8 = RG_rl_138 ;
	7'h4f :
		rl_a18_t8 = RG_rl_138 ;
	7'h50 :
		rl_a18_t8 = RG_rl_138 ;
	7'h51 :
		rl_a18_t8 = RG_rl_138 ;
	7'h52 :
		rl_a18_t8 = RG_rl_138 ;
	7'h53 :
		rl_a18_t8 = RG_rl_138 ;
	7'h54 :
		rl_a18_t8 = RG_rl_138 ;
	7'h55 :
		rl_a18_t8 = RG_rl_138 ;
	7'h56 :
		rl_a18_t8 = RG_rl_138 ;
	7'h57 :
		rl_a18_t8 = RG_rl_138 ;
	7'h58 :
		rl_a18_t8 = RG_rl_138 ;
	7'h59 :
		rl_a18_t8 = RG_rl_138 ;
	7'h5a :
		rl_a18_t8 = RG_rl_138 ;
	7'h5b :
		rl_a18_t8 = RG_rl_138 ;
	7'h5c :
		rl_a18_t8 = RG_rl_138 ;
	7'h5d :
		rl_a18_t8 = RG_rl_138 ;
	7'h5e :
		rl_a18_t8 = RG_rl_138 ;
	7'h5f :
		rl_a18_t8 = RG_rl_138 ;
	7'h60 :
		rl_a18_t8 = RG_rl_138 ;
	7'h61 :
		rl_a18_t8 = RG_rl_138 ;
	7'h62 :
		rl_a18_t8 = RG_rl_138 ;
	7'h63 :
		rl_a18_t8 = RG_rl_138 ;
	7'h64 :
		rl_a18_t8 = RG_rl_138 ;
	7'h65 :
		rl_a18_t8 = RG_rl_138 ;
	7'h66 :
		rl_a18_t8 = RG_rl_138 ;
	7'h67 :
		rl_a18_t8 = RG_rl_138 ;
	7'h68 :
		rl_a18_t8 = RG_rl_138 ;
	7'h69 :
		rl_a18_t8 = RG_rl_138 ;
	7'h6a :
		rl_a18_t8 = RG_rl_138 ;
	7'h6b :
		rl_a18_t8 = RG_rl_138 ;
	7'h6c :
		rl_a18_t8 = RG_rl_138 ;
	7'h6d :
		rl_a18_t8 = RG_rl_138 ;
	7'h6e :
		rl_a18_t8 = RG_rl_138 ;
	7'h6f :
		rl_a18_t8 = RG_rl_138 ;
	7'h70 :
		rl_a18_t8 = RG_rl_138 ;
	7'h71 :
		rl_a18_t8 = RG_rl_138 ;
	7'h72 :
		rl_a18_t8 = RG_rl_138 ;
	7'h73 :
		rl_a18_t8 = RG_rl_138 ;
	7'h74 :
		rl_a18_t8 = RG_rl_138 ;
	7'h75 :
		rl_a18_t8 = RG_rl_138 ;
	7'h76 :
		rl_a18_t8 = RG_rl_138 ;
	7'h77 :
		rl_a18_t8 = RG_rl_138 ;
	7'h78 :
		rl_a18_t8 = RG_rl_138 ;
	7'h79 :
		rl_a18_t8 = RG_rl_138 ;
	7'h7a :
		rl_a18_t8 = RG_rl_138 ;
	7'h7b :
		rl_a18_t8 = RG_rl_138 ;
	7'h7c :
		rl_a18_t8 = RG_rl_138 ;
	7'h7d :
		rl_a18_t8 = RG_rl_138 ;
	7'h7e :
		rl_a18_t8 = RG_rl_138 ;
	7'h7f :
		rl_a18_t8 = RG_rl_138 ;
	default :
		rl_a18_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_7 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h01 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h02 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h03 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h04 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h05 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h06 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h07 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h08 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h09 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h0a :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h0b :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h0c :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h0d :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h0e :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h0f :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h10 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h11 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h12 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h13 :
		rl_a19_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h14 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h15 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h16 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h17 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h18 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h19 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h1a :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h1b :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h1c :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h1d :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h1e :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h1f :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h20 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h21 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h22 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h23 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h24 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h25 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h26 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h27 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h28 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h29 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h2a :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h2b :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h2c :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h2d :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h2e :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h2f :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h30 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h31 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h32 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h33 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h34 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h35 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h36 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h37 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h38 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h39 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h3a :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h3b :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h3c :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h3d :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h3e :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h3f :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h40 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h41 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h42 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h43 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h44 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h45 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h46 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h47 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h48 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h49 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h4a :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h4b :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h4c :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h4d :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h4e :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h4f :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h50 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h51 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h52 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h53 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h54 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h55 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h56 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h57 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h58 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h59 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h5a :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h5b :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h5c :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h5d :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h5e :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h5f :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h60 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h61 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h62 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h63 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h64 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h65 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h66 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h67 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h68 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h69 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h6a :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h6b :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h6c :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h6d :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h6e :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h6f :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h70 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h71 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h72 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h73 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h74 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h75 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h76 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h77 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h78 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h79 :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h7a :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h7b :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h7c :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h7d :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h7e :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	7'h7f :
		rl_a19_t8 = RG_quantized_block_rl_7 ;
	default :
		rl_a19_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_139 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a20_t8 = RG_rl_139 ;
	7'h01 :
		rl_a20_t8 = RG_rl_139 ;
	7'h02 :
		rl_a20_t8 = RG_rl_139 ;
	7'h03 :
		rl_a20_t8 = RG_rl_139 ;
	7'h04 :
		rl_a20_t8 = RG_rl_139 ;
	7'h05 :
		rl_a20_t8 = RG_rl_139 ;
	7'h06 :
		rl_a20_t8 = RG_rl_139 ;
	7'h07 :
		rl_a20_t8 = RG_rl_139 ;
	7'h08 :
		rl_a20_t8 = RG_rl_139 ;
	7'h09 :
		rl_a20_t8 = RG_rl_139 ;
	7'h0a :
		rl_a20_t8 = RG_rl_139 ;
	7'h0b :
		rl_a20_t8 = RG_rl_139 ;
	7'h0c :
		rl_a20_t8 = RG_rl_139 ;
	7'h0d :
		rl_a20_t8 = RG_rl_139 ;
	7'h0e :
		rl_a20_t8 = RG_rl_139 ;
	7'h0f :
		rl_a20_t8 = RG_rl_139 ;
	7'h10 :
		rl_a20_t8 = RG_rl_139 ;
	7'h11 :
		rl_a20_t8 = RG_rl_139 ;
	7'h12 :
		rl_a20_t8 = RG_rl_139 ;
	7'h13 :
		rl_a20_t8 = RG_rl_139 ;
	7'h14 :
		rl_a20_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h15 :
		rl_a20_t8 = RG_rl_139 ;
	7'h16 :
		rl_a20_t8 = RG_rl_139 ;
	7'h17 :
		rl_a20_t8 = RG_rl_139 ;
	7'h18 :
		rl_a20_t8 = RG_rl_139 ;
	7'h19 :
		rl_a20_t8 = RG_rl_139 ;
	7'h1a :
		rl_a20_t8 = RG_rl_139 ;
	7'h1b :
		rl_a20_t8 = RG_rl_139 ;
	7'h1c :
		rl_a20_t8 = RG_rl_139 ;
	7'h1d :
		rl_a20_t8 = RG_rl_139 ;
	7'h1e :
		rl_a20_t8 = RG_rl_139 ;
	7'h1f :
		rl_a20_t8 = RG_rl_139 ;
	7'h20 :
		rl_a20_t8 = RG_rl_139 ;
	7'h21 :
		rl_a20_t8 = RG_rl_139 ;
	7'h22 :
		rl_a20_t8 = RG_rl_139 ;
	7'h23 :
		rl_a20_t8 = RG_rl_139 ;
	7'h24 :
		rl_a20_t8 = RG_rl_139 ;
	7'h25 :
		rl_a20_t8 = RG_rl_139 ;
	7'h26 :
		rl_a20_t8 = RG_rl_139 ;
	7'h27 :
		rl_a20_t8 = RG_rl_139 ;
	7'h28 :
		rl_a20_t8 = RG_rl_139 ;
	7'h29 :
		rl_a20_t8 = RG_rl_139 ;
	7'h2a :
		rl_a20_t8 = RG_rl_139 ;
	7'h2b :
		rl_a20_t8 = RG_rl_139 ;
	7'h2c :
		rl_a20_t8 = RG_rl_139 ;
	7'h2d :
		rl_a20_t8 = RG_rl_139 ;
	7'h2e :
		rl_a20_t8 = RG_rl_139 ;
	7'h2f :
		rl_a20_t8 = RG_rl_139 ;
	7'h30 :
		rl_a20_t8 = RG_rl_139 ;
	7'h31 :
		rl_a20_t8 = RG_rl_139 ;
	7'h32 :
		rl_a20_t8 = RG_rl_139 ;
	7'h33 :
		rl_a20_t8 = RG_rl_139 ;
	7'h34 :
		rl_a20_t8 = RG_rl_139 ;
	7'h35 :
		rl_a20_t8 = RG_rl_139 ;
	7'h36 :
		rl_a20_t8 = RG_rl_139 ;
	7'h37 :
		rl_a20_t8 = RG_rl_139 ;
	7'h38 :
		rl_a20_t8 = RG_rl_139 ;
	7'h39 :
		rl_a20_t8 = RG_rl_139 ;
	7'h3a :
		rl_a20_t8 = RG_rl_139 ;
	7'h3b :
		rl_a20_t8 = RG_rl_139 ;
	7'h3c :
		rl_a20_t8 = RG_rl_139 ;
	7'h3d :
		rl_a20_t8 = RG_rl_139 ;
	7'h3e :
		rl_a20_t8 = RG_rl_139 ;
	7'h3f :
		rl_a20_t8 = RG_rl_139 ;
	7'h40 :
		rl_a20_t8 = RG_rl_139 ;
	7'h41 :
		rl_a20_t8 = RG_rl_139 ;
	7'h42 :
		rl_a20_t8 = RG_rl_139 ;
	7'h43 :
		rl_a20_t8 = RG_rl_139 ;
	7'h44 :
		rl_a20_t8 = RG_rl_139 ;
	7'h45 :
		rl_a20_t8 = RG_rl_139 ;
	7'h46 :
		rl_a20_t8 = RG_rl_139 ;
	7'h47 :
		rl_a20_t8 = RG_rl_139 ;
	7'h48 :
		rl_a20_t8 = RG_rl_139 ;
	7'h49 :
		rl_a20_t8 = RG_rl_139 ;
	7'h4a :
		rl_a20_t8 = RG_rl_139 ;
	7'h4b :
		rl_a20_t8 = RG_rl_139 ;
	7'h4c :
		rl_a20_t8 = RG_rl_139 ;
	7'h4d :
		rl_a20_t8 = RG_rl_139 ;
	7'h4e :
		rl_a20_t8 = RG_rl_139 ;
	7'h4f :
		rl_a20_t8 = RG_rl_139 ;
	7'h50 :
		rl_a20_t8 = RG_rl_139 ;
	7'h51 :
		rl_a20_t8 = RG_rl_139 ;
	7'h52 :
		rl_a20_t8 = RG_rl_139 ;
	7'h53 :
		rl_a20_t8 = RG_rl_139 ;
	7'h54 :
		rl_a20_t8 = RG_rl_139 ;
	7'h55 :
		rl_a20_t8 = RG_rl_139 ;
	7'h56 :
		rl_a20_t8 = RG_rl_139 ;
	7'h57 :
		rl_a20_t8 = RG_rl_139 ;
	7'h58 :
		rl_a20_t8 = RG_rl_139 ;
	7'h59 :
		rl_a20_t8 = RG_rl_139 ;
	7'h5a :
		rl_a20_t8 = RG_rl_139 ;
	7'h5b :
		rl_a20_t8 = RG_rl_139 ;
	7'h5c :
		rl_a20_t8 = RG_rl_139 ;
	7'h5d :
		rl_a20_t8 = RG_rl_139 ;
	7'h5e :
		rl_a20_t8 = RG_rl_139 ;
	7'h5f :
		rl_a20_t8 = RG_rl_139 ;
	7'h60 :
		rl_a20_t8 = RG_rl_139 ;
	7'h61 :
		rl_a20_t8 = RG_rl_139 ;
	7'h62 :
		rl_a20_t8 = RG_rl_139 ;
	7'h63 :
		rl_a20_t8 = RG_rl_139 ;
	7'h64 :
		rl_a20_t8 = RG_rl_139 ;
	7'h65 :
		rl_a20_t8 = RG_rl_139 ;
	7'h66 :
		rl_a20_t8 = RG_rl_139 ;
	7'h67 :
		rl_a20_t8 = RG_rl_139 ;
	7'h68 :
		rl_a20_t8 = RG_rl_139 ;
	7'h69 :
		rl_a20_t8 = RG_rl_139 ;
	7'h6a :
		rl_a20_t8 = RG_rl_139 ;
	7'h6b :
		rl_a20_t8 = RG_rl_139 ;
	7'h6c :
		rl_a20_t8 = RG_rl_139 ;
	7'h6d :
		rl_a20_t8 = RG_rl_139 ;
	7'h6e :
		rl_a20_t8 = RG_rl_139 ;
	7'h6f :
		rl_a20_t8 = RG_rl_139 ;
	7'h70 :
		rl_a20_t8 = RG_rl_139 ;
	7'h71 :
		rl_a20_t8 = RG_rl_139 ;
	7'h72 :
		rl_a20_t8 = RG_rl_139 ;
	7'h73 :
		rl_a20_t8 = RG_rl_139 ;
	7'h74 :
		rl_a20_t8 = RG_rl_139 ;
	7'h75 :
		rl_a20_t8 = RG_rl_139 ;
	7'h76 :
		rl_a20_t8 = RG_rl_139 ;
	7'h77 :
		rl_a20_t8 = RG_rl_139 ;
	7'h78 :
		rl_a20_t8 = RG_rl_139 ;
	7'h79 :
		rl_a20_t8 = RG_rl_139 ;
	7'h7a :
		rl_a20_t8 = RG_rl_139 ;
	7'h7b :
		rl_a20_t8 = RG_rl_139 ;
	7'h7c :
		rl_a20_t8 = RG_rl_139 ;
	7'h7d :
		rl_a20_t8 = RG_rl_139 ;
	7'h7e :
		rl_a20_t8 = RG_rl_139 ;
	7'h7f :
		rl_a20_t8 = RG_rl_139 ;
	default :
		rl_a20_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_8 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h01 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h02 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h03 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h04 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h05 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h06 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h07 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h08 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h09 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h0a :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h0b :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h0c :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h0d :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h0e :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h0f :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h10 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h11 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h12 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h13 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h14 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h15 :
		rl_a21_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h16 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h17 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h18 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h19 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h1a :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h1b :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h1c :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h1d :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h1e :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h1f :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h20 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h21 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h22 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h23 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h24 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h25 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h26 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h27 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h28 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h29 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h2a :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h2b :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h2c :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h2d :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h2e :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h2f :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h30 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h31 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h32 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h33 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h34 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h35 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h36 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h37 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h38 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h39 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h3a :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h3b :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h3c :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h3d :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h3e :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h3f :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h40 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h41 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h42 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h43 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h44 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h45 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h46 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h47 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h48 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h49 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h4a :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h4b :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h4c :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h4d :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h4e :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h4f :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h50 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h51 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h52 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h53 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h54 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h55 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h56 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h57 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h58 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h59 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h5a :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h5b :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h5c :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h5d :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h5e :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h5f :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h60 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h61 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h62 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h63 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h64 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h65 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h66 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h67 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h68 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h69 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h6a :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h6b :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h6c :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h6d :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h6e :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h6f :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h70 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h71 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h72 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h73 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h74 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h75 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h76 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h77 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h78 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h79 :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h7a :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h7b :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h7c :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h7d :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h7e :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	7'h7f :
		rl_a21_t8 = RG_quantized_block_rl_8 ;
	default :
		rl_a21_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_140 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a22_t8 = RG_rl_140 ;
	7'h01 :
		rl_a22_t8 = RG_rl_140 ;
	7'h02 :
		rl_a22_t8 = RG_rl_140 ;
	7'h03 :
		rl_a22_t8 = RG_rl_140 ;
	7'h04 :
		rl_a22_t8 = RG_rl_140 ;
	7'h05 :
		rl_a22_t8 = RG_rl_140 ;
	7'h06 :
		rl_a22_t8 = RG_rl_140 ;
	7'h07 :
		rl_a22_t8 = RG_rl_140 ;
	7'h08 :
		rl_a22_t8 = RG_rl_140 ;
	7'h09 :
		rl_a22_t8 = RG_rl_140 ;
	7'h0a :
		rl_a22_t8 = RG_rl_140 ;
	7'h0b :
		rl_a22_t8 = RG_rl_140 ;
	7'h0c :
		rl_a22_t8 = RG_rl_140 ;
	7'h0d :
		rl_a22_t8 = RG_rl_140 ;
	7'h0e :
		rl_a22_t8 = RG_rl_140 ;
	7'h0f :
		rl_a22_t8 = RG_rl_140 ;
	7'h10 :
		rl_a22_t8 = RG_rl_140 ;
	7'h11 :
		rl_a22_t8 = RG_rl_140 ;
	7'h12 :
		rl_a22_t8 = RG_rl_140 ;
	7'h13 :
		rl_a22_t8 = RG_rl_140 ;
	7'h14 :
		rl_a22_t8 = RG_rl_140 ;
	7'h15 :
		rl_a22_t8 = RG_rl_140 ;
	7'h16 :
		rl_a22_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h17 :
		rl_a22_t8 = RG_rl_140 ;
	7'h18 :
		rl_a22_t8 = RG_rl_140 ;
	7'h19 :
		rl_a22_t8 = RG_rl_140 ;
	7'h1a :
		rl_a22_t8 = RG_rl_140 ;
	7'h1b :
		rl_a22_t8 = RG_rl_140 ;
	7'h1c :
		rl_a22_t8 = RG_rl_140 ;
	7'h1d :
		rl_a22_t8 = RG_rl_140 ;
	7'h1e :
		rl_a22_t8 = RG_rl_140 ;
	7'h1f :
		rl_a22_t8 = RG_rl_140 ;
	7'h20 :
		rl_a22_t8 = RG_rl_140 ;
	7'h21 :
		rl_a22_t8 = RG_rl_140 ;
	7'h22 :
		rl_a22_t8 = RG_rl_140 ;
	7'h23 :
		rl_a22_t8 = RG_rl_140 ;
	7'h24 :
		rl_a22_t8 = RG_rl_140 ;
	7'h25 :
		rl_a22_t8 = RG_rl_140 ;
	7'h26 :
		rl_a22_t8 = RG_rl_140 ;
	7'h27 :
		rl_a22_t8 = RG_rl_140 ;
	7'h28 :
		rl_a22_t8 = RG_rl_140 ;
	7'h29 :
		rl_a22_t8 = RG_rl_140 ;
	7'h2a :
		rl_a22_t8 = RG_rl_140 ;
	7'h2b :
		rl_a22_t8 = RG_rl_140 ;
	7'h2c :
		rl_a22_t8 = RG_rl_140 ;
	7'h2d :
		rl_a22_t8 = RG_rl_140 ;
	7'h2e :
		rl_a22_t8 = RG_rl_140 ;
	7'h2f :
		rl_a22_t8 = RG_rl_140 ;
	7'h30 :
		rl_a22_t8 = RG_rl_140 ;
	7'h31 :
		rl_a22_t8 = RG_rl_140 ;
	7'h32 :
		rl_a22_t8 = RG_rl_140 ;
	7'h33 :
		rl_a22_t8 = RG_rl_140 ;
	7'h34 :
		rl_a22_t8 = RG_rl_140 ;
	7'h35 :
		rl_a22_t8 = RG_rl_140 ;
	7'h36 :
		rl_a22_t8 = RG_rl_140 ;
	7'h37 :
		rl_a22_t8 = RG_rl_140 ;
	7'h38 :
		rl_a22_t8 = RG_rl_140 ;
	7'h39 :
		rl_a22_t8 = RG_rl_140 ;
	7'h3a :
		rl_a22_t8 = RG_rl_140 ;
	7'h3b :
		rl_a22_t8 = RG_rl_140 ;
	7'h3c :
		rl_a22_t8 = RG_rl_140 ;
	7'h3d :
		rl_a22_t8 = RG_rl_140 ;
	7'h3e :
		rl_a22_t8 = RG_rl_140 ;
	7'h3f :
		rl_a22_t8 = RG_rl_140 ;
	7'h40 :
		rl_a22_t8 = RG_rl_140 ;
	7'h41 :
		rl_a22_t8 = RG_rl_140 ;
	7'h42 :
		rl_a22_t8 = RG_rl_140 ;
	7'h43 :
		rl_a22_t8 = RG_rl_140 ;
	7'h44 :
		rl_a22_t8 = RG_rl_140 ;
	7'h45 :
		rl_a22_t8 = RG_rl_140 ;
	7'h46 :
		rl_a22_t8 = RG_rl_140 ;
	7'h47 :
		rl_a22_t8 = RG_rl_140 ;
	7'h48 :
		rl_a22_t8 = RG_rl_140 ;
	7'h49 :
		rl_a22_t8 = RG_rl_140 ;
	7'h4a :
		rl_a22_t8 = RG_rl_140 ;
	7'h4b :
		rl_a22_t8 = RG_rl_140 ;
	7'h4c :
		rl_a22_t8 = RG_rl_140 ;
	7'h4d :
		rl_a22_t8 = RG_rl_140 ;
	7'h4e :
		rl_a22_t8 = RG_rl_140 ;
	7'h4f :
		rl_a22_t8 = RG_rl_140 ;
	7'h50 :
		rl_a22_t8 = RG_rl_140 ;
	7'h51 :
		rl_a22_t8 = RG_rl_140 ;
	7'h52 :
		rl_a22_t8 = RG_rl_140 ;
	7'h53 :
		rl_a22_t8 = RG_rl_140 ;
	7'h54 :
		rl_a22_t8 = RG_rl_140 ;
	7'h55 :
		rl_a22_t8 = RG_rl_140 ;
	7'h56 :
		rl_a22_t8 = RG_rl_140 ;
	7'h57 :
		rl_a22_t8 = RG_rl_140 ;
	7'h58 :
		rl_a22_t8 = RG_rl_140 ;
	7'h59 :
		rl_a22_t8 = RG_rl_140 ;
	7'h5a :
		rl_a22_t8 = RG_rl_140 ;
	7'h5b :
		rl_a22_t8 = RG_rl_140 ;
	7'h5c :
		rl_a22_t8 = RG_rl_140 ;
	7'h5d :
		rl_a22_t8 = RG_rl_140 ;
	7'h5e :
		rl_a22_t8 = RG_rl_140 ;
	7'h5f :
		rl_a22_t8 = RG_rl_140 ;
	7'h60 :
		rl_a22_t8 = RG_rl_140 ;
	7'h61 :
		rl_a22_t8 = RG_rl_140 ;
	7'h62 :
		rl_a22_t8 = RG_rl_140 ;
	7'h63 :
		rl_a22_t8 = RG_rl_140 ;
	7'h64 :
		rl_a22_t8 = RG_rl_140 ;
	7'h65 :
		rl_a22_t8 = RG_rl_140 ;
	7'h66 :
		rl_a22_t8 = RG_rl_140 ;
	7'h67 :
		rl_a22_t8 = RG_rl_140 ;
	7'h68 :
		rl_a22_t8 = RG_rl_140 ;
	7'h69 :
		rl_a22_t8 = RG_rl_140 ;
	7'h6a :
		rl_a22_t8 = RG_rl_140 ;
	7'h6b :
		rl_a22_t8 = RG_rl_140 ;
	7'h6c :
		rl_a22_t8 = RG_rl_140 ;
	7'h6d :
		rl_a22_t8 = RG_rl_140 ;
	7'h6e :
		rl_a22_t8 = RG_rl_140 ;
	7'h6f :
		rl_a22_t8 = RG_rl_140 ;
	7'h70 :
		rl_a22_t8 = RG_rl_140 ;
	7'h71 :
		rl_a22_t8 = RG_rl_140 ;
	7'h72 :
		rl_a22_t8 = RG_rl_140 ;
	7'h73 :
		rl_a22_t8 = RG_rl_140 ;
	7'h74 :
		rl_a22_t8 = RG_rl_140 ;
	7'h75 :
		rl_a22_t8 = RG_rl_140 ;
	7'h76 :
		rl_a22_t8 = RG_rl_140 ;
	7'h77 :
		rl_a22_t8 = RG_rl_140 ;
	7'h78 :
		rl_a22_t8 = RG_rl_140 ;
	7'h79 :
		rl_a22_t8 = RG_rl_140 ;
	7'h7a :
		rl_a22_t8 = RG_rl_140 ;
	7'h7b :
		rl_a22_t8 = RG_rl_140 ;
	7'h7c :
		rl_a22_t8 = RG_rl_140 ;
	7'h7d :
		rl_a22_t8 = RG_rl_140 ;
	7'h7e :
		rl_a22_t8 = RG_rl_140 ;
	7'h7f :
		rl_a22_t8 = RG_rl_140 ;
	default :
		rl_a22_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_9 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h01 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h02 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h03 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h04 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h05 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h06 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h07 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h08 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h09 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h0a :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h0b :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h0c :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h0d :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h0e :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h0f :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h10 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h11 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h12 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h13 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h14 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h15 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h16 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h17 :
		rl_a23_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h18 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h19 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h1a :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h1b :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h1c :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h1d :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h1e :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h1f :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h20 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h21 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h22 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h23 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h24 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h25 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h26 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h27 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h28 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h29 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h2a :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h2b :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h2c :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h2d :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h2e :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h2f :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h30 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h31 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h32 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h33 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h34 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h35 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h36 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h37 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h38 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h39 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h3a :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h3b :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h3c :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h3d :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h3e :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h3f :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h40 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h41 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h42 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h43 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h44 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h45 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h46 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h47 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h48 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h49 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h4a :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h4b :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h4c :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h4d :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h4e :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h4f :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h50 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h51 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h52 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h53 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h54 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h55 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h56 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h57 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h58 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h59 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h5a :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h5b :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h5c :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h5d :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h5e :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h5f :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h60 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h61 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h62 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h63 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h64 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h65 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h66 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h67 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h68 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h69 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h6a :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h6b :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h6c :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h6d :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h6e :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h6f :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h70 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h71 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h72 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h73 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h74 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h75 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h76 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h77 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h78 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h79 :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h7a :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h7b :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h7c :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h7d :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h7e :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	7'h7f :
		rl_a23_t8 = RG_quantized_block_rl_9 ;
	default :
		rl_a23_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_141 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a24_t8 = RG_rl_141 ;
	7'h01 :
		rl_a24_t8 = RG_rl_141 ;
	7'h02 :
		rl_a24_t8 = RG_rl_141 ;
	7'h03 :
		rl_a24_t8 = RG_rl_141 ;
	7'h04 :
		rl_a24_t8 = RG_rl_141 ;
	7'h05 :
		rl_a24_t8 = RG_rl_141 ;
	7'h06 :
		rl_a24_t8 = RG_rl_141 ;
	7'h07 :
		rl_a24_t8 = RG_rl_141 ;
	7'h08 :
		rl_a24_t8 = RG_rl_141 ;
	7'h09 :
		rl_a24_t8 = RG_rl_141 ;
	7'h0a :
		rl_a24_t8 = RG_rl_141 ;
	7'h0b :
		rl_a24_t8 = RG_rl_141 ;
	7'h0c :
		rl_a24_t8 = RG_rl_141 ;
	7'h0d :
		rl_a24_t8 = RG_rl_141 ;
	7'h0e :
		rl_a24_t8 = RG_rl_141 ;
	7'h0f :
		rl_a24_t8 = RG_rl_141 ;
	7'h10 :
		rl_a24_t8 = RG_rl_141 ;
	7'h11 :
		rl_a24_t8 = RG_rl_141 ;
	7'h12 :
		rl_a24_t8 = RG_rl_141 ;
	7'h13 :
		rl_a24_t8 = RG_rl_141 ;
	7'h14 :
		rl_a24_t8 = RG_rl_141 ;
	7'h15 :
		rl_a24_t8 = RG_rl_141 ;
	7'h16 :
		rl_a24_t8 = RG_rl_141 ;
	7'h17 :
		rl_a24_t8 = RG_rl_141 ;
	7'h18 :
		rl_a24_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h19 :
		rl_a24_t8 = RG_rl_141 ;
	7'h1a :
		rl_a24_t8 = RG_rl_141 ;
	7'h1b :
		rl_a24_t8 = RG_rl_141 ;
	7'h1c :
		rl_a24_t8 = RG_rl_141 ;
	7'h1d :
		rl_a24_t8 = RG_rl_141 ;
	7'h1e :
		rl_a24_t8 = RG_rl_141 ;
	7'h1f :
		rl_a24_t8 = RG_rl_141 ;
	7'h20 :
		rl_a24_t8 = RG_rl_141 ;
	7'h21 :
		rl_a24_t8 = RG_rl_141 ;
	7'h22 :
		rl_a24_t8 = RG_rl_141 ;
	7'h23 :
		rl_a24_t8 = RG_rl_141 ;
	7'h24 :
		rl_a24_t8 = RG_rl_141 ;
	7'h25 :
		rl_a24_t8 = RG_rl_141 ;
	7'h26 :
		rl_a24_t8 = RG_rl_141 ;
	7'h27 :
		rl_a24_t8 = RG_rl_141 ;
	7'h28 :
		rl_a24_t8 = RG_rl_141 ;
	7'h29 :
		rl_a24_t8 = RG_rl_141 ;
	7'h2a :
		rl_a24_t8 = RG_rl_141 ;
	7'h2b :
		rl_a24_t8 = RG_rl_141 ;
	7'h2c :
		rl_a24_t8 = RG_rl_141 ;
	7'h2d :
		rl_a24_t8 = RG_rl_141 ;
	7'h2e :
		rl_a24_t8 = RG_rl_141 ;
	7'h2f :
		rl_a24_t8 = RG_rl_141 ;
	7'h30 :
		rl_a24_t8 = RG_rl_141 ;
	7'h31 :
		rl_a24_t8 = RG_rl_141 ;
	7'h32 :
		rl_a24_t8 = RG_rl_141 ;
	7'h33 :
		rl_a24_t8 = RG_rl_141 ;
	7'h34 :
		rl_a24_t8 = RG_rl_141 ;
	7'h35 :
		rl_a24_t8 = RG_rl_141 ;
	7'h36 :
		rl_a24_t8 = RG_rl_141 ;
	7'h37 :
		rl_a24_t8 = RG_rl_141 ;
	7'h38 :
		rl_a24_t8 = RG_rl_141 ;
	7'h39 :
		rl_a24_t8 = RG_rl_141 ;
	7'h3a :
		rl_a24_t8 = RG_rl_141 ;
	7'h3b :
		rl_a24_t8 = RG_rl_141 ;
	7'h3c :
		rl_a24_t8 = RG_rl_141 ;
	7'h3d :
		rl_a24_t8 = RG_rl_141 ;
	7'h3e :
		rl_a24_t8 = RG_rl_141 ;
	7'h3f :
		rl_a24_t8 = RG_rl_141 ;
	7'h40 :
		rl_a24_t8 = RG_rl_141 ;
	7'h41 :
		rl_a24_t8 = RG_rl_141 ;
	7'h42 :
		rl_a24_t8 = RG_rl_141 ;
	7'h43 :
		rl_a24_t8 = RG_rl_141 ;
	7'h44 :
		rl_a24_t8 = RG_rl_141 ;
	7'h45 :
		rl_a24_t8 = RG_rl_141 ;
	7'h46 :
		rl_a24_t8 = RG_rl_141 ;
	7'h47 :
		rl_a24_t8 = RG_rl_141 ;
	7'h48 :
		rl_a24_t8 = RG_rl_141 ;
	7'h49 :
		rl_a24_t8 = RG_rl_141 ;
	7'h4a :
		rl_a24_t8 = RG_rl_141 ;
	7'h4b :
		rl_a24_t8 = RG_rl_141 ;
	7'h4c :
		rl_a24_t8 = RG_rl_141 ;
	7'h4d :
		rl_a24_t8 = RG_rl_141 ;
	7'h4e :
		rl_a24_t8 = RG_rl_141 ;
	7'h4f :
		rl_a24_t8 = RG_rl_141 ;
	7'h50 :
		rl_a24_t8 = RG_rl_141 ;
	7'h51 :
		rl_a24_t8 = RG_rl_141 ;
	7'h52 :
		rl_a24_t8 = RG_rl_141 ;
	7'h53 :
		rl_a24_t8 = RG_rl_141 ;
	7'h54 :
		rl_a24_t8 = RG_rl_141 ;
	7'h55 :
		rl_a24_t8 = RG_rl_141 ;
	7'h56 :
		rl_a24_t8 = RG_rl_141 ;
	7'h57 :
		rl_a24_t8 = RG_rl_141 ;
	7'h58 :
		rl_a24_t8 = RG_rl_141 ;
	7'h59 :
		rl_a24_t8 = RG_rl_141 ;
	7'h5a :
		rl_a24_t8 = RG_rl_141 ;
	7'h5b :
		rl_a24_t8 = RG_rl_141 ;
	7'h5c :
		rl_a24_t8 = RG_rl_141 ;
	7'h5d :
		rl_a24_t8 = RG_rl_141 ;
	7'h5e :
		rl_a24_t8 = RG_rl_141 ;
	7'h5f :
		rl_a24_t8 = RG_rl_141 ;
	7'h60 :
		rl_a24_t8 = RG_rl_141 ;
	7'h61 :
		rl_a24_t8 = RG_rl_141 ;
	7'h62 :
		rl_a24_t8 = RG_rl_141 ;
	7'h63 :
		rl_a24_t8 = RG_rl_141 ;
	7'h64 :
		rl_a24_t8 = RG_rl_141 ;
	7'h65 :
		rl_a24_t8 = RG_rl_141 ;
	7'h66 :
		rl_a24_t8 = RG_rl_141 ;
	7'h67 :
		rl_a24_t8 = RG_rl_141 ;
	7'h68 :
		rl_a24_t8 = RG_rl_141 ;
	7'h69 :
		rl_a24_t8 = RG_rl_141 ;
	7'h6a :
		rl_a24_t8 = RG_rl_141 ;
	7'h6b :
		rl_a24_t8 = RG_rl_141 ;
	7'h6c :
		rl_a24_t8 = RG_rl_141 ;
	7'h6d :
		rl_a24_t8 = RG_rl_141 ;
	7'h6e :
		rl_a24_t8 = RG_rl_141 ;
	7'h6f :
		rl_a24_t8 = RG_rl_141 ;
	7'h70 :
		rl_a24_t8 = RG_rl_141 ;
	7'h71 :
		rl_a24_t8 = RG_rl_141 ;
	7'h72 :
		rl_a24_t8 = RG_rl_141 ;
	7'h73 :
		rl_a24_t8 = RG_rl_141 ;
	7'h74 :
		rl_a24_t8 = RG_rl_141 ;
	7'h75 :
		rl_a24_t8 = RG_rl_141 ;
	7'h76 :
		rl_a24_t8 = RG_rl_141 ;
	7'h77 :
		rl_a24_t8 = RG_rl_141 ;
	7'h78 :
		rl_a24_t8 = RG_rl_141 ;
	7'h79 :
		rl_a24_t8 = RG_rl_141 ;
	7'h7a :
		rl_a24_t8 = RG_rl_141 ;
	7'h7b :
		rl_a24_t8 = RG_rl_141 ;
	7'h7c :
		rl_a24_t8 = RG_rl_141 ;
	7'h7d :
		rl_a24_t8 = RG_rl_141 ;
	7'h7e :
		rl_a24_t8 = RG_rl_141 ;
	7'h7f :
		rl_a24_t8 = RG_rl_141 ;
	default :
		rl_a24_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_10 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h01 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h02 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h03 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h04 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h05 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h06 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h07 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h08 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h09 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h0a :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h0b :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h0c :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h0d :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h0e :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h0f :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h10 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h11 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h12 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h13 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h14 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h15 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h16 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h17 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h18 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h19 :
		rl_a25_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h1a :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h1b :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h1c :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h1d :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h1e :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h1f :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h20 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h21 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h22 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h23 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h24 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h25 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h26 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h27 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h28 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h29 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h2a :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h2b :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h2c :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h2d :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h2e :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h2f :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h30 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h31 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h32 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h33 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h34 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h35 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h36 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h37 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h38 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h39 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h3a :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h3b :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h3c :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h3d :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h3e :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h3f :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h40 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h41 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h42 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h43 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h44 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h45 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h46 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h47 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h48 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h49 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h4a :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h4b :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h4c :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h4d :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h4e :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h4f :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h50 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h51 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h52 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h53 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h54 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h55 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h56 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h57 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h58 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h59 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h5a :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h5b :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h5c :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h5d :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h5e :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h5f :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h60 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h61 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h62 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h63 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h64 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h65 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h66 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h67 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h68 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h69 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h6a :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h6b :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h6c :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h6d :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h6e :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h6f :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h70 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h71 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h72 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h73 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h74 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h75 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h76 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h77 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h78 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h79 :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h7a :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h7b :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h7c :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h7d :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h7e :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	7'h7f :
		rl_a25_t8 = RG_quantized_block_rl_10 ;
	default :
		rl_a25_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_142 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a26_t8 = RG_rl_142 ;
	7'h01 :
		rl_a26_t8 = RG_rl_142 ;
	7'h02 :
		rl_a26_t8 = RG_rl_142 ;
	7'h03 :
		rl_a26_t8 = RG_rl_142 ;
	7'h04 :
		rl_a26_t8 = RG_rl_142 ;
	7'h05 :
		rl_a26_t8 = RG_rl_142 ;
	7'h06 :
		rl_a26_t8 = RG_rl_142 ;
	7'h07 :
		rl_a26_t8 = RG_rl_142 ;
	7'h08 :
		rl_a26_t8 = RG_rl_142 ;
	7'h09 :
		rl_a26_t8 = RG_rl_142 ;
	7'h0a :
		rl_a26_t8 = RG_rl_142 ;
	7'h0b :
		rl_a26_t8 = RG_rl_142 ;
	7'h0c :
		rl_a26_t8 = RG_rl_142 ;
	7'h0d :
		rl_a26_t8 = RG_rl_142 ;
	7'h0e :
		rl_a26_t8 = RG_rl_142 ;
	7'h0f :
		rl_a26_t8 = RG_rl_142 ;
	7'h10 :
		rl_a26_t8 = RG_rl_142 ;
	7'h11 :
		rl_a26_t8 = RG_rl_142 ;
	7'h12 :
		rl_a26_t8 = RG_rl_142 ;
	7'h13 :
		rl_a26_t8 = RG_rl_142 ;
	7'h14 :
		rl_a26_t8 = RG_rl_142 ;
	7'h15 :
		rl_a26_t8 = RG_rl_142 ;
	7'h16 :
		rl_a26_t8 = RG_rl_142 ;
	7'h17 :
		rl_a26_t8 = RG_rl_142 ;
	7'h18 :
		rl_a26_t8 = RG_rl_142 ;
	7'h19 :
		rl_a26_t8 = RG_rl_142 ;
	7'h1a :
		rl_a26_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h1b :
		rl_a26_t8 = RG_rl_142 ;
	7'h1c :
		rl_a26_t8 = RG_rl_142 ;
	7'h1d :
		rl_a26_t8 = RG_rl_142 ;
	7'h1e :
		rl_a26_t8 = RG_rl_142 ;
	7'h1f :
		rl_a26_t8 = RG_rl_142 ;
	7'h20 :
		rl_a26_t8 = RG_rl_142 ;
	7'h21 :
		rl_a26_t8 = RG_rl_142 ;
	7'h22 :
		rl_a26_t8 = RG_rl_142 ;
	7'h23 :
		rl_a26_t8 = RG_rl_142 ;
	7'h24 :
		rl_a26_t8 = RG_rl_142 ;
	7'h25 :
		rl_a26_t8 = RG_rl_142 ;
	7'h26 :
		rl_a26_t8 = RG_rl_142 ;
	7'h27 :
		rl_a26_t8 = RG_rl_142 ;
	7'h28 :
		rl_a26_t8 = RG_rl_142 ;
	7'h29 :
		rl_a26_t8 = RG_rl_142 ;
	7'h2a :
		rl_a26_t8 = RG_rl_142 ;
	7'h2b :
		rl_a26_t8 = RG_rl_142 ;
	7'h2c :
		rl_a26_t8 = RG_rl_142 ;
	7'h2d :
		rl_a26_t8 = RG_rl_142 ;
	7'h2e :
		rl_a26_t8 = RG_rl_142 ;
	7'h2f :
		rl_a26_t8 = RG_rl_142 ;
	7'h30 :
		rl_a26_t8 = RG_rl_142 ;
	7'h31 :
		rl_a26_t8 = RG_rl_142 ;
	7'h32 :
		rl_a26_t8 = RG_rl_142 ;
	7'h33 :
		rl_a26_t8 = RG_rl_142 ;
	7'h34 :
		rl_a26_t8 = RG_rl_142 ;
	7'h35 :
		rl_a26_t8 = RG_rl_142 ;
	7'h36 :
		rl_a26_t8 = RG_rl_142 ;
	7'h37 :
		rl_a26_t8 = RG_rl_142 ;
	7'h38 :
		rl_a26_t8 = RG_rl_142 ;
	7'h39 :
		rl_a26_t8 = RG_rl_142 ;
	7'h3a :
		rl_a26_t8 = RG_rl_142 ;
	7'h3b :
		rl_a26_t8 = RG_rl_142 ;
	7'h3c :
		rl_a26_t8 = RG_rl_142 ;
	7'h3d :
		rl_a26_t8 = RG_rl_142 ;
	7'h3e :
		rl_a26_t8 = RG_rl_142 ;
	7'h3f :
		rl_a26_t8 = RG_rl_142 ;
	7'h40 :
		rl_a26_t8 = RG_rl_142 ;
	7'h41 :
		rl_a26_t8 = RG_rl_142 ;
	7'h42 :
		rl_a26_t8 = RG_rl_142 ;
	7'h43 :
		rl_a26_t8 = RG_rl_142 ;
	7'h44 :
		rl_a26_t8 = RG_rl_142 ;
	7'h45 :
		rl_a26_t8 = RG_rl_142 ;
	7'h46 :
		rl_a26_t8 = RG_rl_142 ;
	7'h47 :
		rl_a26_t8 = RG_rl_142 ;
	7'h48 :
		rl_a26_t8 = RG_rl_142 ;
	7'h49 :
		rl_a26_t8 = RG_rl_142 ;
	7'h4a :
		rl_a26_t8 = RG_rl_142 ;
	7'h4b :
		rl_a26_t8 = RG_rl_142 ;
	7'h4c :
		rl_a26_t8 = RG_rl_142 ;
	7'h4d :
		rl_a26_t8 = RG_rl_142 ;
	7'h4e :
		rl_a26_t8 = RG_rl_142 ;
	7'h4f :
		rl_a26_t8 = RG_rl_142 ;
	7'h50 :
		rl_a26_t8 = RG_rl_142 ;
	7'h51 :
		rl_a26_t8 = RG_rl_142 ;
	7'h52 :
		rl_a26_t8 = RG_rl_142 ;
	7'h53 :
		rl_a26_t8 = RG_rl_142 ;
	7'h54 :
		rl_a26_t8 = RG_rl_142 ;
	7'h55 :
		rl_a26_t8 = RG_rl_142 ;
	7'h56 :
		rl_a26_t8 = RG_rl_142 ;
	7'h57 :
		rl_a26_t8 = RG_rl_142 ;
	7'h58 :
		rl_a26_t8 = RG_rl_142 ;
	7'h59 :
		rl_a26_t8 = RG_rl_142 ;
	7'h5a :
		rl_a26_t8 = RG_rl_142 ;
	7'h5b :
		rl_a26_t8 = RG_rl_142 ;
	7'h5c :
		rl_a26_t8 = RG_rl_142 ;
	7'h5d :
		rl_a26_t8 = RG_rl_142 ;
	7'h5e :
		rl_a26_t8 = RG_rl_142 ;
	7'h5f :
		rl_a26_t8 = RG_rl_142 ;
	7'h60 :
		rl_a26_t8 = RG_rl_142 ;
	7'h61 :
		rl_a26_t8 = RG_rl_142 ;
	7'h62 :
		rl_a26_t8 = RG_rl_142 ;
	7'h63 :
		rl_a26_t8 = RG_rl_142 ;
	7'h64 :
		rl_a26_t8 = RG_rl_142 ;
	7'h65 :
		rl_a26_t8 = RG_rl_142 ;
	7'h66 :
		rl_a26_t8 = RG_rl_142 ;
	7'h67 :
		rl_a26_t8 = RG_rl_142 ;
	7'h68 :
		rl_a26_t8 = RG_rl_142 ;
	7'h69 :
		rl_a26_t8 = RG_rl_142 ;
	7'h6a :
		rl_a26_t8 = RG_rl_142 ;
	7'h6b :
		rl_a26_t8 = RG_rl_142 ;
	7'h6c :
		rl_a26_t8 = RG_rl_142 ;
	7'h6d :
		rl_a26_t8 = RG_rl_142 ;
	7'h6e :
		rl_a26_t8 = RG_rl_142 ;
	7'h6f :
		rl_a26_t8 = RG_rl_142 ;
	7'h70 :
		rl_a26_t8 = RG_rl_142 ;
	7'h71 :
		rl_a26_t8 = RG_rl_142 ;
	7'h72 :
		rl_a26_t8 = RG_rl_142 ;
	7'h73 :
		rl_a26_t8 = RG_rl_142 ;
	7'h74 :
		rl_a26_t8 = RG_rl_142 ;
	7'h75 :
		rl_a26_t8 = RG_rl_142 ;
	7'h76 :
		rl_a26_t8 = RG_rl_142 ;
	7'h77 :
		rl_a26_t8 = RG_rl_142 ;
	7'h78 :
		rl_a26_t8 = RG_rl_142 ;
	7'h79 :
		rl_a26_t8 = RG_rl_142 ;
	7'h7a :
		rl_a26_t8 = RG_rl_142 ;
	7'h7b :
		rl_a26_t8 = RG_rl_142 ;
	7'h7c :
		rl_a26_t8 = RG_rl_142 ;
	7'h7d :
		rl_a26_t8 = RG_rl_142 ;
	7'h7e :
		rl_a26_t8 = RG_rl_142 ;
	7'h7f :
		rl_a26_t8 = RG_rl_142 ;
	default :
		rl_a26_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_11 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h01 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h02 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h03 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h04 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h05 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h06 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h07 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h08 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h09 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h0a :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h0b :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h0c :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h0d :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h0e :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h0f :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h10 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h11 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h12 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h13 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h14 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h15 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h16 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h17 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h18 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h19 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h1a :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h1b :
		rl_a27_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h1c :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h1d :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h1e :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h1f :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h20 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h21 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h22 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h23 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h24 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h25 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h26 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h27 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h28 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h29 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h2a :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h2b :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h2c :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h2d :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h2e :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h2f :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h30 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h31 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h32 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h33 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h34 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h35 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h36 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h37 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h38 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h39 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h3a :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h3b :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h3c :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h3d :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h3e :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h3f :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h40 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h41 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h42 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h43 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h44 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h45 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h46 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h47 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h48 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h49 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h4a :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h4b :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h4c :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h4d :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h4e :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h4f :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h50 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h51 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h52 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h53 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h54 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h55 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h56 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h57 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h58 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h59 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h5a :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h5b :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h5c :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h5d :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h5e :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h5f :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h60 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h61 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h62 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h63 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h64 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h65 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h66 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h67 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h68 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h69 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h6a :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h6b :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h6c :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h6d :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h6e :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h6f :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h70 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h71 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h72 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h73 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h74 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h75 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h76 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h77 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h78 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h79 :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h7a :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h7b :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h7c :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h7d :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h7e :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	7'h7f :
		rl_a27_t8 = RG_quantized_block_rl_11 ;
	default :
		rl_a27_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_143 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a28_t8 = RG_rl_143 ;
	7'h01 :
		rl_a28_t8 = RG_rl_143 ;
	7'h02 :
		rl_a28_t8 = RG_rl_143 ;
	7'h03 :
		rl_a28_t8 = RG_rl_143 ;
	7'h04 :
		rl_a28_t8 = RG_rl_143 ;
	7'h05 :
		rl_a28_t8 = RG_rl_143 ;
	7'h06 :
		rl_a28_t8 = RG_rl_143 ;
	7'h07 :
		rl_a28_t8 = RG_rl_143 ;
	7'h08 :
		rl_a28_t8 = RG_rl_143 ;
	7'h09 :
		rl_a28_t8 = RG_rl_143 ;
	7'h0a :
		rl_a28_t8 = RG_rl_143 ;
	7'h0b :
		rl_a28_t8 = RG_rl_143 ;
	7'h0c :
		rl_a28_t8 = RG_rl_143 ;
	7'h0d :
		rl_a28_t8 = RG_rl_143 ;
	7'h0e :
		rl_a28_t8 = RG_rl_143 ;
	7'h0f :
		rl_a28_t8 = RG_rl_143 ;
	7'h10 :
		rl_a28_t8 = RG_rl_143 ;
	7'h11 :
		rl_a28_t8 = RG_rl_143 ;
	7'h12 :
		rl_a28_t8 = RG_rl_143 ;
	7'h13 :
		rl_a28_t8 = RG_rl_143 ;
	7'h14 :
		rl_a28_t8 = RG_rl_143 ;
	7'h15 :
		rl_a28_t8 = RG_rl_143 ;
	7'h16 :
		rl_a28_t8 = RG_rl_143 ;
	7'h17 :
		rl_a28_t8 = RG_rl_143 ;
	7'h18 :
		rl_a28_t8 = RG_rl_143 ;
	7'h19 :
		rl_a28_t8 = RG_rl_143 ;
	7'h1a :
		rl_a28_t8 = RG_rl_143 ;
	7'h1b :
		rl_a28_t8 = RG_rl_143 ;
	7'h1c :
		rl_a28_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h1d :
		rl_a28_t8 = RG_rl_143 ;
	7'h1e :
		rl_a28_t8 = RG_rl_143 ;
	7'h1f :
		rl_a28_t8 = RG_rl_143 ;
	7'h20 :
		rl_a28_t8 = RG_rl_143 ;
	7'h21 :
		rl_a28_t8 = RG_rl_143 ;
	7'h22 :
		rl_a28_t8 = RG_rl_143 ;
	7'h23 :
		rl_a28_t8 = RG_rl_143 ;
	7'h24 :
		rl_a28_t8 = RG_rl_143 ;
	7'h25 :
		rl_a28_t8 = RG_rl_143 ;
	7'h26 :
		rl_a28_t8 = RG_rl_143 ;
	7'h27 :
		rl_a28_t8 = RG_rl_143 ;
	7'h28 :
		rl_a28_t8 = RG_rl_143 ;
	7'h29 :
		rl_a28_t8 = RG_rl_143 ;
	7'h2a :
		rl_a28_t8 = RG_rl_143 ;
	7'h2b :
		rl_a28_t8 = RG_rl_143 ;
	7'h2c :
		rl_a28_t8 = RG_rl_143 ;
	7'h2d :
		rl_a28_t8 = RG_rl_143 ;
	7'h2e :
		rl_a28_t8 = RG_rl_143 ;
	7'h2f :
		rl_a28_t8 = RG_rl_143 ;
	7'h30 :
		rl_a28_t8 = RG_rl_143 ;
	7'h31 :
		rl_a28_t8 = RG_rl_143 ;
	7'h32 :
		rl_a28_t8 = RG_rl_143 ;
	7'h33 :
		rl_a28_t8 = RG_rl_143 ;
	7'h34 :
		rl_a28_t8 = RG_rl_143 ;
	7'h35 :
		rl_a28_t8 = RG_rl_143 ;
	7'h36 :
		rl_a28_t8 = RG_rl_143 ;
	7'h37 :
		rl_a28_t8 = RG_rl_143 ;
	7'h38 :
		rl_a28_t8 = RG_rl_143 ;
	7'h39 :
		rl_a28_t8 = RG_rl_143 ;
	7'h3a :
		rl_a28_t8 = RG_rl_143 ;
	7'h3b :
		rl_a28_t8 = RG_rl_143 ;
	7'h3c :
		rl_a28_t8 = RG_rl_143 ;
	7'h3d :
		rl_a28_t8 = RG_rl_143 ;
	7'h3e :
		rl_a28_t8 = RG_rl_143 ;
	7'h3f :
		rl_a28_t8 = RG_rl_143 ;
	7'h40 :
		rl_a28_t8 = RG_rl_143 ;
	7'h41 :
		rl_a28_t8 = RG_rl_143 ;
	7'h42 :
		rl_a28_t8 = RG_rl_143 ;
	7'h43 :
		rl_a28_t8 = RG_rl_143 ;
	7'h44 :
		rl_a28_t8 = RG_rl_143 ;
	7'h45 :
		rl_a28_t8 = RG_rl_143 ;
	7'h46 :
		rl_a28_t8 = RG_rl_143 ;
	7'h47 :
		rl_a28_t8 = RG_rl_143 ;
	7'h48 :
		rl_a28_t8 = RG_rl_143 ;
	7'h49 :
		rl_a28_t8 = RG_rl_143 ;
	7'h4a :
		rl_a28_t8 = RG_rl_143 ;
	7'h4b :
		rl_a28_t8 = RG_rl_143 ;
	7'h4c :
		rl_a28_t8 = RG_rl_143 ;
	7'h4d :
		rl_a28_t8 = RG_rl_143 ;
	7'h4e :
		rl_a28_t8 = RG_rl_143 ;
	7'h4f :
		rl_a28_t8 = RG_rl_143 ;
	7'h50 :
		rl_a28_t8 = RG_rl_143 ;
	7'h51 :
		rl_a28_t8 = RG_rl_143 ;
	7'h52 :
		rl_a28_t8 = RG_rl_143 ;
	7'h53 :
		rl_a28_t8 = RG_rl_143 ;
	7'h54 :
		rl_a28_t8 = RG_rl_143 ;
	7'h55 :
		rl_a28_t8 = RG_rl_143 ;
	7'h56 :
		rl_a28_t8 = RG_rl_143 ;
	7'h57 :
		rl_a28_t8 = RG_rl_143 ;
	7'h58 :
		rl_a28_t8 = RG_rl_143 ;
	7'h59 :
		rl_a28_t8 = RG_rl_143 ;
	7'h5a :
		rl_a28_t8 = RG_rl_143 ;
	7'h5b :
		rl_a28_t8 = RG_rl_143 ;
	7'h5c :
		rl_a28_t8 = RG_rl_143 ;
	7'h5d :
		rl_a28_t8 = RG_rl_143 ;
	7'h5e :
		rl_a28_t8 = RG_rl_143 ;
	7'h5f :
		rl_a28_t8 = RG_rl_143 ;
	7'h60 :
		rl_a28_t8 = RG_rl_143 ;
	7'h61 :
		rl_a28_t8 = RG_rl_143 ;
	7'h62 :
		rl_a28_t8 = RG_rl_143 ;
	7'h63 :
		rl_a28_t8 = RG_rl_143 ;
	7'h64 :
		rl_a28_t8 = RG_rl_143 ;
	7'h65 :
		rl_a28_t8 = RG_rl_143 ;
	7'h66 :
		rl_a28_t8 = RG_rl_143 ;
	7'h67 :
		rl_a28_t8 = RG_rl_143 ;
	7'h68 :
		rl_a28_t8 = RG_rl_143 ;
	7'h69 :
		rl_a28_t8 = RG_rl_143 ;
	7'h6a :
		rl_a28_t8 = RG_rl_143 ;
	7'h6b :
		rl_a28_t8 = RG_rl_143 ;
	7'h6c :
		rl_a28_t8 = RG_rl_143 ;
	7'h6d :
		rl_a28_t8 = RG_rl_143 ;
	7'h6e :
		rl_a28_t8 = RG_rl_143 ;
	7'h6f :
		rl_a28_t8 = RG_rl_143 ;
	7'h70 :
		rl_a28_t8 = RG_rl_143 ;
	7'h71 :
		rl_a28_t8 = RG_rl_143 ;
	7'h72 :
		rl_a28_t8 = RG_rl_143 ;
	7'h73 :
		rl_a28_t8 = RG_rl_143 ;
	7'h74 :
		rl_a28_t8 = RG_rl_143 ;
	7'h75 :
		rl_a28_t8 = RG_rl_143 ;
	7'h76 :
		rl_a28_t8 = RG_rl_143 ;
	7'h77 :
		rl_a28_t8 = RG_rl_143 ;
	7'h78 :
		rl_a28_t8 = RG_rl_143 ;
	7'h79 :
		rl_a28_t8 = RG_rl_143 ;
	7'h7a :
		rl_a28_t8 = RG_rl_143 ;
	7'h7b :
		rl_a28_t8 = RG_rl_143 ;
	7'h7c :
		rl_a28_t8 = RG_rl_143 ;
	7'h7d :
		rl_a28_t8 = RG_rl_143 ;
	7'h7e :
		rl_a28_t8 = RG_rl_143 ;
	7'h7f :
		rl_a28_t8 = RG_rl_143 ;
	default :
		rl_a28_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_12 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h01 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h02 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h03 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h04 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h05 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h06 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h07 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h08 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h09 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h0a :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h0b :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h0c :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h0d :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h0e :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h0f :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h10 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h11 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h12 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h13 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h14 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h15 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h16 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h17 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h18 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h19 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h1a :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h1b :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h1c :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h1d :
		rl_a29_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h1e :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h1f :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h20 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h21 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h22 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h23 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h24 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h25 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h26 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h27 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h28 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h29 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h2a :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h2b :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h2c :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h2d :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h2e :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h2f :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h30 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h31 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h32 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h33 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h34 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h35 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h36 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h37 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h38 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h39 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h3a :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h3b :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h3c :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h3d :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h3e :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h3f :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h40 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h41 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h42 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h43 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h44 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h45 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h46 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h47 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h48 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h49 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h4a :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h4b :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h4c :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h4d :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h4e :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h4f :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h50 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h51 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h52 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h53 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h54 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h55 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h56 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h57 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h58 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h59 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h5a :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h5b :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h5c :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h5d :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h5e :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h5f :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h60 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h61 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h62 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h63 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h64 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h65 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h66 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h67 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h68 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h69 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h6a :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h6b :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h6c :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h6d :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h6e :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h6f :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h70 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h71 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h72 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h73 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h74 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h75 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h76 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h77 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h78 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h79 :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h7a :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h7b :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h7c :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h7d :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h7e :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	7'h7f :
		rl_a29_t8 = RG_quantized_block_rl_12 ;
	default :
		rl_a29_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_144 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a30_t8 = RG_rl_144 ;
	7'h01 :
		rl_a30_t8 = RG_rl_144 ;
	7'h02 :
		rl_a30_t8 = RG_rl_144 ;
	7'h03 :
		rl_a30_t8 = RG_rl_144 ;
	7'h04 :
		rl_a30_t8 = RG_rl_144 ;
	7'h05 :
		rl_a30_t8 = RG_rl_144 ;
	7'h06 :
		rl_a30_t8 = RG_rl_144 ;
	7'h07 :
		rl_a30_t8 = RG_rl_144 ;
	7'h08 :
		rl_a30_t8 = RG_rl_144 ;
	7'h09 :
		rl_a30_t8 = RG_rl_144 ;
	7'h0a :
		rl_a30_t8 = RG_rl_144 ;
	7'h0b :
		rl_a30_t8 = RG_rl_144 ;
	7'h0c :
		rl_a30_t8 = RG_rl_144 ;
	7'h0d :
		rl_a30_t8 = RG_rl_144 ;
	7'h0e :
		rl_a30_t8 = RG_rl_144 ;
	7'h0f :
		rl_a30_t8 = RG_rl_144 ;
	7'h10 :
		rl_a30_t8 = RG_rl_144 ;
	7'h11 :
		rl_a30_t8 = RG_rl_144 ;
	7'h12 :
		rl_a30_t8 = RG_rl_144 ;
	7'h13 :
		rl_a30_t8 = RG_rl_144 ;
	7'h14 :
		rl_a30_t8 = RG_rl_144 ;
	7'h15 :
		rl_a30_t8 = RG_rl_144 ;
	7'h16 :
		rl_a30_t8 = RG_rl_144 ;
	7'h17 :
		rl_a30_t8 = RG_rl_144 ;
	7'h18 :
		rl_a30_t8 = RG_rl_144 ;
	7'h19 :
		rl_a30_t8 = RG_rl_144 ;
	7'h1a :
		rl_a30_t8 = RG_rl_144 ;
	7'h1b :
		rl_a30_t8 = RG_rl_144 ;
	7'h1c :
		rl_a30_t8 = RG_rl_144 ;
	7'h1d :
		rl_a30_t8 = RG_rl_144 ;
	7'h1e :
		rl_a30_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h1f :
		rl_a30_t8 = RG_rl_144 ;
	7'h20 :
		rl_a30_t8 = RG_rl_144 ;
	7'h21 :
		rl_a30_t8 = RG_rl_144 ;
	7'h22 :
		rl_a30_t8 = RG_rl_144 ;
	7'h23 :
		rl_a30_t8 = RG_rl_144 ;
	7'h24 :
		rl_a30_t8 = RG_rl_144 ;
	7'h25 :
		rl_a30_t8 = RG_rl_144 ;
	7'h26 :
		rl_a30_t8 = RG_rl_144 ;
	7'h27 :
		rl_a30_t8 = RG_rl_144 ;
	7'h28 :
		rl_a30_t8 = RG_rl_144 ;
	7'h29 :
		rl_a30_t8 = RG_rl_144 ;
	7'h2a :
		rl_a30_t8 = RG_rl_144 ;
	7'h2b :
		rl_a30_t8 = RG_rl_144 ;
	7'h2c :
		rl_a30_t8 = RG_rl_144 ;
	7'h2d :
		rl_a30_t8 = RG_rl_144 ;
	7'h2e :
		rl_a30_t8 = RG_rl_144 ;
	7'h2f :
		rl_a30_t8 = RG_rl_144 ;
	7'h30 :
		rl_a30_t8 = RG_rl_144 ;
	7'h31 :
		rl_a30_t8 = RG_rl_144 ;
	7'h32 :
		rl_a30_t8 = RG_rl_144 ;
	7'h33 :
		rl_a30_t8 = RG_rl_144 ;
	7'h34 :
		rl_a30_t8 = RG_rl_144 ;
	7'h35 :
		rl_a30_t8 = RG_rl_144 ;
	7'h36 :
		rl_a30_t8 = RG_rl_144 ;
	7'h37 :
		rl_a30_t8 = RG_rl_144 ;
	7'h38 :
		rl_a30_t8 = RG_rl_144 ;
	7'h39 :
		rl_a30_t8 = RG_rl_144 ;
	7'h3a :
		rl_a30_t8 = RG_rl_144 ;
	7'h3b :
		rl_a30_t8 = RG_rl_144 ;
	7'h3c :
		rl_a30_t8 = RG_rl_144 ;
	7'h3d :
		rl_a30_t8 = RG_rl_144 ;
	7'h3e :
		rl_a30_t8 = RG_rl_144 ;
	7'h3f :
		rl_a30_t8 = RG_rl_144 ;
	7'h40 :
		rl_a30_t8 = RG_rl_144 ;
	7'h41 :
		rl_a30_t8 = RG_rl_144 ;
	7'h42 :
		rl_a30_t8 = RG_rl_144 ;
	7'h43 :
		rl_a30_t8 = RG_rl_144 ;
	7'h44 :
		rl_a30_t8 = RG_rl_144 ;
	7'h45 :
		rl_a30_t8 = RG_rl_144 ;
	7'h46 :
		rl_a30_t8 = RG_rl_144 ;
	7'h47 :
		rl_a30_t8 = RG_rl_144 ;
	7'h48 :
		rl_a30_t8 = RG_rl_144 ;
	7'h49 :
		rl_a30_t8 = RG_rl_144 ;
	7'h4a :
		rl_a30_t8 = RG_rl_144 ;
	7'h4b :
		rl_a30_t8 = RG_rl_144 ;
	7'h4c :
		rl_a30_t8 = RG_rl_144 ;
	7'h4d :
		rl_a30_t8 = RG_rl_144 ;
	7'h4e :
		rl_a30_t8 = RG_rl_144 ;
	7'h4f :
		rl_a30_t8 = RG_rl_144 ;
	7'h50 :
		rl_a30_t8 = RG_rl_144 ;
	7'h51 :
		rl_a30_t8 = RG_rl_144 ;
	7'h52 :
		rl_a30_t8 = RG_rl_144 ;
	7'h53 :
		rl_a30_t8 = RG_rl_144 ;
	7'h54 :
		rl_a30_t8 = RG_rl_144 ;
	7'h55 :
		rl_a30_t8 = RG_rl_144 ;
	7'h56 :
		rl_a30_t8 = RG_rl_144 ;
	7'h57 :
		rl_a30_t8 = RG_rl_144 ;
	7'h58 :
		rl_a30_t8 = RG_rl_144 ;
	7'h59 :
		rl_a30_t8 = RG_rl_144 ;
	7'h5a :
		rl_a30_t8 = RG_rl_144 ;
	7'h5b :
		rl_a30_t8 = RG_rl_144 ;
	7'h5c :
		rl_a30_t8 = RG_rl_144 ;
	7'h5d :
		rl_a30_t8 = RG_rl_144 ;
	7'h5e :
		rl_a30_t8 = RG_rl_144 ;
	7'h5f :
		rl_a30_t8 = RG_rl_144 ;
	7'h60 :
		rl_a30_t8 = RG_rl_144 ;
	7'h61 :
		rl_a30_t8 = RG_rl_144 ;
	7'h62 :
		rl_a30_t8 = RG_rl_144 ;
	7'h63 :
		rl_a30_t8 = RG_rl_144 ;
	7'h64 :
		rl_a30_t8 = RG_rl_144 ;
	7'h65 :
		rl_a30_t8 = RG_rl_144 ;
	7'h66 :
		rl_a30_t8 = RG_rl_144 ;
	7'h67 :
		rl_a30_t8 = RG_rl_144 ;
	7'h68 :
		rl_a30_t8 = RG_rl_144 ;
	7'h69 :
		rl_a30_t8 = RG_rl_144 ;
	7'h6a :
		rl_a30_t8 = RG_rl_144 ;
	7'h6b :
		rl_a30_t8 = RG_rl_144 ;
	7'h6c :
		rl_a30_t8 = RG_rl_144 ;
	7'h6d :
		rl_a30_t8 = RG_rl_144 ;
	7'h6e :
		rl_a30_t8 = RG_rl_144 ;
	7'h6f :
		rl_a30_t8 = RG_rl_144 ;
	7'h70 :
		rl_a30_t8 = RG_rl_144 ;
	7'h71 :
		rl_a30_t8 = RG_rl_144 ;
	7'h72 :
		rl_a30_t8 = RG_rl_144 ;
	7'h73 :
		rl_a30_t8 = RG_rl_144 ;
	7'h74 :
		rl_a30_t8 = RG_rl_144 ;
	7'h75 :
		rl_a30_t8 = RG_rl_144 ;
	7'h76 :
		rl_a30_t8 = RG_rl_144 ;
	7'h77 :
		rl_a30_t8 = RG_rl_144 ;
	7'h78 :
		rl_a30_t8 = RG_rl_144 ;
	7'h79 :
		rl_a30_t8 = RG_rl_144 ;
	7'h7a :
		rl_a30_t8 = RG_rl_144 ;
	7'h7b :
		rl_a30_t8 = RG_rl_144 ;
	7'h7c :
		rl_a30_t8 = RG_rl_144 ;
	7'h7d :
		rl_a30_t8 = RG_rl_144 ;
	7'h7e :
		rl_a30_t8 = RG_rl_144 ;
	7'h7f :
		rl_a30_t8 = RG_rl_144 ;
	default :
		rl_a30_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_13 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h01 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h02 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h03 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h04 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h05 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h06 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h07 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h08 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h09 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h0a :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h0b :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h0c :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h0d :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h0e :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h0f :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h10 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h11 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h12 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h13 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h14 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h15 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h16 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h17 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h18 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h19 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h1a :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h1b :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h1c :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h1d :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h1e :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h1f :
		rl_a31_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h20 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h21 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h22 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h23 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h24 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h25 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h26 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h27 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h28 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h29 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h2a :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h2b :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h2c :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h2d :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h2e :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h2f :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h30 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h31 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h32 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h33 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h34 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h35 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h36 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h37 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h38 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h39 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h3a :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h3b :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h3c :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h3d :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h3e :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h3f :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h40 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h41 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h42 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h43 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h44 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h45 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h46 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h47 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h48 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h49 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h4a :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h4b :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h4c :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h4d :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h4e :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h4f :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h50 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h51 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h52 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h53 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h54 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h55 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h56 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h57 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h58 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h59 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h5a :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h5b :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h5c :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h5d :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h5e :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h5f :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h60 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h61 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h62 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h63 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h64 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h65 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h66 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h67 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h68 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h69 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h6a :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h6b :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h6c :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h6d :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h6e :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h6f :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h70 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h71 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h72 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h73 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h74 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h75 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h76 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h77 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h78 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h79 :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h7a :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h7b :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h7c :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h7d :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h7e :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	7'h7f :
		rl_a31_t8 = RG_quantized_block_rl_13 ;
	default :
		rl_a31_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_145 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a32_t8 = RG_rl_145 ;
	7'h01 :
		rl_a32_t8 = RG_rl_145 ;
	7'h02 :
		rl_a32_t8 = RG_rl_145 ;
	7'h03 :
		rl_a32_t8 = RG_rl_145 ;
	7'h04 :
		rl_a32_t8 = RG_rl_145 ;
	7'h05 :
		rl_a32_t8 = RG_rl_145 ;
	7'h06 :
		rl_a32_t8 = RG_rl_145 ;
	7'h07 :
		rl_a32_t8 = RG_rl_145 ;
	7'h08 :
		rl_a32_t8 = RG_rl_145 ;
	7'h09 :
		rl_a32_t8 = RG_rl_145 ;
	7'h0a :
		rl_a32_t8 = RG_rl_145 ;
	7'h0b :
		rl_a32_t8 = RG_rl_145 ;
	7'h0c :
		rl_a32_t8 = RG_rl_145 ;
	7'h0d :
		rl_a32_t8 = RG_rl_145 ;
	7'h0e :
		rl_a32_t8 = RG_rl_145 ;
	7'h0f :
		rl_a32_t8 = RG_rl_145 ;
	7'h10 :
		rl_a32_t8 = RG_rl_145 ;
	7'h11 :
		rl_a32_t8 = RG_rl_145 ;
	7'h12 :
		rl_a32_t8 = RG_rl_145 ;
	7'h13 :
		rl_a32_t8 = RG_rl_145 ;
	7'h14 :
		rl_a32_t8 = RG_rl_145 ;
	7'h15 :
		rl_a32_t8 = RG_rl_145 ;
	7'h16 :
		rl_a32_t8 = RG_rl_145 ;
	7'h17 :
		rl_a32_t8 = RG_rl_145 ;
	7'h18 :
		rl_a32_t8 = RG_rl_145 ;
	7'h19 :
		rl_a32_t8 = RG_rl_145 ;
	7'h1a :
		rl_a32_t8 = RG_rl_145 ;
	7'h1b :
		rl_a32_t8 = RG_rl_145 ;
	7'h1c :
		rl_a32_t8 = RG_rl_145 ;
	7'h1d :
		rl_a32_t8 = RG_rl_145 ;
	7'h1e :
		rl_a32_t8 = RG_rl_145 ;
	7'h1f :
		rl_a32_t8 = RG_rl_145 ;
	7'h20 :
		rl_a32_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h21 :
		rl_a32_t8 = RG_rl_145 ;
	7'h22 :
		rl_a32_t8 = RG_rl_145 ;
	7'h23 :
		rl_a32_t8 = RG_rl_145 ;
	7'h24 :
		rl_a32_t8 = RG_rl_145 ;
	7'h25 :
		rl_a32_t8 = RG_rl_145 ;
	7'h26 :
		rl_a32_t8 = RG_rl_145 ;
	7'h27 :
		rl_a32_t8 = RG_rl_145 ;
	7'h28 :
		rl_a32_t8 = RG_rl_145 ;
	7'h29 :
		rl_a32_t8 = RG_rl_145 ;
	7'h2a :
		rl_a32_t8 = RG_rl_145 ;
	7'h2b :
		rl_a32_t8 = RG_rl_145 ;
	7'h2c :
		rl_a32_t8 = RG_rl_145 ;
	7'h2d :
		rl_a32_t8 = RG_rl_145 ;
	7'h2e :
		rl_a32_t8 = RG_rl_145 ;
	7'h2f :
		rl_a32_t8 = RG_rl_145 ;
	7'h30 :
		rl_a32_t8 = RG_rl_145 ;
	7'h31 :
		rl_a32_t8 = RG_rl_145 ;
	7'h32 :
		rl_a32_t8 = RG_rl_145 ;
	7'h33 :
		rl_a32_t8 = RG_rl_145 ;
	7'h34 :
		rl_a32_t8 = RG_rl_145 ;
	7'h35 :
		rl_a32_t8 = RG_rl_145 ;
	7'h36 :
		rl_a32_t8 = RG_rl_145 ;
	7'h37 :
		rl_a32_t8 = RG_rl_145 ;
	7'h38 :
		rl_a32_t8 = RG_rl_145 ;
	7'h39 :
		rl_a32_t8 = RG_rl_145 ;
	7'h3a :
		rl_a32_t8 = RG_rl_145 ;
	7'h3b :
		rl_a32_t8 = RG_rl_145 ;
	7'h3c :
		rl_a32_t8 = RG_rl_145 ;
	7'h3d :
		rl_a32_t8 = RG_rl_145 ;
	7'h3e :
		rl_a32_t8 = RG_rl_145 ;
	7'h3f :
		rl_a32_t8 = RG_rl_145 ;
	7'h40 :
		rl_a32_t8 = RG_rl_145 ;
	7'h41 :
		rl_a32_t8 = RG_rl_145 ;
	7'h42 :
		rl_a32_t8 = RG_rl_145 ;
	7'h43 :
		rl_a32_t8 = RG_rl_145 ;
	7'h44 :
		rl_a32_t8 = RG_rl_145 ;
	7'h45 :
		rl_a32_t8 = RG_rl_145 ;
	7'h46 :
		rl_a32_t8 = RG_rl_145 ;
	7'h47 :
		rl_a32_t8 = RG_rl_145 ;
	7'h48 :
		rl_a32_t8 = RG_rl_145 ;
	7'h49 :
		rl_a32_t8 = RG_rl_145 ;
	7'h4a :
		rl_a32_t8 = RG_rl_145 ;
	7'h4b :
		rl_a32_t8 = RG_rl_145 ;
	7'h4c :
		rl_a32_t8 = RG_rl_145 ;
	7'h4d :
		rl_a32_t8 = RG_rl_145 ;
	7'h4e :
		rl_a32_t8 = RG_rl_145 ;
	7'h4f :
		rl_a32_t8 = RG_rl_145 ;
	7'h50 :
		rl_a32_t8 = RG_rl_145 ;
	7'h51 :
		rl_a32_t8 = RG_rl_145 ;
	7'h52 :
		rl_a32_t8 = RG_rl_145 ;
	7'h53 :
		rl_a32_t8 = RG_rl_145 ;
	7'h54 :
		rl_a32_t8 = RG_rl_145 ;
	7'h55 :
		rl_a32_t8 = RG_rl_145 ;
	7'h56 :
		rl_a32_t8 = RG_rl_145 ;
	7'h57 :
		rl_a32_t8 = RG_rl_145 ;
	7'h58 :
		rl_a32_t8 = RG_rl_145 ;
	7'h59 :
		rl_a32_t8 = RG_rl_145 ;
	7'h5a :
		rl_a32_t8 = RG_rl_145 ;
	7'h5b :
		rl_a32_t8 = RG_rl_145 ;
	7'h5c :
		rl_a32_t8 = RG_rl_145 ;
	7'h5d :
		rl_a32_t8 = RG_rl_145 ;
	7'h5e :
		rl_a32_t8 = RG_rl_145 ;
	7'h5f :
		rl_a32_t8 = RG_rl_145 ;
	7'h60 :
		rl_a32_t8 = RG_rl_145 ;
	7'h61 :
		rl_a32_t8 = RG_rl_145 ;
	7'h62 :
		rl_a32_t8 = RG_rl_145 ;
	7'h63 :
		rl_a32_t8 = RG_rl_145 ;
	7'h64 :
		rl_a32_t8 = RG_rl_145 ;
	7'h65 :
		rl_a32_t8 = RG_rl_145 ;
	7'h66 :
		rl_a32_t8 = RG_rl_145 ;
	7'h67 :
		rl_a32_t8 = RG_rl_145 ;
	7'h68 :
		rl_a32_t8 = RG_rl_145 ;
	7'h69 :
		rl_a32_t8 = RG_rl_145 ;
	7'h6a :
		rl_a32_t8 = RG_rl_145 ;
	7'h6b :
		rl_a32_t8 = RG_rl_145 ;
	7'h6c :
		rl_a32_t8 = RG_rl_145 ;
	7'h6d :
		rl_a32_t8 = RG_rl_145 ;
	7'h6e :
		rl_a32_t8 = RG_rl_145 ;
	7'h6f :
		rl_a32_t8 = RG_rl_145 ;
	7'h70 :
		rl_a32_t8 = RG_rl_145 ;
	7'h71 :
		rl_a32_t8 = RG_rl_145 ;
	7'h72 :
		rl_a32_t8 = RG_rl_145 ;
	7'h73 :
		rl_a32_t8 = RG_rl_145 ;
	7'h74 :
		rl_a32_t8 = RG_rl_145 ;
	7'h75 :
		rl_a32_t8 = RG_rl_145 ;
	7'h76 :
		rl_a32_t8 = RG_rl_145 ;
	7'h77 :
		rl_a32_t8 = RG_rl_145 ;
	7'h78 :
		rl_a32_t8 = RG_rl_145 ;
	7'h79 :
		rl_a32_t8 = RG_rl_145 ;
	7'h7a :
		rl_a32_t8 = RG_rl_145 ;
	7'h7b :
		rl_a32_t8 = RG_rl_145 ;
	7'h7c :
		rl_a32_t8 = RG_rl_145 ;
	7'h7d :
		rl_a32_t8 = RG_rl_145 ;
	7'h7e :
		rl_a32_t8 = RG_rl_145 ;
	7'h7f :
		rl_a32_t8 = RG_rl_145 ;
	default :
		rl_a32_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_14 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h01 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h02 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h03 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h04 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h05 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h06 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h07 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h08 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h09 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h0a :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h0b :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h0c :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h0d :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h0e :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h0f :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h10 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h11 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h12 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h13 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h14 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h15 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h16 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h17 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h18 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h19 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h1a :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h1b :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h1c :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h1d :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h1e :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h1f :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h20 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h21 :
		rl_a33_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h22 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h23 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h24 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h25 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h26 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h27 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h28 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h29 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h2a :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h2b :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h2c :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h2d :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h2e :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h2f :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h30 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h31 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h32 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h33 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h34 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h35 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h36 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h37 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h38 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h39 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h3a :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h3b :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h3c :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h3d :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h3e :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h3f :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h40 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h41 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h42 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h43 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h44 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h45 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h46 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h47 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h48 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h49 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h4a :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h4b :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h4c :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h4d :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h4e :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h4f :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h50 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h51 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h52 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h53 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h54 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h55 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h56 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h57 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h58 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h59 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h5a :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h5b :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h5c :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h5d :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h5e :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h5f :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h60 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h61 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h62 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h63 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h64 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h65 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h66 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h67 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h68 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h69 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h6a :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h6b :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h6c :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h6d :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h6e :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h6f :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h70 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h71 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h72 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h73 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h74 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h75 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h76 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h77 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h78 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h79 :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h7a :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h7b :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h7c :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h7d :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h7e :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	7'h7f :
		rl_a33_t8 = RG_quantized_block_rl_14 ;
	default :
		rl_a33_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_146 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a34_t8 = RG_rl_146 ;
	7'h01 :
		rl_a34_t8 = RG_rl_146 ;
	7'h02 :
		rl_a34_t8 = RG_rl_146 ;
	7'h03 :
		rl_a34_t8 = RG_rl_146 ;
	7'h04 :
		rl_a34_t8 = RG_rl_146 ;
	7'h05 :
		rl_a34_t8 = RG_rl_146 ;
	7'h06 :
		rl_a34_t8 = RG_rl_146 ;
	7'h07 :
		rl_a34_t8 = RG_rl_146 ;
	7'h08 :
		rl_a34_t8 = RG_rl_146 ;
	7'h09 :
		rl_a34_t8 = RG_rl_146 ;
	7'h0a :
		rl_a34_t8 = RG_rl_146 ;
	7'h0b :
		rl_a34_t8 = RG_rl_146 ;
	7'h0c :
		rl_a34_t8 = RG_rl_146 ;
	7'h0d :
		rl_a34_t8 = RG_rl_146 ;
	7'h0e :
		rl_a34_t8 = RG_rl_146 ;
	7'h0f :
		rl_a34_t8 = RG_rl_146 ;
	7'h10 :
		rl_a34_t8 = RG_rl_146 ;
	7'h11 :
		rl_a34_t8 = RG_rl_146 ;
	7'h12 :
		rl_a34_t8 = RG_rl_146 ;
	7'h13 :
		rl_a34_t8 = RG_rl_146 ;
	7'h14 :
		rl_a34_t8 = RG_rl_146 ;
	7'h15 :
		rl_a34_t8 = RG_rl_146 ;
	7'h16 :
		rl_a34_t8 = RG_rl_146 ;
	7'h17 :
		rl_a34_t8 = RG_rl_146 ;
	7'h18 :
		rl_a34_t8 = RG_rl_146 ;
	7'h19 :
		rl_a34_t8 = RG_rl_146 ;
	7'h1a :
		rl_a34_t8 = RG_rl_146 ;
	7'h1b :
		rl_a34_t8 = RG_rl_146 ;
	7'h1c :
		rl_a34_t8 = RG_rl_146 ;
	7'h1d :
		rl_a34_t8 = RG_rl_146 ;
	7'h1e :
		rl_a34_t8 = RG_rl_146 ;
	7'h1f :
		rl_a34_t8 = RG_rl_146 ;
	7'h20 :
		rl_a34_t8 = RG_rl_146 ;
	7'h21 :
		rl_a34_t8 = RG_rl_146 ;
	7'h22 :
		rl_a34_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h23 :
		rl_a34_t8 = RG_rl_146 ;
	7'h24 :
		rl_a34_t8 = RG_rl_146 ;
	7'h25 :
		rl_a34_t8 = RG_rl_146 ;
	7'h26 :
		rl_a34_t8 = RG_rl_146 ;
	7'h27 :
		rl_a34_t8 = RG_rl_146 ;
	7'h28 :
		rl_a34_t8 = RG_rl_146 ;
	7'h29 :
		rl_a34_t8 = RG_rl_146 ;
	7'h2a :
		rl_a34_t8 = RG_rl_146 ;
	7'h2b :
		rl_a34_t8 = RG_rl_146 ;
	7'h2c :
		rl_a34_t8 = RG_rl_146 ;
	7'h2d :
		rl_a34_t8 = RG_rl_146 ;
	7'h2e :
		rl_a34_t8 = RG_rl_146 ;
	7'h2f :
		rl_a34_t8 = RG_rl_146 ;
	7'h30 :
		rl_a34_t8 = RG_rl_146 ;
	7'h31 :
		rl_a34_t8 = RG_rl_146 ;
	7'h32 :
		rl_a34_t8 = RG_rl_146 ;
	7'h33 :
		rl_a34_t8 = RG_rl_146 ;
	7'h34 :
		rl_a34_t8 = RG_rl_146 ;
	7'h35 :
		rl_a34_t8 = RG_rl_146 ;
	7'h36 :
		rl_a34_t8 = RG_rl_146 ;
	7'h37 :
		rl_a34_t8 = RG_rl_146 ;
	7'h38 :
		rl_a34_t8 = RG_rl_146 ;
	7'h39 :
		rl_a34_t8 = RG_rl_146 ;
	7'h3a :
		rl_a34_t8 = RG_rl_146 ;
	7'h3b :
		rl_a34_t8 = RG_rl_146 ;
	7'h3c :
		rl_a34_t8 = RG_rl_146 ;
	7'h3d :
		rl_a34_t8 = RG_rl_146 ;
	7'h3e :
		rl_a34_t8 = RG_rl_146 ;
	7'h3f :
		rl_a34_t8 = RG_rl_146 ;
	7'h40 :
		rl_a34_t8 = RG_rl_146 ;
	7'h41 :
		rl_a34_t8 = RG_rl_146 ;
	7'h42 :
		rl_a34_t8 = RG_rl_146 ;
	7'h43 :
		rl_a34_t8 = RG_rl_146 ;
	7'h44 :
		rl_a34_t8 = RG_rl_146 ;
	7'h45 :
		rl_a34_t8 = RG_rl_146 ;
	7'h46 :
		rl_a34_t8 = RG_rl_146 ;
	7'h47 :
		rl_a34_t8 = RG_rl_146 ;
	7'h48 :
		rl_a34_t8 = RG_rl_146 ;
	7'h49 :
		rl_a34_t8 = RG_rl_146 ;
	7'h4a :
		rl_a34_t8 = RG_rl_146 ;
	7'h4b :
		rl_a34_t8 = RG_rl_146 ;
	7'h4c :
		rl_a34_t8 = RG_rl_146 ;
	7'h4d :
		rl_a34_t8 = RG_rl_146 ;
	7'h4e :
		rl_a34_t8 = RG_rl_146 ;
	7'h4f :
		rl_a34_t8 = RG_rl_146 ;
	7'h50 :
		rl_a34_t8 = RG_rl_146 ;
	7'h51 :
		rl_a34_t8 = RG_rl_146 ;
	7'h52 :
		rl_a34_t8 = RG_rl_146 ;
	7'h53 :
		rl_a34_t8 = RG_rl_146 ;
	7'h54 :
		rl_a34_t8 = RG_rl_146 ;
	7'h55 :
		rl_a34_t8 = RG_rl_146 ;
	7'h56 :
		rl_a34_t8 = RG_rl_146 ;
	7'h57 :
		rl_a34_t8 = RG_rl_146 ;
	7'h58 :
		rl_a34_t8 = RG_rl_146 ;
	7'h59 :
		rl_a34_t8 = RG_rl_146 ;
	7'h5a :
		rl_a34_t8 = RG_rl_146 ;
	7'h5b :
		rl_a34_t8 = RG_rl_146 ;
	7'h5c :
		rl_a34_t8 = RG_rl_146 ;
	7'h5d :
		rl_a34_t8 = RG_rl_146 ;
	7'h5e :
		rl_a34_t8 = RG_rl_146 ;
	7'h5f :
		rl_a34_t8 = RG_rl_146 ;
	7'h60 :
		rl_a34_t8 = RG_rl_146 ;
	7'h61 :
		rl_a34_t8 = RG_rl_146 ;
	7'h62 :
		rl_a34_t8 = RG_rl_146 ;
	7'h63 :
		rl_a34_t8 = RG_rl_146 ;
	7'h64 :
		rl_a34_t8 = RG_rl_146 ;
	7'h65 :
		rl_a34_t8 = RG_rl_146 ;
	7'h66 :
		rl_a34_t8 = RG_rl_146 ;
	7'h67 :
		rl_a34_t8 = RG_rl_146 ;
	7'h68 :
		rl_a34_t8 = RG_rl_146 ;
	7'h69 :
		rl_a34_t8 = RG_rl_146 ;
	7'h6a :
		rl_a34_t8 = RG_rl_146 ;
	7'h6b :
		rl_a34_t8 = RG_rl_146 ;
	7'h6c :
		rl_a34_t8 = RG_rl_146 ;
	7'h6d :
		rl_a34_t8 = RG_rl_146 ;
	7'h6e :
		rl_a34_t8 = RG_rl_146 ;
	7'h6f :
		rl_a34_t8 = RG_rl_146 ;
	7'h70 :
		rl_a34_t8 = RG_rl_146 ;
	7'h71 :
		rl_a34_t8 = RG_rl_146 ;
	7'h72 :
		rl_a34_t8 = RG_rl_146 ;
	7'h73 :
		rl_a34_t8 = RG_rl_146 ;
	7'h74 :
		rl_a34_t8 = RG_rl_146 ;
	7'h75 :
		rl_a34_t8 = RG_rl_146 ;
	7'h76 :
		rl_a34_t8 = RG_rl_146 ;
	7'h77 :
		rl_a34_t8 = RG_rl_146 ;
	7'h78 :
		rl_a34_t8 = RG_rl_146 ;
	7'h79 :
		rl_a34_t8 = RG_rl_146 ;
	7'h7a :
		rl_a34_t8 = RG_rl_146 ;
	7'h7b :
		rl_a34_t8 = RG_rl_146 ;
	7'h7c :
		rl_a34_t8 = RG_rl_146 ;
	7'h7d :
		rl_a34_t8 = RG_rl_146 ;
	7'h7e :
		rl_a34_t8 = RG_rl_146 ;
	7'h7f :
		rl_a34_t8 = RG_rl_146 ;
	default :
		rl_a34_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_15 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h01 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h02 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h03 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h04 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h05 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h06 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h07 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h08 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h09 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h0a :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h0b :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h0c :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h0d :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h0e :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h0f :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h10 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h11 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h12 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h13 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h14 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h15 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h16 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h17 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h18 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h19 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h1a :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h1b :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h1c :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h1d :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h1e :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h1f :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h20 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h21 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h22 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h23 :
		rl_a35_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h24 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h25 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h26 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h27 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h28 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h29 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h2a :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h2b :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h2c :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h2d :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h2e :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h2f :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h30 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h31 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h32 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h33 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h34 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h35 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h36 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h37 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h38 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h39 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h3a :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h3b :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h3c :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h3d :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h3e :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h3f :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h40 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h41 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h42 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h43 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h44 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h45 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h46 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h47 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h48 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h49 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h4a :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h4b :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h4c :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h4d :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h4e :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h4f :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h50 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h51 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h52 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h53 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h54 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h55 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h56 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h57 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h58 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h59 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h5a :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h5b :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h5c :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h5d :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h5e :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h5f :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h60 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h61 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h62 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h63 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h64 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h65 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h66 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h67 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h68 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h69 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h6a :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h6b :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h6c :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h6d :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h6e :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h6f :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h70 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h71 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h72 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h73 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h74 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h75 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h76 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h77 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h78 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h79 :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h7a :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h7b :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h7c :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h7d :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h7e :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	7'h7f :
		rl_a35_t8 = RG_quantized_block_rl_15 ;
	default :
		rl_a35_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_147 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a36_t8 = RG_rl_147 ;
	7'h01 :
		rl_a36_t8 = RG_rl_147 ;
	7'h02 :
		rl_a36_t8 = RG_rl_147 ;
	7'h03 :
		rl_a36_t8 = RG_rl_147 ;
	7'h04 :
		rl_a36_t8 = RG_rl_147 ;
	7'h05 :
		rl_a36_t8 = RG_rl_147 ;
	7'h06 :
		rl_a36_t8 = RG_rl_147 ;
	7'h07 :
		rl_a36_t8 = RG_rl_147 ;
	7'h08 :
		rl_a36_t8 = RG_rl_147 ;
	7'h09 :
		rl_a36_t8 = RG_rl_147 ;
	7'h0a :
		rl_a36_t8 = RG_rl_147 ;
	7'h0b :
		rl_a36_t8 = RG_rl_147 ;
	7'h0c :
		rl_a36_t8 = RG_rl_147 ;
	7'h0d :
		rl_a36_t8 = RG_rl_147 ;
	7'h0e :
		rl_a36_t8 = RG_rl_147 ;
	7'h0f :
		rl_a36_t8 = RG_rl_147 ;
	7'h10 :
		rl_a36_t8 = RG_rl_147 ;
	7'h11 :
		rl_a36_t8 = RG_rl_147 ;
	7'h12 :
		rl_a36_t8 = RG_rl_147 ;
	7'h13 :
		rl_a36_t8 = RG_rl_147 ;
	7'h14 :
		rl_a36_t8 = RG_rl_147 ;
	7'h15 :
		rl_a36_t8 = RG_rl_147 ;
	7'h16 :
		rl_a36_t8 = RG_rl_147 ;
	7'h17 :
		rl_a36_t8 = RG_rl_147 ;
	7'h18 :
		rl_a36_t8 = RG_rl_147 ;
	7'h19 :
		rl_a36_t8 = RG_rl_147 ;
	7'h1a :
		rl_a36_t8 = RG_rl_147 ;
	7'h1b :
		rl_a36_t8 = RG_rl_147 ;
	7'h1c :
		rl_a36_t8 = RG_rl_147 ;
	7'h1d :
		rl_a36_t8 = RG_rl_147 ;
	7'h1e :
		rl_a36_t8 = RG_rl_147 ;
	7'h1f :
		rl_a36_t8 = RG_rl_147 ;
	7'h20 :
		rl_a36_t8 = RG_rl_147 ;
	7'h21 :
		rl_a36_t8 = RG_rl_147 ;
	7'h22 :
		rl_a36_t8 = RG_rl_147 ;
	7'h23 :
		rl_a36_t8 = RG_rl_147 ;
	7'h24 :
		rl_a36_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h25 :
		rl_a36_t8 = RG_rl_147 ;
	7'h26 :
		rl_a36_t8 = RG_rl_147 ;
	7'h27 :
		rl_a36_t8 = RG_rl_147 ;
	7'h28 :
		rl_a36_t8 = RG_rl_147 ;
	7'h29 :
		rl_a36_t8 = RG_rl_147 ;
	7'h2a :
		rl_a36_t8 = RG_rl_147 ;
	7'h2b :
		rl_a36_t8 = RG_rl_147 ;
	7'h2c :
		rl_a36_t8 = RG_rl_147 ;
	7'h2d :
		rl_a36_t8 = RG_rl_147 ;
	7'h2e :
		rl_a36_t8 = RG_rl_147 ;
	7'h2f :
		rl_a36_t8 = RG_rl_147 ;
	7'h30 :
		rl_a36_t8 = RG_rl_147 ;
	7'h31 :
		rl_a36_t8 = RG_rl_147 ;
	7'h32 :
		rl_a36_t8 = RG_rl_147 ;
	7'h33 :
		rl_a36_t8 = RG_rl_147 ;
	7'h34 :
		rl_a36_t8 = RG_rl_147 ;
	7'h35 :
		rl_a36_t8 = RG_rl_147 ;
	7'h36 :
		rl_a36_t8 = RG_rl_147 ;
	7'h37 :
		rl_a36_t8 = RG_rl_147 ;
	7'h38 :
		rl_a36_t8 = RG_rl_147 ;
	7'h39 :
		rl_a36_t8 = RG_rl_147 ;
	7'h3a :
		rl_a36_t8 = RG_rl_147 ;
	7'h3b :
		rl_a36_t8 = RG_rl_147 ;
	7'h3c :
		rl_a36_t8 = RG_rl_147 ;
	7'h3d :
		rl_a36_t8 = RG_rl_147 ;
	7'h3e :
		rl_a36_t8 = RG_rl_147 ;
	7'h3f :
		rl_a36_t8 = RG_rl_147 ;
	7'h40 :
		rl_a36_t8 = RG_rl_147 ;
	7'h41 :
		rl_a36_t8 = RG_rl_147 ;
	7'h42 :
		rl_a36_t8 = RG_rl_147 ;
	7'h43 :
		rl_a36_t8 = RG_rl_147 ;
	7'h44 :
		rl_a36_t8 = RG_rl_147 ;
	7'h45 :
		rl_a36_t8 = RG_rl_147 ;
	7'h46 :
		rl_a36_t8 = RG_rl_147 ;
	7'h47 :
		rl_a36_t8 = RG_rl_147 ;
	7'h48 :
		rl_a36_t8 = RG_rl_147 ;
	7'h49 :
		rl_a36_t8 = RG_rl_147 ;
	7'h4a :
		rl_a36_t8 = RG_rl_147 ;
	7'h4b :
		rl_a36_t8 = RG_rl_147 ;
	7'h4c :
		rl_a36_t8 = RG_rl_147 ;
	7'h4d :
		rl_a36_t8 = RG_rl_147 ;
	7'h4e :
		rl_a36_t8 = RG_rl_147 ;
	7'h4f :
		rl_a36_t8 = RG_rl_147 ;
	7'h50 :
		rl_a36_t8 = RG_rl_147 ;
	7'h51 :
		rl_a36_t8 = RG_rl_147 ;
	7'h52 :
		rl_a36_t8 = RG_rl_147 ;
	7'h53 :
		rl_a36_t8 = RG_rl_147 ;
	7'h54 :
		rl_a36_t8 = RG_rl_147 ;
	7'h55 :
		rl_a36_t8 = RG_rl_147 ;
	7'h56 :
		rl_a36_t8 = RG_rl_147 ;
	7'h57 :
		rl_a36_t8 = RG_rl_147 ;
	7'h58 :
		rl_a36_t8 = RG_rl_147 ;
	7'h59 :
		rl_a36_t8 = RG_rl_147 ;
	7'h5a :
		rl_a36_t8 = RG_rl_147 ;
	7'h5b :
		rl_a36_t8 = RG_rl_147 ;
	7'h5c :
		rl_a36_t8 = RG_rl_147 ;
	7'h5d :
		rl_a36_t8 = RG_rl_147 ;
	7'h5e :
		rl_a36_t8 = RG_rl_147 ;
	7'h5f :
		rl_a36_t8 = RG_rl_147 ;
	7'h60 :
		rl_a36_t8 = RG_rl_147 ;
	7'h61 :
		rl_a36_t8 = RG_rl_147 ;
	7'h62 :
		rl_a36_t8 = RG_rl_147 ;
	7'h63 :
		rl_a36_t8 = RG_rl_147 ;
	7'h64 :
		rl_a36_t8 = RG_rl_147 ;
	7'h65 :
		rl_a36_t8 = RG_rl_147 ;
	7'h66 :
		rl_a36_t8 = RG_rl_147 ;
	7'h67 :
		rl_a36_t8 = RG_rl_147 ;
	7'h68 :
		rl_a36_t8 = RG_rl_147 ;
	7'h69 :
		rl_a36_t8 = RG_rl_147 ;
	7'h6a :
		rl_a36_t8 = RG_rl_147 ;
	7'h6b :
		rl_a36_t8 = RG_rl_147 ;
	7'h6c :
		rl_a36_t8 = RG_rl_147 ;
	7'h6d :
		rl_a36_t8 = RG_rl_147 ;
	7'h6e :
		rl_a36_t8 = RG_rl_147 ;
	7'h6f :
		rl_a36_t8 = RG_rl_147 ;
	7'h70 :
		rl_a36_t8 = RG_rl_147 ;
	7'h71 :
		rl_a36_t8 = RG_rl_147 ;
	7'h72 :
		rl_a36_t8 = RG_rl_147 ;
	7'h73 :
		rl_a36_t8 = RG_rl_147 ;
	7'h74 :
		rl_a36_t8 = RG_rl_147 ;
	7'h75 :
		rl_a36_t8 = RG_rl_147 ;
	7'h76 :
		rl_a36_t8 = RG_rl_147 ;
	7'h77 :
		rl_a36_t8 = RG_rl_147 ;
	7'h78 :
		rl_a36_t8 = RG_rl_147 ;
	7'h79 :
		rl_a36_t8 = RG_rl_147 ;
	7'h7a :
		rl_a36_t8 = RG_rl_147 ;
	7'h7b :
		rl_a36_t8 = RG_rl_147 ;
	7'h7c :
		rl_a36_t8 = RG_rl_147 ;
	7'h7d :
		rl_a36_t8 = RG_rl_147 ;
	7'h7e :
		rl_a36_t8 = RG_rl_147 ;
	7'h7f :
		rl_a36_t8 = RG_rl_147 ;
	default :
		rl_a36_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_16 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h01 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h02 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h03 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h04 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h05 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h06 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h07 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h08 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h09 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h0a :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h0b :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h0c :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h0d :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h0e :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h0f :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h10 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h11 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h12 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h13 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h14 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h15 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h16 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h17 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h18 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h19 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h1a :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h1b :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h1c :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h1d :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h1e :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h1f :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h20 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h21 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h22 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h23 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h24 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h25 :
		rl_a37_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h26 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h27 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h28 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h29 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h2a :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h2b :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h2c :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h2d :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h2e :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h2f :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h30 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h31 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h32 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h33 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h34 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h35 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h36 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h37 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h38 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h39 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h3a :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h3b :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h3c :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h3d :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h3e :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h3f :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h40 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h41 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h42 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h43 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h44 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h45 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h46 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h47 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h48 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h49 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h4a :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h4b :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h4c :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h4d :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h4e :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h4f :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h50 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h51 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h52 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h53 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h54 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h55 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h56 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h57 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h58 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h59 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h5a :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h5b :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h5c :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h5d :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h5e :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h5f :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h60 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h61 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h62 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h63 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h64 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h65 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h66 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h67 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h68 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h69 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h6a :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h6b :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h6c :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h6d :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h6e :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h6f :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h70 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h71 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h72 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h73 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h74 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h75 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h76 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h77 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h78 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h79 :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h7a :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h7b :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h7c :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h7d :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h7e :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	7'h7f :
		rl_a37_t8 = RG_quantized_block_rl_16 ;
	default :
		rl_a37_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_148 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a38_t8 = RG_rl_148 ;
	7'h01 :
		rl_a38_t8 = RG_rl_148 ;
	7'h02 :
		rl_a38_t8 = RG_rl_148 ;
	7'h03 :
		rl_a38_t8 = RG_rl_148 ;
	7'h04 :
		rl_a38_t8 = RG_rl_148 ;
	7'h05 :
		rl_a38_t8 = RG_rl_148 ;
	7'h06 :
		rl_a38_t8 = RG_rl_148 ;
	7'h07 :
		rl_a38_t8 = RG_rl_148 ;
	7'h08 :
		rl_a38_t8 = RG_rl_148 ;
	7'h09 :
		rl_a38_t8 = RG_rl_148 ;
	7'h0a :
		rl_a38_t8 = RG_rl_148 ;
	7'h0b :
		rl_a38_t8 = RG_rl_148 ;
	7'h0c :
		rl_a38_t8 = RG_rl_148 ;
	7'h0d :
		rl_a38_t8 = RG_rl_148 ;
	7'h0e :
		rl_a38_t8 = RG_rl_148 ;
	7'h0f :
		rl_a38_t8 = RG_rl_148 ;
	7'h10 :
		rl_a38_t8 = RG_rl_148 ;
	7'h11 :
		rl_a38_t8 = RG_rl_148 ;
	7'h12 :
		rl_a38_t8 = RG_rl_148 ;
	7'h13 :
		rl_a38_t8 = RG_rl_148 ;
	7'h14 :
		rl_a38_t8 = RG_rl_148 ;
	7'h15 :
		rl_a38_t8 = RG_rl_148 ;
	7'h16 :
		rl_a38_t8 = RG_rl_148 ;
	7'h17 :
		rl_a38_t8 = RG_rl_148 ;
	7'h18 :
		rl_a38_t8 = RG_rl_148 ;
	7'h19 :
		rl_a38_t8 = RG_rl_148 ;
	7'h1a :
		rl_a38_t8 = RG_rl_148 ;
	7'h1b :
		rl_a38_t8 = RG_rl_148 ;
	7'h1c :
		rl_a38_t8 = RG_rl_148 ;
	7'h1d :
		rl_a38_t8 = RG_rl_148 ;
	7'h1e :
		rl_a38_t8 = RG_rl_148 ;
	7'h1f :
		rl_a38_t8 = RG_rl_148 ;
	7'h20 :
		rl_a38_t8 = RG_rl_148 ;
	7'h21 :
		rl_a38_t8 = RG_rl_148 ;
	7'h22 :
		rl_a38_t8 = RG_rl_148 ;
	7'h23 :
		rl_a38_t8 = RG_rl_148 ;
	7'h24 :
		rl_a38_t8 = RG_rl_148 ;
	7'h25 :
		rl_a38_t8 = RG_rl_148 ;
	7'h26 :
		rl_a38_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h27 :
		rl_a38_t8 = RG_rl_148 ;
	7'h28 :
		rl_a38_t8 = RG_rl_148 ;
	7'h29 :
		rl_a38_t8 = RG_rl_148 ;
	7'h2a :
		rl_a38_t8 = RG_rl_148 ;
	7'h2b :
		rl_a38_t8 = RG_rl_148 ;
	7'h2c :
		rl_a38_t8 = RG_rl_148 ;
	7'h2d :
		rl_a38_t8 = RG_rl_148 ;
	7'h2e :
		rl_a38_t8 = RG_rl_148 ;
	7'h2f :
		rl_a38_t8 = RG_rl_148 ;
	7'h30 :
		rl_a38_t8 = RG_rl_148 ;
	7'h31 :
		rl_a38_t8 = RG_rl_148 ;
	7'h32 :
		rl_a38_t8 = RG_rl_148 ;
	7'h33 :
		rl_a38_t8 = RG_rl_148 ;
	7'h34 :
		rl_a38_t8 = RG_rl_148 ;
	7'h35 :
		rl_a38_t8 = RG_rl_148 ;
	7'h36 :
		rl_a38_t8 = RG_rl_148 ;
	7'h37 :
		rl_a38_t8 = RG_rl_148 ;
	7'h38 :
		rl_a38_t8 = RG_rl_148 ;
	7'h39 :
		rl_a38_t8 = RG_rl_148 ;
	7'h3a :
		rl_a38_t8 = RG_rl_148 ;
	7'h3b :
		rl_a38_t8 = RG_rl_148 ;
	7'h3c :
		rl_a38_t8 = RG_rl_148 ;
	7'h3d :
		rl_a38_t8 = RG_rl_148 ;
	7'h3e :
		rl_a38_t8 = RG_rl_148 ;
	7'h3f :
		rl_a38_t8 = RG_rl_148 ;
	7'h40 :
		rl_a38_t8 = RG_rl_148 ;
	7'h41 :
		rl_a38_t8 = RG_rl_148 ;
	7'h42 :
		rl_a38_t8 = RG_rl_148 ;
	7'h43 :
		rl_a38_t8 = RG_rl_148 ;
	7'h44 :
		rl_a38_t8 = RG_rl_148 ;
	7'h45 :
		rl_a38_t8 = RG_rl_148 ;
	7'h46 :
		rl_a38_t8 = RG_rl_148 ;
	7'h47 :
		rl_a38_t8 = RG_rl_148 ;
	7'h48 :
		rl_a38_t8 = RG_rl_148 ;
	7'h49 :
		rl_a38_t8 = RG_rl_148 ;
	7'h4a :
		rl_a38_t8 = RG_rl_148 ;
	7'h4b :
		rl_a38_t8 = RG_rl_148 ;
	7'h4c :
		rl_a38_t8 = RG_rl_148 ;
	7'h4d :
		rl_a38_t8 = RG_rl_148 ;
	7'h4e :
		rl_a38_t8 = RG_rl_148 ;
	7'h4f :
		rl_a38_t8 = RG_rl_148 ;
	7'h50 :
		rl_a38_t8 = RG_rl_148 ;
	7'h51 :
		rl_a38_t8 = RG_rl_148 ;
	7'h52 :
		rl_a38_t8 = RG_rl_148 ;
	7'h53 :
		rl_a38_t8 = RG_rl_148 ;
	7'h54 :
		rl_a38_t8 = RG_rl_148 ;
	7'h55 :
		rl_a38_t8 = RG_rl_148 ;
	7'h56 :
		rl_a38_t8 = RG_rl_148 ;
	7'h57 :
		rl_a38_t8 = RG_rl_148 ;
	7'h58 :
		rl_a38_t8 = RG_rl_148 ;
	7'h59 :
		rl_a38_t8 = RG_rl_148 ;
	7'h5a :
		rl_a38_t8 = RG_rl_148 ;
	7'h5b :
		rl_a38_t8 = RG_rl_148 ;
	7'h5c :
		rl_a38_t8 = RG_rl_148 ;
	7'h5d :
		rl_a38_t8 = RG_rl_148 ;
	7'h5e :
		rl_a38_t8 = RG_rl_148 ;
	7'h5f :
		rl_a38_t8 = RG_rl_148 ;
	7'h60 :
		rl_a38_t8 = RG_rl_148 ;
	7'h61 :
		rl_a38_t8 = RG_rl_148 ;
	7'h62 :
		rl_a38_t8 = RG_rl_148 ;
	7'h63 :
		rl_a38_t8 = RG_rl_148 ;
	7'h64 :
		rl_a38_t8 = RG_rl_148 ;
	7'h65 :
		rl_a38_t8 = RG_rl_148 ;
	7'h66 :
		rl_a38_t8 = RG_rl_148 ;
	7'h67 :
		rl_a38_t8 = RG_rl_148 ;
	7'h68 :
		rl_a38_t8 = RG_rl_148 ;
	7'h69 :
		rl_a38_t8 = RG_rl_148 ;
	7'h6a :
		rl_a38_t8 = RG_rl_148 ;
	7'h6b :
		rl_a38_t8 = RG_rl_148 ;
	7'h6c :
		rl_a38_t8 = RG_rl_148 ;
	7'h6d :
		rl_a38_t8 = RG_rl_148 ;
	7'h6e :
		rl_a38_t8 = RG_rl_148 ;
	7'h6f :
		rl_a38_t8 = RG_rl_148 ;
	7'h70 :
		rl_a38_t8 = RG_rl_148 ;
	7'h71 :
		rl_a38_t8 = RG_rl_148 ;
	7'h72 :
		rl_a38_t8 = RG_rl_148 ;
	7'h73 :
		rl_a38_t8 = RG_rl_148 ;
	7'h74 :
		rl_a38_t8 = RG_rl_148 ;
	7'h75 :
		rl_a38_t8 = RG_rl_148 ;
	7'h76 :
		rl_a38_t8 = RG_rl_148 ;
	7'h77 :
		rl_a38_t8 = RG_rl_148 ;
	7'h78 :
		rl_a38_t8 = RG_rl_148 ;
	7'h79 :
		rl_a38_t8 = RG_rl_148 ;
	7'h7a :
		rl_a38_t8 = RG_rl_148 ;
	7'h7b :
		rl_a38_t8 = RG_rl_148 ;
	7'h7c :
		rl_a38_t8 = RG_rl_148 ;
	7'h7d :
		rl_a38_t8 = RG_rl_148 ;
	7'h7e :
		rl_a38_t8 = RG_rl_148 ;
	7'h7f :
		rl_a38_t8 = RG_rl_148 ;
	default :
		rl_a38_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_17 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h01 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h02 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h03 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h04 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h05 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h06 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h07 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h08 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h09 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h0a :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h0b :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h0c :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h0d :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h0e :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h0f :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h10 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h11 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h12 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h13 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h14 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h15 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h16 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h17 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h18 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h19 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h1a :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h1b :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h1c :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h1d :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h1e :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h1f :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h20 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h21 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h22 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h23 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h24 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h25 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h26 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h27 :
		rl_a39_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h28 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h29 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h2a :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h2b :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h2c :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h2d :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h2e :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h2f :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h30 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h31 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h32 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h33 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h34 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h35 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h36 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h37 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h38 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h39 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h3a :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h3b :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h3c :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h3d :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h3e :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h3f :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h40 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h41 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h42 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h43 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h44 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h45 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h46 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h47 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h48 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h49 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h4a :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h4b :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h4c :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h4d :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h4e :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h4f :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h50 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h51 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h52 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h53 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h54 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h55 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h56 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h57 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h58 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h59 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h5a :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h5b :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h5c :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h5d :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h5e :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h5f :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h60 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h61 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h62 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h63 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h64 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h65 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h66 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h67 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h68 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h69 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h6a :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h6b :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h6c :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h6d :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h6e :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h6f :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h70 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h71 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h72 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h73 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h74 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h75 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h76 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h77 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h78 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h79 :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h7a :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h7b :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h7c :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h7d :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h7e :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	7'h7f :
		rl_a39_t8 = RG_quantized_block_rl_17 ;
	default :
		rl_a39_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_149 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a40_t8 = RG_rl_149 ;
	7'h01 :
		rl_a40_t8 = RG_rl_149 ;
	7'h02 :
		rl_a40_t8 = RG_rl_149 ;
	7'h03 :
		rl_a40_t8 = RG_rl_149 ;
	7'h04 :
		rl_a40_t8 = RG_rl_149 ;
	7'h05 :
		rl_a40_t8 = RG_rl_149 ;
	7'h06 :
		rl_a40_t8 = RG_rl_149 ;
	7'h07 :
		rl_a40_t8 = RG_rl_149 ;
	7'h08 :
		rl_a40_t8 = RG_rl_149 ;
	7'h09 :
		rl_a40_t8 = RG_rl_149 ;
	7'h0a :
		rl_a40_t8 = RG_rl_149 ;
	7'h0b :
		rl_a40_t8 = RG_rl_149 ;
	7'h0c :
		rl_a40_t8 = RG_rl_149 ;
	7'h0d :
		rl_a40_t8 = RG_rl_149 ;
	7'h0e :
		rl_a40_t8 = RG_rl_149 ;
	7'h0f :
		rl_a40_t8 = RG_rl_149 ;
	7'h10 :
		rl_a40_t8 = RG_rl_149 ;
	7'h11 :
		rl_a40_t8 = RG_rl_149 ;
	7'h12 :
		rl_a40_t8 = RG_rl_149 ;
	7'h13 :
		rl_a40_t8 = RG_rl_149 ;
	7'h14 :
		rl_a40_t8 = RG_rl_149 ;
	7'h15 :
		rl_a40_t8 = RG_rl_149 ;
	7'h16 :
		rl_a40_t8 = RG_rl_149 ;
	7'h17 :
		rl_a40_t8 = RG_rl_149 ;
	7'h18 :
		rl_a40_t8 = RG_rl_149 ;
	7'h19 :
		rl_a40_t8 = RG_rl_149 ;
	7'h1a :
		rl_a40_t8 = RG_rl_149 ;
	7'h1b :
		rl_a40_t8 = RG_rl_149 ;
	7'h1c :
		rl_a40_t8 = RG_rl_149 ;
	7'h1d :
		rl_a40_t8 = RG_rl_149 ;
	7'h1e :
		rl_a40_t8 = RG_rl_149 ;
	7'h1f :
		rl_a40_t8 = RG_rl_149 ;
	7'h20 :
		rl_a40_t8 = RG_rl_149 ;
	7'h21 :
		rl_a40_t8 = RG_rl_149 ;
	7'h22 :
		rl_a40_t8 = RG_rl_149 ;
	7'h23 :
		rl_a40_t8 = RG_rl_149 ;
	7'h24 :
		rl_a40_t8 = RG_rl_149 ;
	7'h25 :
		rl_a40_t8 = RG_rl_149 ;
	7'h26 :
		rl_a40_t8 = RG_rl_149 ;
	7'h27 :
		rl_a40_t8 = RG_rl_149 ;
	7'h28 :
		rl_a40_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h29 :
		rl_a40_t8 = RG_rl_149 ;
	7'h2a :
		rl_a40_t8 = RG_rl_149 ;
	7'h2b :
		rl_a40_t8 = RG_rl_149 ;
	7'h2c :
		rl_a40_t8 = RG_rl_149 ;
	7'h2d :
		rl_a40_t8 = RG_rl_149 ;
	7'h2e :
		rl_a40_t8 = RG_rl_149 ;
	7'h2f :
		rl_a40_t8 = RG_rl_149 ;
	7'h30 :
		rl_a40_t8 = RG_rl_149 ;
	7'h31 :
		rl_a40_t8 = RG_rl_149 ;
	7'h32 :
		rl_a40_t8 = RG_rl_149 ;
	7'h33 :
		rl_a40_t8 = RG_rl_149 ;
	7'h34 :
		rl_a40_t8 = RG_rl_149 ;
	7'h35 :
		rl_a40_t8 = RG_rl_149 ;
	7'h36 :
		rl_a40_t8 = RG_rl_149 ;
	7'h37 :
		rl_a40_t8 = RG_rl_149 ;
	7'h38 :
		rl_a40_t8 = RG_rl_149 ;
	7'h39 :
		rl_a40_t8 = RG_rl_149 ;
	7'h3a :
		rl_a40_t8 = RG_rl_149 ;
	7'h3b :
		rl_a40_t8 = RG_rl_149 ;
	7'h3c :
		rl_a40_t8 = RG_rl_149 ;
	7'h3d :
		rl_a40_t8 = RG_rl_149 ;
	7'h3e :
		rl_a40_t8 = RG_rl_149 ;
	7'h3f :
		rl_a40_t8 = RG_rl_149 ;
	7'h40 :
		rl_a40_t8 = RG_rl_149 ;
	7'h41 :
		rl_a40_t8 = RG_rl_149 ;
	7'h42 :
		rl_a40_t8 = RG_rl_149 ;
	7'h43 :
		rl_a40_t8 = RG_rl_149 ;
	7'h44 :
		rl_a40_t8 = RG_rl_149 ;
	7'h45 :
		rl_a40_t8 = RG_rl_149 ;
	7'h46 :
		rl_a40_t8 = RG_rl_149 ;
	7'h47 :
		rl_a40_t8 = RG_rl_149 ;
	7'h48 :
		rl_a40_t8 = RG_rl_149 ;
	7'h49 :
		rl_a40_t8 = RG_rl_149 ;
	7'h4a :
		rl_a40_t8 = RG_rl_149 ;
	7'h4b :
		rl_a40_t8 = RG_rl_149 ;
	7'h4c :
		rl_a40_t8 = RG_rl_149 ;
	7'h4d :
		rl_a40_t8 = RG_rl_149 ;
	7'h4e :
		rl_a40_t8 = RG_rl_149 ;
	7'h4f :
		rl_a40_t8 = RG_rl_149 ;
	7'h50 :
		rl_a40_t8 = RG_rl_149 ;
	7'h51 :
		rl_a40_t8 = RG_rl_149 ;
	7'h52 :
		rl_a40_t8 = RG_rl_149 ;
	7'h53 :
		rl_a40_t8 = RG_rl_149 ;
	7'h54 :
		rl_a40_t8 = RG_rl_149 ;
	7'h55 :
		rl_a40_t8 = RG_rl_149 ;
	7'h56 :
		rl_a40_t8 = RG_rl_149 ;
	7'h57 :
		rl_a40_t8 = RG_rl_149 ;
	7'h58 :
		rl_a40_t8 = RG_rl_149 ;
	7'h59 :
		rl_a40_t8 = RG_rl_149 ;
	7'h5a :
		rl_a40_t8 = RG_rl_149 ;
	7'h5b :
		rl_a40_t8 = RG_rl_149 ;
	7'h5c :
		rl_a40_t8 = RG_rl_149 ;
	7'h5d :
		rl_a40_t8 = RG_rl_149 ;
	7'h5e :
		rl_a40_t8 = RG_rl_149 ;
	7'h5f :
		rl_a40_t8 = RG_rl_149 ;
	7'h60 :
		rl_a40_t8 = RG_rl_149 ;
	7'h61 :
		rl_a40_t8 = RG_rl_149 ;
	7'h62 :
		rl_a40_t8 = RG_rl_149 ;
	7'h63 :
		rl_a40_t8 = RG_rl_149 ;
	7'h64 :
		rl_a40_t8 = RG_rl_149 ;
	7'h65 :
		rl_a40_t8 = RG_rl_149 ;
	7'h66 :
		rl_a40_t8 = RG_rl_149 ;
	7'h67 :
		rl_a40_t8 = RG_rl_149 ;
	7'h68 :
		rl_a40_t8 = RG_rl_149 ;
	7'h69 :
		rl_a40_t8 = RG_rl_149 ;
	7'h6a :
		rl_a40_t8 = RG_rl_149 ;
	7'h6b :
		rl_a40_t8 = RG_rl_149 ;
	7'h6c :
		rl_a40_t8 = RG_rl_149 ;
	7'h6d :
		rl_a40_t8 = RG_rl_149 ;
	7'h6e :
		rl_a40_t8 = RG_rl_149 ;
	7'h6f :
		rl_a40_t8 = RG_rl_149 ;
	7'h70 :
		rl_a40_t8 = RG_rl_149 ;
	7'h71 :
		rl_a40_t8 = RG_rl_149 ;
	7'h72 :
		rl_a40_t8 = RG_rl_149 ;
	7'h73 :
		rl_a40_t8 = RG_rl_149 ;
	7'h74 :
		rl_a40_t8 = RG_rl_149 ;
	7'h75 :
		rl_a40_t8 = RG_rl_149 ;
	7'h76 :
		rl_a40_t8 = RG_rl_149 ;
	7'h77 :
		rl_a40_t8 = RG_rl_149 ;
	7'h78 :
		rl_a40_t8 = RG_rl_149 ;
	7'h79 :
		rl_a40_t8 = RG_rl_149 ;
	7'h7a :
		rl_a40_t8 = RG_rl_149 ;
	7'h7b :
		rl_a40_t8 = RG_rl_149 ;
	7'h7c :
		rl_a40_t8 = RG_rl_149 ;
	7'h7d :
		rl_a40_t8 = RG_rl_149 ;
	7'h7e :
		rl_a40_t8 = RG_rl_149 ;
	7'h7f :
		rl_a40_t8 = RG_rl_149 ;
	default :
		rl_a40_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_18 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h01 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h02 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h03 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h04 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h05 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h06 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h07 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h08 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h09 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h0a :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h0b :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h0c :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h0d :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h0e :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h0f :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h10 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h11 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h12 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h13 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h14 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h15 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h16 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h17 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h18 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h19 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h1a :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h1b :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h1c :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h1d :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h1e :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h1f :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h20 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h21 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h22 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h23 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h24 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h25 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h26 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h27 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h28 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h29 :
		rl_a41_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h2a :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h2b :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h2c :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h2d :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h2e :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h2f :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h30 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h31 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h32 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h33 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h34 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h35 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h36 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h37 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h38 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h39 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h3a :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h3b :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h3c :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h3d :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h3e :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h3f :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h40 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h41 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h42 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h43 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h44 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h45 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h46 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h47 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h48 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h49 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h4a :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h4b :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h4c :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h4d :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h4e :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h4f :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h50 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h51 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h52 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h53 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h54 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h55 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h56 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h57 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h58 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h59 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h5a :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h5b :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h5c :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h5d :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h5e :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h5f :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h60 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h61 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h62 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h63 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h64 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h65 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h66 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h67 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h68 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h69 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h6a :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h6b :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h6c :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h6d :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h6e :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h6f :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h70 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h71 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h72 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h73 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h74 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h75 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h76 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h77 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h78 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h79 :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h7a :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h7b :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h7c :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h7d :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h7e :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	7'h7f :
		rl_a41_t8 = RG_quantized_block_rl_18 ;
	default :
		rl_a41_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_150 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a42_t8 = RG_rl_150 ;
	7'h01 :
		rl_a42_t8 = RG_rl_150 ;
	7'h02 :
		rl_a42_t8 = RG_rl_150 ;
	7'h03 :
		rl_a42_t8 = RG_rl_150 ;
	7'h04 :
		rl_a42_t8 = RG_rl_150 ;
	7'h05 :
		rl_a42_t8 = RG_rl_150 ;
	7'h06 :
		rl_a42_t8 = RG_rl_150 ;
	7'h07 :
		rl_a42_t8 = RG_rl_150 ;
	7'h08 :
		rl_a42_t8 = RG_rl_150 ;
	7'h09 :
		rl_a42_t8 = RG_rl_150 ;
	7'h0a :
		rl_a42_t8 = RG_rl_150 ;
	7'h0b :
		rl_a42_t8 = RG_rl_150 ;
	7'h0c :
		rl_a42_t8 = RG_rl_150 ;
	7'h0d :
		rl_a42_t8 = RG_rl_150 ;
	7'h0e :
		rl_a42_t8 = RG_rl_150 ;
	7'h0f :
		rl_a42_t8 = RG_rl_150 ;
	7'h10 :
		rl_a42_t8 = RG_rl_150 ;
	7'h11 :
		rl_a42_t8 = RG_rl_150 ;
	7'h12 :
		rl_a42_t8 = RG_rl_150 ;
	7'h13 :
		rl_a42_t8 = RG_rl_150 ;
	7'h14 :
		rl_a42_t8 = RG_rl_150 ;
	7'h15 :
		rl_a42_t8 = RG_rl_150 ;
	7'h16 :
		rl_a42_t8 = RG_rl_150 ;
	7'h17 :
		rl_a42_t8 = RG_rl_150 ;
	7'h18 :
		rl_a42_t8 = RG_rl_150 ;
	7'h19 :
		rl_a42_t8 = RG_rl_150 ;
	7'h1a :
		rl_a42_t8 = RG_rl_150 ;
	7'h1b :
		rl_a42_t8 = RG_rl_150 ;
	7'h1c :
		rl_a42_t8 = RG_rl_150 ;
	7'h1d :
		rl_a42_t8 = RG_rl_150 ;
	7'h1e :
		rl_a42_t8 = RG_rl_150 ;
	7'h1f :
		rl_a42_t8 = RG_rl_150 ;
	7'h20 :
		rl_a42_t8 = RG_rl_150 ;
	7'h21 :
		rl_a42_t8 = RG_rl_150 ;
	7'h22 :
		rl_a42_t8 = RG_rl_150 ;
	7'h23 :
		rl_a42_t8 = RG_rl_150 ;
	7'h24 :
		rl_a42_t8 = RG_rl_150 ;
	7'h25 :
		rl_a42_t8 = RG_rl_150 ;
	7'h26 :
		rl_a42_t8 = RG_rl_150 ;
	7'h27 :
		rl_a42_t8 = RG_rl_150 ;
	7'h28 :
		rl_a42_t8 = RG_rl_150 ;
	7'h29 :
		rl_a42_t8 = RG_rl_150 ;
	7'h2a :
		rl_a42_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h2b :
		rl_a42_t8 = RG_rl_150 ;
	7'h2c :
		rl_a42_t8 = RG_rl_150 ;
	7'h2d :
		rl_a42_t8 = RG_rl_150 ;
	7'h2e :
		rl_a42_t8 = RG_rl_150 ;
	7'h2f :
		rl_a42_t8 = RG_rl_150 ;
	7'h30 :
		rl_a42_t8 = RG_rl_150 ;
	7'h31 :
		rl_a42_t8 = RG_rl_150 ;
	7'h32 :
		rl_a42_t8 = RG_rl_150 ;
	7'h33 :
		rl_a42_t8 = RG_rl_150 ;
	7'h34 :
		rl_a42_t8 = RG_rl_150 ;
	7'h35 :
		rl_a42_t8 = RG_rl_150 ;
	7'h36 :
		rl_a42_t8 = RG_rl_150 ;
	7'h37 :
		rl_a42_t8 = RG_rl_150 ;
	7'h38 :
		rl_a42_t8 = RG_rl_150 ;
	7'h39 :
		rl_a42_t8 = RG_rl_150 ;
	7'h3a :
		rl_a42_t8 = RG_rl_150 ;
	7'h3b :
		rl_a42_t8 = RG_rl_150 ;
	7'h3c :
		rl_a42_t8 = RG_rl_150 ;
	7'h3d :
		rl_a42_t8 = RG_rl_150 ;
	7'h3e :
		rl_a42_t8 = RG_rl_150 ;
	7'h3f :
		rl_a42_t8 = RG_rl_150 ;
	7'h40 :
		rl_a42_t8 = RG_rl_150 ;
	7'h41 :
		rl_a42_t8 = RG_rl_150 ;
	7'h42 :
		rl_a42_t8 = RG_rl_150 ;
	7'h43 :
		rl_a42_t8 = RG_rl_150 ;
	7'h44 :
		rl_a42_t8 = RG_rl_150 ;
	7'h45 :
		rl_a42_t8 = RG_rl_150 ;
	7'h46 :
		rl_a42_t8 = RG_rl_150 ;
	7'h47 :
		rl_a42_t8 = RG_rl_150 ;
	7'h48 :
		rl_a42_t8 = RG_rl_150 ;
	7'h49 :
		rl_a42_t8 = RG_rl_150 ;
	7'h4a :
		rl_a42_t8 = RG_rl_150 ;
	7'h4b :
		rl_a42_t8 = RG_rl_150 ;
	7'h4c :
		rl_a42_t8 = RG_rl_150 ;
	7'h4d :
		rl_a42_t8 = RG_rl_150 ;
	7'h4e :
		rl_a42_t8 = RG_rl_150 ;
	7'h4f :
		rl_a42_t8 = RG_rl_150 ;
	7'h50 :
		rl_a42_t8 = RG_rl_150 ;
	7'h51 :
		rl_a42_t8 = RG_rl_150 ;
	7'h52 :
		rl_a42_t8 = RG_rl_150 ;
	7'h53 :
		rl_a42_t8 = RG_rl_150 ;
	7'h54 :
		rl_a42_t8 = RG_rl_150 ;
	7'h55 :
		rl_a42_t8 = RG_rl_150 ;
	7'h56 :
		rl_a42_t8 = RG_rl_150 ;
	7'h57 :
		rl_a42_t8 = RG_rl_150 ;
	7'h58 :
		rl_a42_t8 = RG_rl_150 ;
	7'h59 :
		rl_a42_t8 = RG_rl_150 ;
	7'h5a :
		rl_a42_t8 = RG_rl_150 ;
	7'h5b :
		rl_a42_t8 = RG_rl_150 ;
	7'h5c :
		rl_a42_t8 = RG_rl_150 ;
	7'h5d :
		rl_a42_t8 = RG_rl_150 ;
	7'h5e :
		rl_a42_t8 = RG_rl_150 ;
	7'h5f :
		rl_a42_t8 = RG_rl_150 ;
	7'h60 :
		rl_a42_t8 = RG_rl_150 ;
	7'h61 :
		rl_a42_t8 = RG_rl_150 ;
	7'h62 :
		rl_a42_t8 = RG_rl_150 ;
	7'h63 :
		rl_a42_t8 = RG_rl_150 ;
	7'h64 :
		rl_a42_t8 = RG_rl_150 ;
	7'h65 :
		rl_a42_t8 = RG_rl_150 ;
	7'h66 :
		rl_a42_t8 = RG_rl_150 ;
	7'h67 :
		rl_a42_t8 = RG_rl_150 ;
	7'h68 :
		rl_a42_t8 = RG_rl_150 ;
	7'h69 :
		rl_a42_t8 = RG_rl_150 ;
	7'h6a :
		rl_a42_t8 = RG_rl_150 ;
	7'h6b :
		rl_a42_t8 = RG_rl_150 ;
	7'h6c :
		rl_a42_t8 = RG_rl_150 ;
	7'h6d :
		rl_a42_t8 = RG_rl_150 ;
	7'h6e :
		rl_a42_t8 = RG_rl_150 ;
	7'h6f :
		rl_a42_t8 = RG_rl_150 ;
	7'h70 :
		rl_a42_t8 = RG_rl_150 ;
	7'h71 :
		rl_a42_t8 = RG_rl_150 ;
	7'h72 :
		rl_a42_t8 = RG_rl_150 ;
	7'h73 :
		rl_a42_t8 = RG_rl_150 ;
	7'h74 :
		rl_a42_t8 = RG_rl_150 ;
	7'h75 :
		rl_a42_t8 = RG_rl_150 ;
	7'h76 :
		rl_a42_t8 = RG_rl_150 ;
	7'h77 :
		rl_a42_t8 = RG_rl_150 ;
	7'h78 :
		rl_a42_t8 = RG_rl_150 ;
	7'h79 :
		rl_a42_t8 = RG_rl_150 ;
	7'h7a :
		rl_a42_t8 = RG_rl_150 ;
	7'h7b :
		rl_a42_t8 = RG_rl_150 ;
	7'h7c :
		rl_a42_t8 = RG_rl_150 ;
	7'h7d :
		rl_a42_t8 = RG_rl_150 ;
	7'h7e :
		rl_a42_t8 = RG_rl_150 ;
	7'h7f :
		rl_a42_t8 = RG_rl_150 ;
	default :
		rl_a42_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_19 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h01 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h02 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h03 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h04 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h05 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h06 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h07 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h08 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h09 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h0a :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h0b :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h0c :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h0d :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h0e :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h0f :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h10 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h11 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h12 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h13 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h14 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h15 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h16 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h17 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h18 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h19 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h1a :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h1b :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h1c :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h1d :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h1e :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h1f :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h20 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h21 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h22 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h23 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h24 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h25 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h26 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h27 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h28 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h29 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h2a :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h2b :
		rl_a43_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h2c :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h2d :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h2e :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h2f :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h30 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h31 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h32 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h33 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h34 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h35 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h36 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h37 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h38 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h39 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h3a :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h3b :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h3c :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h3d :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h3e :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h3f :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h40 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h41 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h42 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h43 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h44 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h45 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h46 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h47 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h48 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h49 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h4a :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h4b :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h4c :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h4d :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h4e :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h4f :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h50 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h51 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h52 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h53 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h54 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h55 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h56 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h57 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h58 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h59 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h5a :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h5b :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h5c :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h5d :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h5e :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h5f :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h60 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h61 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h62 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h63 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h64 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h65 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h66 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h67 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h68 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h69 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h6a :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h6b :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h6c :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h6d :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h6e :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h6f :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h70 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h71 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h72 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h73 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h74 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h75 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h76 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h77 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h78 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h79 :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h7a :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h7b :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h7c :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h7d :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h7e :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	7'h7f :
		rl_a43_t8 = RG_quantized_block_rl_19 ;
	default :
		rl_a43_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_151 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a44_t8 = RG_rl_151 ;
	7'h01 :
		rl_a44_t8 = RG_rl_151 ;
	7'h02 :
		rl_a44_t8 = RG_rl_151 ;
	7'h03 :
		rl_a44_t8 = RG_rl_151 ;
	7'h04 :
		rl_a44_t8 = RG_rl_151 ;
	7'h05 :
		rl_a44_t8 = RG_rl_151 ;
	7'h06 :
		rl_a44_t8 = RG_rl_151 ;
	7'h07 :
		rl_a44_t8 = RG_rl_151 ;
	7'h08 :
		rl_a44_t8 = RG_rl_151 ;
	7'h09 :
		rl_a44_t8 = RG_rl_151 ;
	7'h0a :
		rl_a44_t8 = RG_rl_151 ;
	7'h0b :
		rl_a44_t8 = RG_rl_151 ;
	7'h0c :
		rl_a44_t8 = RG_rl_151 ;
	7'h0d :
		rl_a44_t8 = RG_rl_151 ;
	7'h0e :
		rl_a44_t8 = RG_rl_151 ;
	7'h0f :
		rl_a44_t8 = RG_rl_151 ;
	7'h10 :
		rl_a44_t8 = RG_rl_151 ;
	7'h11 :
		rl_a44_t8 = RG_rl_151 ;
	7'h12 :
		rl_a44_t8 = RG_rl_151 ;
	7'h13 :
		rl_a44_t8 = RG_rl_151 ;
	7'h14 :
		rl_a44_t8 = RG_rl_151 ;
	7'h15 :
		rl_a44_t8 = RG_rl_151 ;
	7'h16 :
		rl_a44_t8 = RG_rl_151 ;
	7'h17 :
		rl_a44_t8 = RG_rl_151 ;
	7'h18 :
		rl_a44_t8 = RG_rl_151 ;
	7'h19 :
		rl_a44_t8 = RG_rl_151 ;
	7'h1a :
		rl_a44_t8 = RG_rl_151 ;
	7'h1b :
		rl_a44_t8 = RG_rl_151 ;
	7'h1c :
		rl_a44_t8 = RG_rl_151 ;
	7'h1d :
		rl_a44_t8 = RG_rl_151 ;
	7'h1e :
		rl_a44_t8 = RG_rl_151 ;
	7'h1f :
		rl_a44_t8 = RG_rl_151 ;
	7'h20 :
		rl_a44_t8 = RG_rl_151 ;
	7'h21 :
		rl_a44_t8 = RG_rl_151 ;
	7'h22 :
		rl_a44_t8 = RG_rl_151 ;
	7'h23 :
		rl_a44_t8 = RG_rl_151 ;
	7'h24 :
		rl_a44_t8 = RG_rl_151 ;
	7'h25 :
		rl_a44_t8 = RG_rl_151 ;
	7'h26 :
		rl_a44_t8 = RG_rl_151 ;
	7'h27 :
		rl_a44_t8 = RG_rl_151 ;
	7'h28 :
		rl_a44_t8 = RG_rl_151 ;
	7'h29 :
		rl_a44_t8 = RG_rl_151 ;
	7'h2a :
		rl_a44_t8 = RG_rl_151 ;
	7'h2b :
		rl_a44_t8 = RG_rl_151 ;
	7'h2c :
		rl_a44_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h2d :
		rl_a44_t8 = RG_rl_151 ;
	7'h2e :
		rl_a44_t8 = RG_rl_151 ;
	7'h2f :
		rl_a44_t8 = RG_rl_151 ;
	7'h30 :
		rl_a44_t8 = RG_rl_151 ;
	7'h31 :
		rl_a44_t8 = RG_rl_151 ;
	7'h32 :
		rl_a44_t8 = RG_rl_151 ;
	7'h33 :
		rl_a44_t8 = RG_rl_151 ;
	7'h34 :
		rl_a44_t8 = RG_rl_151 ;
	7'h35 :
		rl_a44_t8 = RG_rl_151 ;
	7'h36 :
		rl_a44_t8 = RG_rl_151 ;
	7'h37 :
		rl_a44_t8 = RG_rl_151 ;
	7'h38 :
		rl_a44_t8 = RG_rl_151 ;
	7'h39 :
		rl_a44_t8 = RG_rl_151 ;
	7'h3a :
		rl_a44_t8 = RG_rl_151 ;
	7'h3b :
		rl_a44_t8 = RG_rl_151 ;
	7'h3c :
		rl_a44_t8 = RG_rl_151 ;
	7'h3d :
		rl_a44_t8 = RG_rl_151 ;
	7'h3e :
		rl_a44_t8 = RG_rl_151 ;
	7'h3f :
		rl_a44_t8 = RG_rl_151 ;
	7'h40 :
		rl_a44_t8 = RG_rl_151 ;
	7'h41 :
		rl_a44_t8 = RG_rl_151 ;
	7'h42 :
		rl_a44_t8 = RG_rl_151 ;
	7'h43 :
		rl_a44_t8 = RG_rl_151 ;
	7'h44 :
		rl_a44_t8 = RG_rl_151 ;
	7'h45 :
		rl_a44_t8 = RG_rl_151 ;
	7'h46 :
		rl_a44_t8 = RG_rl_151 ;
	7'h47 :
		rl_a44_t8 = RG_rl_151 ;
	7'h48 :
		rl_a44_t8 = RG_rl_151 ;
	7'h49 :
		rl_a44_t8 = RG_rl_151 ;
	7'h4a :
		rl_a44_t8 = RG_rl_151 ;
	7'h4b :
		rl_a44_t8 = RG_rl_151 ;
	7'h4c :
		rl_a44_t8 = RG_rl_151 ;
	7'h4d :
		rl_a44_t8 = RG_rl_151 ;
	7'h4e :
		rl_a44_t8 = RG_rl_151 ;
	7'h4f :
		rl_a44_t8 = RG_rl_151 ;
	7'h50 :
		rl_a44_t8 = RG_rl_151 ;
	7'h51 :
		rl_a44_t8 = RG_rl_151 ;
	7'h52 :
		rl_a44_t8 = RG_rl_151 ;
	7'h53 :
		rl_a44_t8 = RG_rl_151 ;
	7'h54 :
		rl_a44_t8 = RG_rl_151 ;
	7'h55 :
		rl_a44_t8 = RG_rl_151 ;
	7'h56 :
		rl_a44_t8 = RG_rl_151 ;
	7'h57 :
		rl_a44_t8 = RG_rl_151 ;
	7'h58 :
		rl_a44_t8 = RG_rl_151 ;
	7'h59 :
		rl_a44_t8 = RG_rl_151 ;
	7'h5a :
		rl_a44_t8 = RG_rl_151 ;
	7'h5b :
		rl_a44_t8 = RG_rl_151 ;
	7'h5c :
		rl_a44_t8 = RG_rl_151 ;
	7'h5d :
		rl_a44_t8 = RG_rl_151 ;
	7'h5e :
		rl_a44_t8 = RG_rl_151 ;
	7'h5f :
		rl_a44_t8 = RG_rl_151 ;
	7'h60 :
		rl_a44_t8 = RG_rl_151 ;
	7'h61 :
		rl_a44_t8 = RG_rl_151 ;
	7'h62 :
		rl_a44_t8 = RG_rl_151 ;
	7'h63 :
		rl_a44_t8 = RG_rl_151 ;
	7'h64 :
		rl_a44_t8 = RG_rl_151 ;
	7'h65 :
		rl_a44_t8 = RG_rl_151 ;
	7'h66 :
		rl_a44_t8 = RG_rl_151 ;
	7'h67 :
		rl_a44_t8 = RG_rl_151 ;
	7'h68 :
		rl_a44_t8 = RG_rl_151 ;
	7'h69 :
		rl_a44_t8 = RG_rl_151 ;
	7'h6a :
		rl_a44_t8 = RG_rl_151 ;
	7'h6b :
		rl_a44_t8 = RG_rl_151 ;
	7'h6c :
		rl_a44_t8 = RG_rl_151 ;
	7'h6d :
		rl_a44_t8 = RG_rl_151 ;
	7'h6e :
		rl_a44_t8 = RG_rl_151 ;
	7'h6f :
		rl_a44_t8 = RG_rl_151 ;
	7'h70 :
		rl_a44_t8 = RG_rl_151 ;
	7'h71 :
		rl_a44_t8 = RG_rl_151 ;
	7'h72 :
		rl_a44_t8 = RG_rl_151 ;
	7'h73 :
		rl_a44_t8 = RG_rl_151 ;
	7'h74 :
		rl_a44_t8 = RG_rl_151 ;
	7'h75 :
		rl_a44_t8 = RG_rl_151 ;
	7'h76 :
		rl_a44_t8 = RG_rl_151 ;
	7'h77 :
		rl_a44_t8 = RG_rl_151 ;
	7'h78 :
		rl_a44_t8 = RG_rl_151 ;
	7'h79 :
		rl_a44_t8 = RG_rl_151 ;
	7'h7a :
		rl_a44_t8 = RG_rl_151 ;
	7'h7b :
		rl_a44_t8 = RG_rl_151 ;
	7'h7c :
		rl_a44_t8 = RG_rl_151 ;
	7'h7d :
		rl_a44_t8 = RG_rl_151 ;
	7'h7e :
		rl_a44_t8 = RG_rl_151 ;
	7'h7f :
		rl_a44_t8 = RG_rl_151 ;
	default :
		rl_a44_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_20 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h01 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h02 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h03 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h04 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h05 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h06 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h07 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h08 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h09 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h0a :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h0b :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h0c :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h0d :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h0e :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h0f :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h10 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h11 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h12 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h13 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h14 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h15 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h16 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h17 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h18 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h19 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h1a :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h1b :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h1c :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h1d :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h1e :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h1f :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h20 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h21 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h22 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h23 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h24 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h25 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h26 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h27 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h28 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h29 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h2a :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h2b :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h2c :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h2d :
		rl_a45_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h2e :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h2f :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h30 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h31 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h32 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h33 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h34 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h35 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h36 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h37 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h38 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h39 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h3a :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h3b :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h3c :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h3d :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h3e :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h3f :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h40 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h41 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h42 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h43 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h44 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h45 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h46 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h47 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h48 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h49 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h4a :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h4b :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h4c :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h4d :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h4e :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h4f :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h50 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h51 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h52 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h53 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h54 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h55 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h56 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h57 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h58 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h59 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h5a :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h5b :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h5c :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h5d :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h5e :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h5f :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h60 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h61 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h62 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h63 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h64 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h65 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h66 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h67 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h68 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h69 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h6a :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h6b :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h6c :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h6d :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h6e :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h6f :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h70 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h71 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h72 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h73 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h74 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h75 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h76 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h77 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h78 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h79 :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h7a :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h7b :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h7c :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h7d :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h7e :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	7'h7f :
		rl_a45_t8 = RG_quantized_block_rl_20 ;
	default :
		rl_a45_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_152 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a46_t8 = RG_rl_152 ;
	7'h01 :
		rl_a46_t8 = RG_rl_152 ;
	7'h02 :
		rl_a46_t8 = RG_rl_152 ;
	7'h03 :
		rl_a46_t8 = RG_rl_152 ;
	7'h04 :
		rl_a46_t8 = RG_rl_152 ;
	7'h05 :
		rl_a46_t8 = RG_rl_152 ;
	7'h06 :
		rl_a46_t8 = RG_rl_152 ;
	7'h07 :
		rl_a46_t8 = RG_rl_152 ;
	7'h08 :
		rl_a46_t8 = RG_rl_152 ;
	7'h09 :
		rl_a46_t8 = RG_rl_152 ;
	7'h0a :
		rl_a46_t8 = RG_rl_152 ;
	7'h0b :
		rl_a46_t8 = RG_rl_152 ;
	7'h0c :
		rl_a46_t8 = RG_rl_152 ;
	7'h0d :
		rl_a46_t8 = RG_rl_152 ;
	7'h0e :
		rl_a46_t8 = RG_rl_152 ;
	7'h0f :
		rl_a46_t8 = RG_rl_152 ;
	7'h10 :
		rl_a46_t8 = RG_rl_152 ;
	7'h11 :
		rl_a46_t8 = RG_rl_152 ;
	7'h12 :
		rl_a46_t8 = RG_rl_152 ;
	7'h13 :
		rl_a46_t8 = RG_rl_152 ;
	7'h14 :
		rl_a46_t8 = RG_rl_152 ;
	7'h15 :
		rl_a46_t8 = RG_rl_152 ;
	7'h16 :
		rl_a46_t8 = RG_rl_152 ;
	7'h17 :
		rl_a46_t8 = RG_rl_152 ;
	7'h18 :
		rl_a46_t8 = RG_rl_152 ;
	7'h19 :
		rl_a46_t8 = RG_rl_152 ;
	7'h1a :
		rl_a46_t8 = RG_rl_152 ;
	7'h1b :
		rl_a46_t8 = RG_rl_152 ;
	7'h1c :
		rl_a46_t8 = RG_rl_152 ;
	7'h1d :
		rl_a46_t8 = RG_rl_152 ;
	7'h1e :
		rl_a46_t8 = RG_rl_152 ;
	7'h1f :
		rl_a46_t8 = RG_rl_152 ;
	7'h20 :
		rl_a46_t8 = RG_rl_152 ;
	7'h21 :
		rl_a46_t8 = RG_rl_152 ;
	7'h22 :
		rl_a46_t8 = RG_rl_152 ;
	7'h23 :
		rl_a46_t8 = RG_rl_152 ;
	7'h24 :
		rl_a46_t8 = RG_rl_152 ;
	7'h25 :
		rl_a46_t8 = RG_rl_152 ;
	7'h26 :
		rl_a46_t8 = RG_rl_152 ;
	7'h27 :
		rl_a46_t8 = RG_rl_152 ;
	7'h28 :
		rl_a46_t8 = RG_rl_152 ;
	7'h29 :
		rl_a46_t8 = RG_rl_152 ;
	7'h2a :
		rl_a46_t8 = RG_rl_152 ;
	7'h2b :
		rl_a46_t8 = RG_rl_152 ;
	7'h2c :
		rl_a46_t8 = RG_rl_152 ;
	7'h2d :
		rl_a46_t8 = RG_rl_152 ;
	7'h2e :
		rl_a46_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h2f :
		rl_a46_t8 = RG_rl_152 ;
	7'h30 :
		rl_a46_t8 = RG_rl_152 ;
	7'h31 :
		rl_a46_t8 = RG_rl_152 ;
	7'h32 :
		rl_a46_t8 = RG_rl_152 ;
	7'h33 :
		rl_a46_t8 = RG_rl_152 ;
	7'h34 :
		rl_a46_t8 = RG_rl_152 ;
	7'h35 :
		rl_a46_t8 = RG_rl_152 ;
	7'h36 :
		rl_a46_t8 = RG_rl_152 ;
	7'h37 :
		rl_a46_t8 = RG_rl_152 ;
	7'h38 :
		rl_a46_t8 = RG_rl_152 ;
	7'h39 :
		rl_a46_t8 = RG_rl_152 ;
	7'h3a :
		rl_a46_t8 = RG_rl_152 ;
	7'h3b :
		rl_a46_t8 = RG_rl_152 ;
	7'h3c :
		rl_a46_t8 = RG_rl_152 ;
	7'h3d :
		rl_a46_t8 = RG_rl_152 ;
	7'h3e :
		rl_a46_t8 = RG_rl_152 ;
	7'h3f :
		rl_a46_t8 = RG_rl_152 ;
	7'h40 :
		rl_a46_t8 = RG_rl_152 ;
	7'h41 :
		rl_a46_t8 = RG_rl_152 ;
	7'h42 :
		rl_a46_t8 = RG_rl_152 ;
	7'h43 :
		rl_a46_t8 = RG_rl_152 ;
	7'h44 :
		rl_a46_t8 = RG_rl_152 ;
	7'h45 :
		rl_a46_t8 = RG_rl_152 ;
	7'h46 :
		rl_a46_t8 = RG_rl_152 ;
	7'h47 :
		rl_a46_t8 = RG_rl_152 ;
	7'h48 :
		rl_a46_t8 = RG_rl_152 ;
	7'h49 :
		rl_a46_t8 = RG_rl_152 ;
	7'h4a :
		rl_a46_t8 = RG_rl_152 ;
	7'h4b :
		rl_a46_t8 = RG_rl_152 ;
	7'h4c :
		rl_a46_t8 = RG_rl_152 ;
	7'h4d :
		rl_a46_t8 = RG_rl_152 ;
	7'h4e :
		rl_a46_t8 = RG_rl_152 ;
	7'h4f :
		rl_a46_t8 = RG_rl_152 ;
	7'h50 :
		rl_a46_t8 = RG_rl_152 ;
	7'h51 :
		rl_a46_t8 = RG_rl_152 ;
	7'h52 :
		rl_a46_t8 = RG_rl_152 ;
	7'h53 :
		rl_a46_t8 = RG_rl_152 ;
	7'h54 :
		rl_a46_t8 = RG_rl_152 ;
	7'h55 :
		rl_a46_t8 = RG_rl_152 ;
	7'h56 :
		rl_a46_t8 = RG_rl_152 ;
	7'h57 :
		rl_a46_t8 = RG_rl_152 ;
	7'h58 :
		rl_a46_t8 = RG_rl_152 ;
	7'h59 :
		rl_a46_t8 = RG_rl_152 ;
	7'h5a :
		rl_a46_t8 = RG_rl_152 ;
	7'h5b :
		rl_a46_t8 = RG_rl_152 ;
	7'h5c :
		rl_a46_t8 = RG_rl_152 ;
	7'h5d :
		rl_a46_t8 = RG_rl_152 ;
	7'h5e :
		rl_a46_t8 = RG_rl_152 ;
	7'h5f :
		rl_a46_t8 = RG_rl_152 ;
	7'h60 :
		rl_a46_t8 = RG_rl_152 ;
	7'h61 :
		rl_a46_t8 = RG_rl_152 ;
	7'h62 :
		rl_a46_t8 = RG_rl_152 ;
	7'h63 :
		rl_a46_t8 = RG_rl_152 ;
	7'h64 :
		rl_a46_t8 = RG_rl_152 ;
	7'h65 :
		rl_a46_t8 = RG_rl_152 ;
	7'h66 :
		rl_a46_t8 = RG_rl_152 ;
	7'h67 :
		rl_a46_t8 = RG_rl_152 ;
	7'h68 :
		rl_a46_t8 = RG_rl_152 ;
	7'h69 :
		rl_a46_t8 = RG_rl_152 ;
	7'h6a :
		rl_a46_t8 = RG_rl_152 ;
	7'h6b :
		rl_a46_t8 = RG_rl_152 ;
	7'h6c :
		rl_a46_t8 = RG_rl_152 ;
	7'h6d :
		rl_a46_t8 = RG_rl_152 ;
	7'h6e :
		rl_a46_t8 = RG_rl_152 ;
	7'h6f :
		rl_a46_t8 = RG_rl_152 ;
	7'h70 :
		rl_a46_t8 = RG_rl_152 ;
	7'h71 :
		rl_a46_t8 = RG_rl_152 ;
	7'h72 :
		rl_a46_t8 = RG_rl_152 ;
	7'h73 :
		rl_a46_t8 = RG_rl_152 ;
	7'h74 :
		rl_a46_t8 = RG_rl_152 ;
	7'h75 :
		rl_a46_t8 = RG_rl_152 ;
	7'h76 :
		rl_a46_t8 = RG_rl_152 ;
	7'h77 :
		rl_a46_t8 = RG_rl_152 ;
	7'h78 :
		rl_a46_t8 = RG_rl_152 ;
	7'h79 :
		rl_a46_t8 = RG_rl_152 ;
	7'h7a :
		rl_a46_t8 = RG_rl_152 ;
	7'h7b :
		rl_a46_t8 = RG_rl_152 ;
	7'h7c :
		rl_a46_t8 = RG_rl_152 ;
	7'h7d :
		rl_a46_t8 = RG_rl_152 ;
	7'h7e :
		rl_a46_t8 = RG_rl_152 ;
	7'h7f :
		rl_a46_t8 = RG_rl_152 ;
	default :
		rl_a46_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_21 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h01 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h02 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h03 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h04 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h05 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h06 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h07 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h08 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h09 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h0a :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h0b :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h0c :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h0d :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h0e :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h0f :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h10 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h11 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h12 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h13 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h14 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h15 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h16 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h17 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h18 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h19 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h1a :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h1b :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h1c :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h1d :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h1e :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h1f :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h20 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h21 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h22 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h23 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h24 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h25 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h26 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h27 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h28 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h29 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h2a :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h2b :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h2c :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h2d :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h2e :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h2f :
		rl_a47_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h30 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h31 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h32 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h33 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h34 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h35 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h36 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h37 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h38 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h39 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h3a :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h3b :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h3c :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h3d :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h3e :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h3f :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h40 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h41 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h42 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h43 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h44 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h45 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h46 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h47 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h48 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h49 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h4a :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h4b :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h4c :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h4d :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h4e :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h4f :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h50 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h51 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h52 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h53 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h54 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h55 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h56 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h57 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h58 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h59 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h5a :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h5b :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h5c :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h5d :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h5e :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h5f :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h60 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h61 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h62 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h63 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h64 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h65 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h66 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h67 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h68 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h69 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h6a :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h6b :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h6c :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h6d :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h6e :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h6f :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h70 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h71 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h72 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h73 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h74 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h75 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h76 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h77 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h78 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h79 :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h7a :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h7b :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h7c :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h7d :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h7e :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	7'h7f :
		rl_a47_t8 = RG_quantized_block_rl_21 ;
	default :
		rl_a47_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_153 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a48_t8 = RG_rl_153 ;
	7'h01 :
		rl_a48_t8 = RG_rl_153 ;
	7'h02 :
		rl_a48_t8 = RG_rl_153 ;
	7'h03 :
		rl_a48_t8 = RG_rl_153 ;
	7'h04 :
		rl_a48_t8 = RG_rl_153 ;
	7'h05 :
		rl_a48_t8 = RG_rl_153 ;
	7'h06 :
		rl_a48_t8 = RG_rl_153 ;
	7'h07 :
		rl_a48_t8 = RG_rl_153 ;
	7'h08 :
		rl_a48_t8 = RG_rl_153 ;
	7'h09 :
		rl_a48_t8 = RG_rl_153 ;
	7'h0a :
		rl_a48_t8 = RG_rl_153 ;
	7'h0b :
		rl_a48_t8 = RG_rl_153 ;
	7'h0c :
		rl_a48_t8 = RG_rl_153 ;
	7'h0d :
		rl_a48_t8 = RG_rl_153 ;
	7'h0e :
		rl_a48_t8 = RG_rl_153 ;
	7'h0f :
		rl_a48_t8 = RG_rl_153 ;
	7'h10 :
		rl_a48_t8 = RG_rl_153 ;
	7'h11 :
		rl_a48_t8 = RG_rl_153 ;
	7'h12 :
		rl_a48_t8 = RG_rl_153 ;
	7'h13 :
		rl_a48_t8 = RG_rl_153 ;
	7'h14 :
		rl_a48_t8 = RG_rl_153 ;
	7'h15 :
		rl_a48_t8 = RG_rl_153 ;
	7'h16 :
		rl_a48_t8 = RG_rl_153 ;
	7'h17 :
		rl_a48_t8 = RG_rl_153 ;
	7'h18 :
		rl_a48_t8 = RG_rl_153 ;
	7'h19 :
		rl_a48_t8 = RG_rl_153 ;
	7'h1a :
		rl_a48_t8 = RG_rl_153 ;
	7'h1b :
		rl_a48_t8 = RG_rl_153 ;
	7'h1c :
		rl_a48_t8 = RG_rl_153 ;
	7'h1d :
		rl_a48_t8 = RG_rl_153 ;
	7'h1e :
		rl_a48_t8 = RG_rl_153 ;
	7'h1f :
		rl_a48_t8 = RG_rl_153 ;
	7'h20 :
		rl_a48_t8 = RG_rl_153 ;
	7'h21 :
		rl_a48_t8 = RG_rl_153 ;
	7'h22 :
		rl_a48_t8 = RG_rl_153 ;
	7'h23 :
		rl_a48_t8 = RG_rl_153 ;
	7'h24 :
		rl_a48_t8 = RG_rl_153 ;
	7'h25 :
		rl_a48_t8 = RG_rl_153 ;
	7'h26 :
		rl_a48_t8 = RG_rl_153 ;
	7'h27 :
		rl_a48_t8 = RG_rl_153 ;
	7'h28 :
		rl_a48_t8 = RG_rl_153 ;
	7'h29 :
		rl_a48_t8 = RG_rl_153 ;
	7'h2a :
		rl_a48_t8 = RG_rl_153 ;
	7'h2b :
		rl_a48_t8 = RG_rl_153 ;
	7'h2c :
		rl_a48_t8 = RG_rl_153 ;
	7'h2d :
		rl_a48_t8 = RG_rl_153 ;
	7'h2e :
		rl_a48_t8 = RG_rl_153 ;
	7'h2f :
		rl_a48_t8 = RG_rl_153 ;
	7'h30 :
		rl_a48_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h31 :
		rl_a48_t8 = RG_rl_153 ;
	7'h32 :
		rl_a48_t8 = RG_rl_153 ;
	7'h33 :
		rl_a48_t8 = RG_rl_153 ;
	7'h34 :
		rl_a48_t8 = RG_rl_153 ;
	7'h35 :
		rl_a48_t8 = RG_rl_153 ;
	7'h36 :
		rl_a48_t8 = RG_rl_153 ;
	7'h37 :
		rl_a48_t8 = RG_rl_153 ;
	7'h38 :
		rl_a48_t8 = RG_rl_153 ;
	7'h39 :
		rl_a48_t8 = RG_rl_153 ;
	7'h3a :
		rl_a48_t8 = RG_rl_153 ;
	7'h3b :
		rl_a48_t8 = RG_rl_153 ;
	7'h3c :
		rl_a48_t8 = RG_rl_153 ;
	7'h3d :
		rl_a48_t8 = RG_rl_153 ;
	7'h3e :
		rl_a48_t8 = RG_rl_153 ;
	7'h3f :
		rl_a48_t8 = RG_rl_153 ;
	7'h40 :
		rl_a48_t8 = RG_rl_153 ;
	7'h41 :
		rl_a48_t8 = RG_rl_153 ;
	7'h42 :
		rl_a48_t8 = RG_rl_153 ;
	7'h43 :
		rl_a48_t8 = RG_rl_153 ;
	7'h44 :
		rl_a48_t8 = RG_rl_153 ;
	7'h45 :
		rl_a48_t8 = RG_rl_153 ;
	7'h46 :
		rl_a48_t8 = RG_rl_153 ;
	7'h47 :
		rl_a48_t8 = RG_rl_153 ;
	7'h48 :
		rl_a48_t8 = RG_rl_153 ;
	7'h49 :
		rl_a48_t8 = RG_rl_153 ;
	7'h4a :
		rl_a48_t8 = RG_rl_153 ;
	7'h4b :
		rl_a48_t8 = RG_rl_153 ;
	7'h4c :
		rl_a48_t8 = RG_rl_153 ;
	7'h4d :
		rl_a48_t8 = RG_rl_153 ;
	7'h4e :
		rl_a48_t8 = RG_rl_153 ;
	7'h4f :
		rl_a48_t8 = RG_rl_153 ;
	7'h50 :
		rl_a48_t8 = RG_rl_153 ;
	7'h51 :
		rl_a48_t8 = RG_rl_153 ;
	7'h52 :
		rl_a48_t8 = RG_rl_153 ;
	7'h53 :
		rl_a48_t8 = RG_rl_153 ;
	7'h54 :
		rl_a48_t8 = RG_rl_153 ;
	7'h55 :
		rl_a48_t8 = RG_rl_153 ;
	7'h56 :
		rl_a48_t8 = RG_rl_153 ;
	7'h57 :
		rl_a48_t8 = RG_rl_153 ;
	7'h58 :
		rl_a48_t8 = RG_rl_153 ;
	7'h59 :
		rl_a48_t8 = RG_rl_153 ;
	7'h5a :
		rl_a48_t8 = RG_rl_153 ;
	7'h5b :
		rl_a48_t8 = RG_rl_153 ;
	7'h5c :
		rl_a48_t8 = RG_rl_153 ;
	7'h5d :
		rl_a48_t8 = RG_rl_153 ;
	7'h5e :
		rl_a48_t8 = RG_rl_153 ;
	7'h5f :
		rl_a48_t8 = RG_rl_153 ;
	7'h60 :
		rl_a48_t8 = RG_rl_153 ;
	7'h61 :
		rl_a48_t8 = RG_rl_153 ;
	7'h62 :
		rl_a48_t8 = RG_rl_153 ;
	7'h63 :
		rl_a48_t8 = RG_rl_153 ;
	7'h64 :
		rl_a48_t8 = RG_rl_153 ;
	7'h65 :
		rl_a48_t8 = RG_rl_153 ;
	7'h66 :
		rl_a48_t8 = RG_rl_153 ;
	7'h67 :
		rl_a48_t8 = RG_rl_153 ;
	7'h68 :
		rl_a48_t8 = RG_rl_153 ;
	7'h69 :
		rl_a48_t8 = RG_rl_153 ;
	7'h6a :
		rl_a48_t8 = RG_rl_153 ;
	7'h6b :
		rl_a48_t8 = RG_rl_153 ;
	7'h6c :
		rl_a48_t8 = RG_rl_153 ;
	7'h6d :
		rl_a48_t8 = RG_rl_153 ;
	7'h6e :
		rl_a48_t8 = RG_rl_153 ;
	7'h6f :
		rl_a48_t8 = RG_rl_153 ;
	7'h70 :
		rl_a48_t8 = RG_rl_153 ;
	7'h71 :
		rl_a48_t8 = RG_rl_153 ;
	7'h72 :
		rl_a48_t8 = RG_rl_153 ;
	7'h73 :
		rl_a48_t8 = RG_rl_153 ;
	7'h74 :
		rl_a48_t8 = RG_rl_153 ;
	7'h75 :
		rl_a48_t8 = RG_rl_153 ;
	7'h76 :
		rl_a48_t8 = RG_rl_153 ;
	7'h77 :
		rl_a48_t8 = RG_rl_153 ;
	7'h78 :
		rl_a48_t8 = RG_rl_153 ;
	7'h79 :
		rl_a48_t8 = RG_rl_153 ;
	7'h7a :
		rl_a48_t8 = RG_rl_153 ;
	7'h7b :
		rl_a48_t8 = RG_rl_153 ;
	7'h7c :
		rl_a48_t8 = RG_rl_153 ;
	7'h7d :
		rl_a48_t8 = RG_rl_153 ;
	7'h7e :
		rl_a48_t8 = RG_rl_153 ;
	7'h7f :
		rl_a48_t8 = RG_rl_153 ;
	default :
		rl_a48_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_22 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h01 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h02 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h03 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h04 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h05 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h06 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h07 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h08 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h09 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h0a :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h0b :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h0c :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h0d :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h0e :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h0f :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h10 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h11 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h12 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h13 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h14 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h15 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h16 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h17 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h18 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h19 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h1a :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h1b :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h1c :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h1d :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h1e :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h1f :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h20 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h21 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h22 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h23 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h24 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h25 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h26 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h27 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h28 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h29 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h2a :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h2b :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h2c :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h2d :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h2e :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h2f :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h30 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h31 :
		rl_a49_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h32 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h33 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h34 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h35 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h36 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h37 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h38 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h39 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h3a :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h3b :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h3c :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h3d :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h3e :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h3f :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h40 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h41 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h42 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h43 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h44 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h45 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h46 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h47 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h48 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h49 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h4a :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h4b :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h4c :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h4d :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h4e :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h4f :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h50 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h51 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h52 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h53 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h54 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h55 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h56 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h57 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h58 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h59 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h5a :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h5b :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h5c :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h5d :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h5e :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h5f :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h60 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h61 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h62 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h63 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h64 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h65 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h66 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h67 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h68 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h69 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h6a :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h6b :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h6c :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h6d :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h6e :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h6f :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h70 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h71 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h72 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h73 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h74 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h75 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h76 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h77 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h78 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h79 :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h7a :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h7b :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h7c :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h7d :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h7e :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	7'h7f :
		rl_a49_t8 = RG_quantized_block_rl_22 ;
	default :
		rl_a49_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_154 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a50_t8 = RG_rl_154 ;
	7'h01 :
		rl_a50_t8 = RG_rl_154 ;
	7'h02 :
		rl_a50_t8 = RG_rl_154 ;
	7'h03 :
		rl_a50_t8 = RG_rl_154 ;
	7'h04 :
		rl_a50_t8 = RG_rl_154 ;
	7'h05 :
		rl_a50_t8 = RG_rl_154 ;
	7'h06 :
		rl_a50_t8 = RG_rl_154 ;
	7'h07 :
		rl_a50_t8 = RG_rl_154 ;
	7'h08 :
		rl_a50_t8 = RG_rl_154 ;
	7'h09 :
		rl_a50_t8 = RG_rl_154 ;
	7'h0a :
		rl_a50_t8 = RG_rl_154 ;
	7'h0b :
		rl_a50_t8 = RG_rl_154 ;
	7'h0c :
		rl_a50_t8 = RG_rl_154 ;
	7'h0d :
		rl_a50_t8 = RG_rl_154 ;
	7'h0e :
		rl_a50_t8 = RG_rl_154 ;
	7'h0f :
		rl_a50_t8 = RG_rl_154 ;
	7'h10 :
		rl_a50_t8 = RG_rl_154 ;
	7'h11 :
		rl_a50_t8 = RG_rl_154 ;
	7'h12 :
		rl_a50_t8 = RG_rl_154 ;
	7'h13 :
		rl_a50_t8 = RG_rl_154 ;
	7'h14 :
		rl_a50_t8 = RG_rl_154 ;
	7'h15 :
		rl_a50_t8 = RG_rl_154 ;
	7'h16 :
		rl_a50_t8 = RG_rl_154 ;
	7'h17 :
		rl_a50_t8 = RG_rl_154 ;
	7'h18 :
		rl_a50_t8 = RG_rl_154 ;
	7'h19 :
		rl_a50_t8 = RG_rl_154 ;
	7'h1a :
		rl_a50_t8 = RG_rl_154 ;
	7'h1b :
		rl_a50_t8 = RG_rl_154 ;
	7'h1c :
		rl_a50_t8 = RG_rl_154 ;
	7'h1d :
		rl_a50_t8 = RG_rl_154 ;
	7'h1e :
		rl_a50_t8 = RG_rl_154 ;
	7'h1f :
		rl_a50_t8 = RG_rl_154 ;
	7'h20 :
		rl_a50_t8 = RG_rl_154 ;
	7'h21 :
		rl_a50_t8 = RG_rl_154 ;
	7'h22 :
		rl_a50_t8 = RG_rl_154 ;
	7'h23 :
		rl_a50_t8 = RG_rl_154 ;
	7'h24 :
		rl_a50_t8 = RG_rl_154 ;
	7'h25 :
		rl_a50_t8 = RG_rl_154 ;
	7'h26 :
		rl_a50_t8 = RG_rl_154 ;
	7'h27 :
		rl_a50_t8 = RG_rl_154 ;
	7'h28 :
		rl_a50_t8 = RG_rl_154 ;
	7'h29 :
		rl_a50_t8 = RG_rl_154 ;
	7'h2a :
		rl_a50_t8 = RG_rl_154 ;
	7'h2b :
		rl_a50_t8 = RG_rl_154 ;
	7'h2c :
		rl_a50_t8 = RG_rl_154 ;
	7'h2d :
		rl_a50_t8 = RG_rl_154 ;
	7'h2e :
		rl_a50_t8 = RG_rl_154 ;
	7'h2f :
		rl_a50_t8 = RG_rl_154 ;
	7'h30 :
		rl_a50_t8 = RG_rl_154 ;
	7'h31 :
		rl_a50_t8 = RG_rl_154 ;
	7'h32 :
		rl_a50_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h33 :
		rl_a50_t8 = RG_rl_154 ;
	7'h34 :
		rl_a50_t8 = RG_rl_154 ;
	7'h35 :
		rl_a50_t8 = RG_rl_154 ;
	7'h36 :
		rl_a50_t8 = RG_rl_154 ;
	7'h37 :
		rl_a50_t8 = RG_rl_154 ;
	7'h38 :
		rl_a50_t8 = RG_rl_154 ;
	7'h39 :
		rl_a50_t8 = RG_rl_154 ;
	7'h3a :
		rl_a50_t8 = RG_rl_154 ;
	7'h3b :
		rl_a50_t8 = RG_rl_154 ;
	7'h3c :
		rl_a50_t8 = RG_rl_154 ;
	7'h3d :
		rl_a50_t8 = RG_rl_154 ;
	7'h3e :
		rl_a50_t8 = RG_rl_154 ;
	7'h3f :
		rl_a50_t8 = RG_rl_154 ;
	7'h40 :
		rl_a50_t8 = RG_rl_154 ;
	7'h41 :
		rl_a50_t8 = RG_rl_154 ;
	7'h42 :
		rl_a50_t8 = RG_rl_154 ;
	7'h43 :
		rl_a50_t8 = RG_rl_154 ;
	7'h44 :
		rl_a50_t8 = RG_rl_154 ;
	7'h45 :
		rl_a50_t8 = RG_rl_154 ;
	7'h46 :
		rl_a50_t8 = RG_rl_154 ;
	7'h47 :
		rl_a50_t8 = RG_rl_154 ;
	7'h48 :
		rl_a50_t8 = RG_rl_154 ;
	7'h49 :
		rl_a50_t8 = RG_rl_154 ;
	7'h4a :
		rl_a50_t8 = RG_rl_154 ;
	7'h4b :
		rl_a50_t8 = RG_rl_154 ;
	7'h4c :
		rl_a50_t8 = RG_rl_154 ;
	7'h4d :
		rl_a50_t8 = RG_rl_154 ;
	7'h4e :
		rl_a50_t8 = RG_rl_154 ;
	7'h4f :
		rl_a50_t8 = RG_rl_154 ;
	7'h50 :
		rl_a50_t8 = RG_rl_154 ;
	7'h51 :
		rl_a50_t8 = RG_rl_154 ;
	7'h52 :
		rl_a50_t8 = RG_rl_154 ;
	7'h53 :
		rl_a50_t8 = RG_rl_154 ;
	7'h54 :
		rl_a50_t8 = RG_rl_154 ;
	7'h55 :
		rl_a50_t8 = RG_rl_154 ;
	7'h56 :
		rl_a50_t8 = RG_rl_154 ;
	7'h57 :
		rl_a50_t8 = RG_rl_154 ;
	7'h58 :
		rl_a50_t8 = RG_rl_154 ;
	7'h59 :
		rl_a50_t8 = RG_rl_154 ;
	7'h5a :
		rl_a50_t8 = RG_rl_154 ;
	7'h5b :
		rl_a50_t8 = RG_rl_154 ;
	7'h5c :
		rl_a50_t8 = RG_rl_154 ;
	7'h5d :
		rl_a50_t8 = RG_rl_154 ;
	7'h5e :
		rl_a50_t8 = RG_rl_154 ;
	7'h5f :
		rl_a50_t8 = RG_rl_154 ;
	7'h60 :
		rl_a50_t8 = RG_rl_154 ;
	7'h61 :
		rl_a50_t8 = RG_rl_154 ;
	7'h62 :
		rl_a50_t8 = RG_rl_154 ;
	7'h63 :
		rl_a50_t8 = RG_rl_154 ;
	7'h64 :
		rl_a50_t8 = RG_rl_154 ;
	7'h65 :
		rl_a50_t8 = RG_rl_154 ;
	7'h66 :
		rl_a50_t8 = RG_rl_154 ;
	7'h67 :
		rl_a50_t8 = RG_rl_154 ;
	7'h68 :
		rl_a50_t8 = RG_rl_154 ;
	7'h69 :
		rl_a50_t8 = RG_rl_154 ;
	7'h6a :
		rl_a50_t8 = RG_rl_154 ;
	7'h6b :
		rl_a50_t8 = RG_rl_154 ;
	7'h6c :
		rl_a50_t8 = RG_rl_154 ;
	7'h6d :
		rl_a50_t8 = RG_rl_154 ;
	7'h6e :
		rl_a50_t8 = RG_rl_154 ;
	7'h6f :
		rl_a50_t8 = RG_rl_154 ;
	7'h70 :
		rl_a50_t8 = RG_rl_154 ;
	7'h71 :
		rl_a50_t8 = RG_rl_154 ;
	7'h72 :
		rl_a50_t8 = RG_rl_154 ;
	7'h73 :
		rl_a50_t8 = RG_rl_154 ;
	7'h74 :
		rl_a50_t8 = RG_rl_154 ;
	7'h75 :
		rl_a50_t8 = RG_rl_154 ;
	7'h76 :
		rl_a50_t8 = RG_rl_154 ;
	7'h77 :
		rl_a50_t8 = RG_rl_154 ;
	7'h78 :
		rl_a50_t8 = RG_rl_154 ;
	7'h79 :
		rl_a50_t8 = RG_rl_154 ;
	7'h7a :
		rl_a50_t8 = RG_rl_154 ;
	7'h7b :
		rl_a50_t8 = RG_rl_154 ;
	7'h7c :
		rl_a50_t8 = RG_rl_154 ;
	7'h7d :
		rl_a50_t8 = RG_rl_154 ;
	7'h7e :
		rl_a50_t8 = RG_rl_154 ;
	7'h7f :
		rl_a50_t8 = RG_rl_154 ;
	default :
		rl_a50_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_23 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h01 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h02 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h03 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h04 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h05 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h06 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h07 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h08 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h09 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h0a :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h0b :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h0c :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h0d :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h0e :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h0f :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h10 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h11 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h12 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h13 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h14 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h15 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h16 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h17 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h18 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h19 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h1a :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h1b :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h1c :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h1d :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h1e :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h1f :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h20 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h21 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h22 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h23 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h24 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h25 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h26 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h27 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h28 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h29 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h2a :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h2b :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h2c :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h2d :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h2e :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h2f :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h30 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h31 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h32 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h33 :
		rl_a51_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h34 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h35 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h36 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h37 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h38 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h39 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h3a :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h3b :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h3c :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h3d :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h3e :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h3f :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h40 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h41 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h42 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h43 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h44 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h45 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h46 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h47 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h48 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h49 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h4a :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h4b :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h4c :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h4d :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h4e :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h4f :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h50 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h51 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h52 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h53 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h54 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h55 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h56 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h57 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h58 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h59 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h5a :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h5b :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h5c :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h5d :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h5e :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h5f :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h60 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h61 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h62 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h63 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h64 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h65 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h66 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h67 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h68 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h69 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h6a :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h6b :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h6c :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h6d :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h6e :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h6f :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h70 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h71 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h72 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h73 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h74 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h75 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h76 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h77 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h78 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h79 :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h7a :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h7b :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h7c :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h7d :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h7e :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	7'h7f :
		rl_a51_t8 = RG_quantized_block_rl_23 ;
	default :
		rl_a51_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_155 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a52_t8 = RG_rl_155 ;
	7'h01 :
		rl_a52_t8 = RG_rl_155 ;
	7'h02 :
		rl_a52_t8 = RG_rl_155 ;
	7'h03 :
		rl_a52_t8 = RG_rl_155 ;
	7'h04 :
		rl_a52_t8 = RG_rl_155 ;
	7'h05 :
		rl_a52_t8 = RG_rl_155 ;
	7'h06 :
		rl_a52_t8 = RG_rl_155 ;
	7'h07 :
		rl_a52_t8 = RG_rl_155 ;
	7'h08 :
		rl_a52_t8 = RG_rl_155 ;
	7'h09 :
		rl_a52_t8 = RG_rl_155 ;
	7'h0a :
		rl_a52_t8 = RG_rl_155 ;
	7'h0b :
		rl_a52_t8 = RG_rl_155 ;
	7'h0c :
		rl_a52_t8 = RG_rl_155 ;
	7'h0d :
		rl_a52_t8 = RG_rl_155 ;
	7'h0e :
		rl_a52_t8 = RG_rl_155 ;
	7'h0f :
		rl_a52_t8 = RG_rl_155 ;
	7'h10 :
		rl_a52_t8 = RG_rl_155 ;
	7'h11 :
		rl_a52_t8 = RG_rl_155 ;
	7'h12 :
		rl_a52_t8 = RG_rl_155 ;
	7'h13 :
		rl_a52_t8 = RG_rl_155 ;
	7'h14 :
		rl_a52_t8 = RG_rl_155 ;
	7'h15 :
		rl_a52_t8 = RG_rl_155 ;
	7'h16 :
		rl_a52_t8 = RG_rl_155 ;
	7'h17 :
		rl_a52_t8 = RG_rl_155 ;
	7'h18 :
		rl_a52_t8 = RG_rl_155 ;
	7'h19 :
		rl_a52_t8 = RG_rl_155 ;
	7'h1a :
		rl_a52_t8 = RG_rl_155 ;
	7'h1b :
		rl_a52_t8 = RG_rl_155 ;
	7'h1c :
		rl_a52_t8 = RG_rl_155 ;
	7'h1d :
		rl_a52_t8 = RG_rl_155 ;
	7'h1e :
		rl_a52_t8 = RG_rl_155 ;
	7'h1f :
		rl_a52_t8 = RG_rl_155 ;
	7'h20 :
		rl_a52_t8 = RG_rl_155 ;
	7'h21 :
		rl_a52_t8 = RG_rl_155 ;
	7'h22 :
		rl_a52_t8 = RG_rl_155 ;
	7'h23 :
		rl_a52_t8 = RG_rl_155 ;
	7'h24 :
		rl_a52_t8 = RG_rl_155 ;
	7'h25 :
		rl_a52_t8 = RG_rl_155 ;
	7'h26 :
		rl_a52_t8 = RG_rl_155 ;
	7'h27 :
		rl_a52_t8 = RG_rl_155 ;
	7'h28 :
		rl_a52_t8 = RG_rl_155 ;
	7'h29 :
		rl_a52_t8 = RG_rl_155 ;
	7'h2a :
		rl_a52_t8 = RG_rl_155 ;
	7'h2b :
		rl_a52_t8 = RG_rl_155 ;
	7'h2c :
		rl_a52_t8 = RG_rl_155 ;
	7'h2d :
		rl_a52_t8 = RG_rl_155 ;
	7'h2e :
		rl_a52_t8 = RG_rl_155 ;
	7'h2f :
		rl_a52_t8 = RG_rl_155 ;
	7'h30 :
		rl_a52_t8 = RG_rl_155 ;
	7'h31 :
		rl_a52_t8 = RG_rl_155 ;
	7'h32 :
		rl_a52_t8 = RG_rl_155 ;
	7'h33 :
		rl_a52_t8 = RG_rl_155 ;
	7'h34 :
		rl_a52_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h35 :
		rl_a52_t8 = RG_rl_155 ;
	7'h36 :
		rl_a52_t8 = RG_rl_155 ;
	7'h37 :
		rl_a52_t8 = RG_rl_155 ;
	7'h38 :
		rl_a52_t8 = RG_rl_155 ;
	7'h39 :
		rl_a52_t8 = RG_rl_155 ;
	7'h3a :
		rl_a52_t8 = RG_rl_155 ;
	7'h3b :
		rl_a52_t8 = RG_rl_155 ;
	7'h3c :
		rl_a52_t8 = RG_rl_155 ;
	7'h3d :
		rl_a52_t8 = RG_rl_155 ;
	7'h3e :
		rl_a52_t8 = RG_rl_155 ;
	7'h3f :
		rl_a52_t8 = RG_rl_155 ;
	7'h40 :
		rl_a52_t8 = RG_rl_155 ;
	7'h41 :
		rl_a52_t8 = RG_rl_155 ;
	7'h42 :
		rl_a52_t8 = RG_rl_155 ;
	7'h43 :
		rl_a52_t8 = RG_rl_155 ;
	7'h44 :
		rl_a52_t8 = RG_rl_155 ;
	7'h45 :
		rl_a52_t8 = RG_rl_155 ;
	7'h46 :
		rl_a52_t8 = RG_rl_155 ;
	7'h47 :
		rl_a52_t8 = RG_rl_155 ;
	7'h48 :
		rl_a52_t8 = RG_rl_155 ;
	7'h49 :
		rl_a52_t8 = RG_rl_155 ;
	7'h4a :
		rl_a52_t8 = RG_rl_155 ;
	7'h4b :
		rl_a52_t8 = RG_rl_155 ;
	7'h4c :
		rl_a52_t8 = RG_rl_155 ;
	7'h4d :
		rl_a52_t8 = RG_rl_155 ;
	7'h4e :
		rl_a52_t8 = RG_rl_155 ;
	7'h4f :
		rl_a52_t8 = RG_rl_155 ;
	7'h50 :
		rl_a52_t8 = RG_rl_155 ;
	7'h51 :
		rl_a52_t8 = RG_rl_155 ;
	7'h52 :
		rl_a52_t8 = RG_rl_155 ;
	7'h53 :
		rl_a52_t8 = RG_rl_155 ;
	7'h54 :
		rl_a52_t8 = RG_rl_155 ;
	7'h55 :
		rl_a52_t8 = RG_rl_155 ;
	7'h56 :
		rl_a52_t8 = RG_rl_155 ;
	7'h57 :
		rl_a52_t8 = RG_rl_155 ;
	7'h58 :
		rl_a52_t8 = RG_rl_155 ;
	7'h59 :
		rl_a52_t8 = RG_rl_155 ;
	7'h5a :
		rl_a52_t8 = RG_rl_155 ;
	7'h5b :
		rl_a52_t8 = RG_rl_155 ;
	7'h5c :
		rl_a52_t8 = RG_rl_155 ;
	7'h5d :
		rl_a52_t8 = RG_rl_155 ;
	7'h5e :
		rl_a52_t8 = RG_rl_155 ;
	7'h5f :
		rl_a52_t8 = RG_rl_155 ;
	7'h60 :
		rl_a52_t8 = RG_rl_155 ;
	7'h61 :
		rl_a52_t8 = RG_rl_155 ;
	7'h62 :
		rl_a52_t8 = RG_rl_155 ;
	7'h63 :
		rl_a52_t8 = RG_rl_155 ;
	7'h64 :
		rl_a52_t8 = RG_rl_155 ;
	7'h65 :
		rl_a52_t8 = RG_rl_155 ;
	7'h66 :
		rl_a52_t8 = RG_rl_155 ;
	7'h67 :
		rl_a52_t8 = RG_rl_155 ;
	7'h68 :
		rl_a52_t8 = RG_rl_155 ;
	7'h69 :
		rl_a52_t8 = RG_rl_155 ;
	7'h6a :
		rl_a52_t8 = RG_rl_155 ;
	7'h6b :
		rl_a52_t8 = RG_rl_155 ;
	7'h6c :
		rl_a52_t8 = RG_rl_155 ;
	7'h6d :
		rl_a52_t8 = RG_rl_155 ;
	7'h6e :
		rl_a52_t8 = RG_rl_155 ;
	7'h6f :
		rl_a52_t8 = RG_rl_155 ;
	7'h70 :
		rl_a52_t8 = RG_rl_155 ;
	7'h71 :
		rl_a52_t8 = RG_rl_155 ;
	7'h72 :
		rl_a52_t8 = RG_rl_155 ;
	7'h73 :
		rl_a52_t8 = RG_rl_155 ;
	7'h74 :
		rl_a52_t8 = RG_rl_155 ;
	7'h75 :
		rl_a52_t8 = RG_rl_155 ;
	7'h76 :
		rl_a52_t8 = RG_rl_155 ;
	7'h77 :
		rl_a52_t8 = RG_rl_155 ;
	7'h78 :
		rl_a52_t8 = RG_rl_155 ;
	7'h79 :
		rl_a52_t8 = RG_rl_155 ;
	7'h7a :
		rl_a52_t8 = RG_rl_155 ;
	7'h7b :
		rl_a52_t8 = RG_rl_155 ;
	7'h7c :
		rl_a52_t8 = RG_rl_155 ;
	7'h7d :
		rl_a52_t8 = RG_rl_155 ;
	7'h7e :
		rl_a52_t8 = RG_rl_155 ;
	7'h7f :
		rl_a52_t8 = RG_rl_155 ;
	default :
		rl_a52_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_24 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h01 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h02 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h03 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h04 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h05 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h06 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h07 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h08 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h09 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h0a :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h0b :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h0c :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h0d :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h0e :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h0f :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h10 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h11 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h12 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h13 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h14 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h15 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h16 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h17 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h18 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h19 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h1a :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h1b :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h1c :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h1d :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h1e :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h1f :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h20 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h21 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h22 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h23 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h24 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h25 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h26 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h27 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h28 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h29 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h2a :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h2b :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h2c :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h2d :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h2e :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h2f :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h30 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h31 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h32 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h33 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h34 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h35 :
		rl_a53_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h36 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h37 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h38 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h39 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h3a :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h3b :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h3c :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h3d :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h3e :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h3f :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h40 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h41 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h42 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h43 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h44 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h45 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h46 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h47 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h48 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h49 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h4a :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h4b :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h4c :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h4d :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h4e :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h4f :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h50 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h51 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h52 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h53 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h54 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h55 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h56 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h57 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h58 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h59 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h5a :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h5b :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h5c :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h5d :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h5e :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h5f :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h60 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h61 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h62 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h63 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h64 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h65 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h66 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h67 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h68 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h69 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h6a :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h6b :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h6c :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h6d :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h6e :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h6f :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h70 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h71 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h72 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h73 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h74 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h75 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h76 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h77 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h78 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h79 :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h7a :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h7b :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h7c :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h7d :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h7e :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	7'h7f :
		rl_a53_t8 = RG_quantized_block_rl_24 ;
	default :
		rl_a53_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_156 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a54_t8 = RG_rl_156 ;
	7'h01 :
		rl_a54_t8 = RG_rl_156 ;
	7'h02 :
		rl_a54_t8 = RG_rl_156 ;
	7'h03 :
		rl_a54_t8 = RG_rl_156 ;
	7'h04 :
		rl_a54_t8 = RG_rl_156 ;
	7'h05 :
		rl_a54_t8 = RG_rl_156 ;
	7'h06 :
		rl_a54_t8 = RG_rl_156 ;
	7'h07 :
		rl_a54_t8 = RG_rl_156 ;
	7'h08 :
		rl_a54_t8 = RG_rl_156 ;
	7'h09 :
		rl_a54_t8 = RG_rl_156 ;
	7'h0a :
		rl_a54_t8 = RG_rl_156 ;
	7'h0b :
		rl_a54_t8 = RG_rl_156 ;
	7'h0c :
		rl_a54_t8 = RG_rl_156 ;
	7'h0d :
		rl_a54_t8 = RG_rl_156 ;
	7'h0e :
		rl_a54_t8 = RG_rl_156 ;
	7'h0f :
		rl_a54_t8 = RG_rl_156 ;
	7'h10 :
		rl_a54_t8 = RG_rl_156 ;
	7'h11 :
		rl_a54_t8 = RG_rl_156 ;
	7'h12 :
		rl_a54_t8 = RG_rl_156 ;
	7'h13 :
		rl_a54_t8 = RG_rl_156 ;
	7'h14 :
		rl_a54_t8 = RG_rl_156 ;
	7'h15 :
		rl_a54_t8 = RG_rl_156 ;
	7'h16 :
		rl_a54_t8 = RG_rl_156 ;
	7'h17 :
		rl_a54_t8 = RG_rl_156 ;
	7'h18 :
		rl_a54_t8 = RG_rl_156 ;
	7'h19 :
		rl_a54_t8 = RG_rl_156 ;
	7'h1a :
		rl_a54_t8 = RG_rl_156 ;
	7'h1b :
		rl_a54_t8 = RG_rl_156 ;
	7'h1c :
		rl_a54_t8 = RG_rl_156 ;
	7'h1d :
		rl_a54_t8 = RG_rl_156 ;
	7'h1e :
		rl_a54_t8 = RG_rl_156 ;
	7'h1f :
		rl_a54_t8 = RG_rl_156 ;
	7'h20 :
		rl_a54_t8 = RG_rl_156 ;
	7'h21 :
		rl_a54_t8 = RG_rl_156 ;
	7'h22 :
		rl_a54_t8 = RG_rl_156 ;
	7'h23 :
		rl_a54_t8 = RG_rl_156 ;
	7'h24 :
		rl_a54_t8 = RG_rl_156 ;
	7'h25 :
		rl_a54_t8 = RG_rl_156 ;
	7'h26 :
		rl_a54_t8 = RG_rl_156 ;
	7'h27 :
		rl_a54_t8 = RG_rl_156 ;
	7'h28 :
		rl_a54_t8 = RG_rl_156 ;
	7'h29 :
		rl_a54_t8 = RG_rl_156 ;
	7'h2a :
		rl_a54_t8 = RG_rl_156 ;
	7'h2b :
		rl_a54_t8 = RG_rl_156 ;
	7'h2c :
		rl_a54_t8 = RG_rl_156 ;
	7'h2d :
		rl_a54_t8 = RG_rl_156 ;
	7'h2e :
		rl_a54_t8 = RG_rl_156 ;
	7'h2f :
		rl_a54_t8 = RG_rl_156 ;
	7'h30 :
		rl_a54_t8 = RG_rl_156 ;
	7'h31 :
		rl_a54_t8 = RG_rl_156 ;
	7'h32 :
		rl_a54_t8 = RG_rl_156 ;
	7'h33 :
		rl_a54_t8 = RG_rl_156 ;
	7'h34 :
		rl_a54_t8 = RG_rl_156 ;
	7'h35 :
		rl_a54_t8 = RG_rl_156 ;
	7'h36 :
		rl_a54_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h37 :
		rl_a54_t8 = RG_rl_156 ;
	7'h38 :
		rl_a54_t8 = RG_rl_156 ;
	7'h39 :
		rl_a54_t8 = RG_rl_156 ;
	7'h3a :
		rl_a54_t8 = RG_rl_156 ;
	7'h3b :
		rl_a54_t8 = RG_rl_156 ;
	7'h3c :
		rl_a54_t8 = RG_rl_156 ;
	7'h3d :
		rl_a54_t8 = RG_rl_156 ;
	7'h3e :
		rl_a54_t8 = RG_rl_156 ;
	7'h3f :
		rl_a54_t8 = RG_rl_156 ;
	7'h40 :
		rl_a54_t8 = RG_rl_156 ;
	7'h41 :
		rl_a54_t8 = RG_rl_156 ;
	7'h42 :
		rl_a54_t8 = RG_rl_156 ;
	7'h43 :
		rl_a54_t8 = RG_rl_156 ;
	7'h44 :
		rl_a54_t8 = RG_rl_156 ;
	7'h45 :
		rl_a54_t8 = RG_rl_156 ;
	7'h46 :
		rl_a54_t8 = RG_rl_156 ;
	7'h47 :
		rl_a54_t8 = RG_rl_156 ;
	7'h48 :
		rl_a54_t8 = RG_rl_156 ;
	7'h49 :
		rl_a54_t8 = RG_rl_156 ;
	7'h4a :
		rl_a54_t8 = RG_rl_156 ;
	7'h4b :
		rl_a54_t8 = RG_rl_156 ;
	7'h4c :
		rl_a54_t8 = RG_rl_156 ;
	7'h4d :
		rl_a54_t8 = RG_rl_156 ;
	7'h4e :
		rl_a54_t8 = RG_rl_156 ;
	7'h4f :
		rl_a54_t8 = RG_rl_156 ;
	7'h50 :
		rl_a54_t8 = RG_rl_156 ;
	7'h51 :
		rl_a54_t8 = RG_rl_156 ;
	7'h52 :
		rl_a54_t8 = RG_rl_156 ;
	7'h53 :
		rl_a54_t8 = RG_rl_156 ;
	7'h54 :
		rl_a54_t8 = RG_rl_156 ;
	7'h55 :
		rl_a54_t8 = RG_rl_156 ;
	7'h56 :
		rl_a54_t8 = RG_rl_156 ;
	7'h57 :
		rl_a54_t8 = RG_rl_156 ;
	7'h58 :
		rl_a54_t8 = RG_rl_156 ;
	7'h59 :
		rl_a54_t8 = RG_rl_156 ;
	7'h5a :
		rl_a54_t8 = RG_rl_156 ;
	7'h5b :
		rl_a54_t8 = RG_rl_156 ;
	7'h5c :
		rl_a54_t8 = RG_rl_156 ;
	7'h5d :
		rl_a54_t8 = RG_rl_156 ;
	7'h5e :
		rl_a54_t8 = RG_rl_156 ;
	7'h5f :
		rl_a54_t8 = RG_rl_156 ;
	7'h60 :
		rl_a54_t8 = RG_rl_156 ;
	7'h61 :
		rl_a54_t8 = RG_rl_156 ;
	7'h62 :
		rl_a54_t8 = RG_rl_156 ;
	7'h63 :
		rl_a54_t8 = RG_rl_156 ;
	7'h64 :
		rl_a54_t8 = RG_rl_156 ;
	7'h65 :
		rl_a54_t8 = RG_rl_156 ;
	7'h66 :
		rl_a54_t8 = RG_rl_156 ;
	7'h67 :
		rl_a54_t8 = RG_rl_156 ;
	7'h68 :
		rl_a54_t8 = RG_rl_156 ;
	7'h69 :
		rl_a54_t8 = RG_rl_156 ;
	7'h6a :
		rl_a54_t8 = RG_rl_156 ;
	7'h6b :
		rl_a54_t8 = RG_rl_156 ;
	7'h6c :
		rl_a54_t8 = RG_rl_156 ;
	7'h6d :
		rl_a54_t8 = RG_rl_156 ;
	7'h6e :
		rl_a54_t8 = RG_rl_156 ;
	7'h6f :
		rl_a54_t8 = RG_rl_156 ;
	7'h70 :
		rl_a54_t8 = RG_rl_156 ;
	7'h71 :
		rl_a54_t8 = RG_rl_156 ;
	7'h72 :
		rl_a54_t8 = RG_rl_156 ;
	7'h73 :
		rl_a54_t8 = RG_rl_156 ;
	7'h74 :
		rl_a54_t8 = RG_rl_156 ;
	7'h75 :
		rl_a54_t8 = RG_rl_156 ;
	7'h76 :
		rl_a54_t8 = RG_rl_156 ;
	7'h77 :
		rl_a54_t8 = RG_rl_156 ;
	7'h78 :
		rl_a54_t8 = RG_rl_156 ;
	7'h79 :
		rl_a54_t8 = RG_rl_156 ;
	7'h7a :
		rl_a54_t8 = RG_rl_156 ;
	7'h7b :
		rl_a54_t8 = RG_rl_156 ;
	7'h7c :
		rl_a54_t8 = RG_rl_156 ;
	7'h7d :
		rl_a54_t8 = RG_rl_156 ;
	7'h7e :
		rl_a54_t8 = RG_rl_156 ;
	7'h7f :
		rl_a54_t8 = RG_rl_156 ;
	default :
		rl_a54_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_25 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h01 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h02 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h03 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h04 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h05 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h06 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h07 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h08 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h09 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h0a :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h0b :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h0c :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h0d :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h0e :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h0f :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h10 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h11 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h12 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h13 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h14 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h15 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h16 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h17 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h18 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h19 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h1a :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h1b :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h1c :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h1d :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h1e :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h1f :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h20 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h21 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h22 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h23 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h24 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h25 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h26 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h27 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h28 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h29 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h2a :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h2b :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h2c :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h2d :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h2e :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h2f :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h30 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h31 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h32 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h33 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h34 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h35 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h36 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h37 :
		rl_a55_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h38 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h39 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h3a :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h3b :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h3c :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h3d :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h3e :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h3f :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h40 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h41 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h42 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h43 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h44 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h45 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h46 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h47 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h48 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h49 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h4a :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h4b :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h4c :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h4d :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h4e :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h4f :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h50 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h51 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h52 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h53 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h54 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h55 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h56 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h57 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h58 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h59 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h5a :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h5b :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h5c :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h5d :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h5e :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h5f :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h60 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h61 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h62 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h63 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h64 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h65 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h66 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h67 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h68 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h69 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h6a :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h6b :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h6c :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h6d :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h6e :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h6f :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h70 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h71 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h72 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h73 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h74 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h75 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h76 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h77 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h78 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h79 :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h7a :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h7b :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h7c :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h7d :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h7e :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	7'h7f :
		rl_a55_t8 = RG_quantized_block_rl_25 ;
	default :
		rl_a55_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_157 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a56_t8 = RG_rl_157 ;
	7'h01 :
		rl_a56_t8 = RG_rl_157 ;
	7'h02 :
		rl_a56_t8 = RG_rl_157 ;
	7'h03 :
		rl_a56_t8 = RG_rl_157 ;
	7'h04 :
		rl_a56_t8 = RG_rl_157 ;
	7'h05 :
		rl_a56_t8 = RG_rl_157 ;
	7'h06 :
		rl_a56_t8 = RG_rl_157 ;
	7'h07 :
		rl_a56_t8 = RG_rl_157 ;
	7'h08 :
		rl_a56_t8 = RG_rl_157 ;
	7'h09 :
		rl_a56_t8 = RG_rl_157 ;
	7'h0a :
		rl_a56_t8 = RG_rl_157 ;
	7'h0b :
		rl_a56_t8 = RG_rl_157 ;
	7'h0c :
		rl_a56_t8 = RG_rl_157 ;
	7'h0d :
		rl_a56_t8 = RG_rl_157 ;
	7'h0e :
		rl_a56_t8 = RG_rl_157 ;
	7'h0f :
		rl_a56_t8 = RG_rl_157 ;
	7'h10 :
		rl_a56_t8 = RG_rl_157 ;
	7'h11 :
		rl_a56_t8 = RG_rl_157 ;
	7'h12 :
		rl_a56_t8 = RG_rl_157 ;
	7'h13 :
		rl_a56_t8 = RG_rl_157 ;
	7'h14 :
		rl_a56_t8 = RG_rl_157 ;
	7'h15 :
		rl_a56_t8 = RG_rl_157 ;
	7'h16 :
		rl_a56_t8 = RG_rl_157 ;
	7'h17 :
		rl_a56_t8 = RG_rl_157 ;
	7'h18 :
		rl_a56_t8 = RG_rl_157 ;
	7'h19 :
		rl_a56_t8 = RG_rl_157 ;
	7'h1a :
		rl_a56_t8 = RG_rl_157 ;
	7'h1b :
		rl_a56_t8 = RG_rl_157 ;
	7'h1c :
		rl_a56_t8 = RG_rl_157 ;
	7'h1d :
		rl_a56_t8 = RG_rl_157 ;
	7'h1e :
		rl_a56_t8 = RG_rl_157 ;
	7'h1f :
		rl_a56_t8 = RG_rl_157 ;
	7'h20 :
		rl_a56_t8 = RG_rl_157 ;
	7'h21 :
		rl_a56_t8 = RG_rl_157 ;
	7'h22 :
		rl_a56_t8 = RG_rl_157 ;
	7'h23 :
		rl_a56_t8 = RG_rl_157 ;
	7'h24 :
		rl_a56_t8 = RG_rl_157 ;
	7'h25 :
		rl_a56_t8 = RG_rl_157 ;
	7'h26 :
		rl_a56_t8 = RG_rl_157 ;
	7'h27 :
		rl_a56_t8 = RG_rl_157 ;
	7'h28 :
		rl_a56_t8 = RG_rl_157 ;
	7'h29 :
		rl_a56_t8 = RG_rl_157 ;
	7'h2a :
		rl_a56_t8 = RG_rl_157 ;
	7'h2b :
		rl_a56_t8 = RG_rl_157 ;
	7'h2c :
		rl_a56_t8 = RG_rl_157 ;
	7'h2d :
		rl_a56_t8 = RG_rl_157 ;
	7'h2e :
		rl_a56_t8 = RG_rl_157 ;
	7'h2f :
		rl_a56_t8 = RG_rl_157 ;
	7'h30 :
		rl_a56_t8 = RG_rl_157 ;
	7'h31 :
		rl_a56_t8 = RG_rl_157 ;
	7'h32 :
		rl_a56_t8 = RG_rl_157 ;
	7'h33 :
		rl_a56_t8 = RG_rl_157 ;
	7'h34 :
		rl_a56_t8 = RG_rl_157 ;
	7'h35 :
		rl_a56_t8 = RG_rl_157 ;
	7'h36 :
		rl_a56_t8 = RG_rl_157 ;
	7'h37 :
		rl_a56_t8 = RG_rl_157 ;
	7'h38 :
		rl_a56_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h39 :
		rl_a56_t8 = RG_rl_157 ;
	7'h3a :
		rl_a56_t8 = RG_rl_157 ;
	7'h3b :
		rl_a56_t8 = RG_rl_157 ;
	7'h3c :
		rl_a56_t8 = RG_rl_157 ;
	7'h3d :
		rl_a56_t8 = RG_rl_157 ;
	7'h3e :
		rl_a56_t8 = RG_rl_157 ;
	7'h3f :
		rl_a56_t8 = RG_rl_157 ;
	7'h40 :
		rl_a56_t8 = RG_rl_157 ;
	7'h41 :
		rl_a56_t8 = RG_rl_157 ;
	7'h42 :
		rl_a56_t8 = RG_rl_157 ;
	7'h43 :
		rl_a56_t8 = RG_rl_157 ;
	7'h44 :
		rl_a56_t8 = RG_rl_157 ;
	7'h45 :
		rl_a56_t8 = RG_rl_157 ;
	7'h46 :
		rl_a56_t8 = RG_rl_157 ;
	7'h47 :
		rl_a56_t8 = RG_rl_157 ;
	7'h48 :
		rl_a56_t8 = RG_rl_157 ;
	7'h49 :
		rl_a56_t8 = RG_rl_157 ;
	7'h4a :
		rl_a56_t8 = RG_rl_157 ;
	7'h4b :
		rl_a56_t8 = RG_rl_157 ;
	7'h4c :
		rl_a56_t8 = RG_rl_157 ;
	7'h4d :
		rl_a56_t8 = RG_rl_157 ;
	7'h4e :
		rl_a56_t8 = RG_rl_157 ;
	7'h4f :
		rl_a56_t8 = RG_rl_157 ;
	7'h50 :
		rl_a56_t8 = RG_rl_157 ;
	7'h51 :
		rl_a56_t8 = RG_rl_157 ;
	7'h52 :
		rl_a56_t8 = RG_rl_157 ;
	7'h53 :
		rl_a56_t8 = RG_rl_157 ;
	7'h54 :
		rl_a56_t8 = RG_rl_157 ;
	7'h55 :
		rl_a56_t8 = RG_rl_157 ;
	7'h56 :
		rl_a56_t8 = RG_rl_157 ;
	7'h57 :
		rl_a56_t8 = RG_rl_157 ;
	7'h58 :
		rl_a56_t8 = RG_rl_157 ;
	7'h59 :
		rl_a56_t8 = RG_rl_157 ;
	7'h5a :
		rl_a56_t8 = RG_rl_157 ;
	7'h5b :
		rl_a56_t8 = RG_rl_157 ;
	7'h5c :
		rl_a56_t8 = RG_rl_157 ;
	7'h5d :
		rl_a56_t8 = RG_rl_157 ;
	7'h5e :
		rl_a56_t8 = RG_rl_157 ;
	7'h5f :
		rl_a56_t8 = RG_rl_157 ;
	7'h60 :
		rl_a56_t8 = RG_rl_157 ;
	7'h61 :
		rl_a56_t8 = RG_rl_157 ;
	7'h62 :
		rl_a56_t8 = RG_rl_157 ;
	7'h63 :
		rl_a56_t8 = RG_rl_157 ;
	7'h64 :
		rl_a56_t8 = RG_rl_157 ;
	7'h65 :
		rl_a56_t8 = RG_rl_157 ;
	7'h66 :
		rl_a56_t8 = RG_rl_157 ;
	7'h67 :
		rl_a56_t8 = RG_rl_157 ;
	7'h68 :
		rl_a56_t8 = RG_rl_157 ;
	7'h69 :
		rl_a56_t8 = RG_rl_157 ;
	7'h6a :
		rl_a56_t8 = RG_rl_157 ;
	7'h6b :
		rl_a56_t8 = RG_rl_157 ;
	7'h6c :
		rl_a56_t8 = RG_rl_157 ;
	7'h6d :
		rl_a56_t8 = RG_rl_157 ;
	7'h6e :
		rl_a56_t8 = RG_rl_157 ;
	7'h6f :
		rl_a56_t8 = RG_rl_157 ;
	7'h70 :
		rl_a56_t8 = RG_rl_157 ;
	7'h71 :
		rl_a56_t8 = RG_rl_157 ;
	7'h72 :
		rl_a56_t8 = RG_rl_157 ;
	7'h73 :
		rl_a56_t8 = RG_rl_157 ;
	7'h74 :
		rl_a56_t8 = RG_rl_157 ;
	7'h75 :
		rl_a56_t8 = RG_rl_157 ;
	7'h76 :
		rl_a56_t8 = RG_rl_157 ;
	7'h77 :
		rl_a56_t8 = RG_rl_157 ;
	7'h78 :
		rl_a56_t8 = RG_rl_157 ;
	7'h79 :
		rl_a56_t8 = RG_rl_157 ;
	7'h7a :
		rl_a56_t8 = RG_rl_157 ;
	7'h7b :
		rl_a56_t8 = RG_rl_157 ;
	7'h7c :
		rl_a56_t8 = RG_rl_157 ;
	7'h7d :
		rl_a56_t8 = RG_rl_157 ;
	7'h7e :
		rl_a56_t8 = RG_rl_157 ;
	7'h7f :
		rl_a56_t8 = RG_rl_157 ;
	default :
		rl_a56_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_26 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h01 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h02 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h03 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h04 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h05 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h06 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h07 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h08 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h09 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h0a :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h0b :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h0c :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h0d :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h0e :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h0f :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h10 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h11 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h12 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h13 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h14 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h15 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h16 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h17 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h18 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h19 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h1a :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h1b :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h1c :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h1d :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h1e :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h1f :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h20 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h21 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h22 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h23 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h24 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h25 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h26 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h27 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h28 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h29 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h2a :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h2b :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h2c :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h2d :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h2e :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h2f :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h30 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h31 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h32 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h33 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h34 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h35 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h36 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h37 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h38 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h39 :
		rl_a57_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h3a :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h3b :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h3c :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h3d :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h3e :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h3f :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h40 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h41 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h42 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h43 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h44 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h45 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h46 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h47 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h48 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h49 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h4a :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h4b :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h4c :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h4d :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h4e :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h4f :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h50 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h51 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h52 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h53 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h54 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h55 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h56 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h57 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h58 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h59 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h5a :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h5b :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h5c :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h5d :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h5e :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h5f :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h60 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h61 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h62 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h63 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h64 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h65 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h66 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h67 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h68 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h69 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h6a :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h6b :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h6c :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h6d :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h6e :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h6f :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h70 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h71 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h72 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h73 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h74 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h75 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h76 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h77 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h78 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h79 :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h7a :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h7b :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h7c :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h7d :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h7e :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	7'h7f :
		rl_a57_t8 = RG_quantized_block_rl_26 ;
	default :
		rl_a57_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_158 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a58_t8 = RG_rl_158 ;
	7'h01 :
		rl_a58_t8 = RG_rl_158 ;
	7'h02 :
		rl_a58_t8 = RG_rl_158 ;
	7'h03 :
		rl_a58_t8 = RG_rl_158 ;
	7'h04 :
		rl_a58_t8 = RG_rl_158 ;
	7'h05 :
		rl_a58_t8 = RG_rl_158 ;
	7'h06 :
		rl_a58_t8 = RG_rl_158 ;
	7'h07 :
		rl_a58_t8 = RG_rl_158 ;
	7'h08 :
		rl_a58_t8 = RG_rl_158 ;
	7'h09 :
		rl_a58_t8 = RG_rl_158 ;
	7'h0a :
		rl_a58_t8 = RG_rl_158 ;
	7'h0b :
		rl_a58_t8 = RG_rl_158 ;
	7'h0c :
		rl_a58_t8 = RG_rl_158 ;
	7'h0d :
		rl_a58_t8 = RG_rl_158 ;
	7'h0e :
		rl_a58_t8 = RG_rl_158 ;
	7'h0f :
		rl_a58_t8 = RG_rl_158 ;
	7'h10 :
		rl_a58_t8 = RG_rl_158 ;
	7'h11 :
		rl_a58_t8 = RG_rl_158 ;
	7'h12 :
		rl_a58_t8 = RG_rl_158 ;
	7'h13 :
		rl_a58_t8 = RG_rl_158 ;
	7'h14 :
		rl_a58_t8 = RG_rl_158 ;
	7'h15 :
		rl_a58_t8 = RG_rl_158 ;
	7'h16 :
		rl_a58_t8 = RG_rl_158 ;
	7'h17 :
		rl_a58_t8 = RG_rl_158 ;
	7'h18 :
		rl_a58_t8 = RG_rl_158 ;
	7'h19 :
		rl_a58_t8 = RG_rl_158 ;
	7'h1a :
		rl_a58_t8 = RG_rl_158 ;
	7'h1b :
		rl_a58_t8 = RG_rl_158 ;
	7'h1c :
		rl_a58_t8 = RG_rl_158 ;
	7'h1d :
		rl_a58_t8 = RG_rl_158 ;
	7'h1e :
		rl_a58_t8 = RG_rl_158 ;
	7'h1f :
		rl_a58_t8 = RG_rl_158 ;
	7'h20 :
		rl_a58_t8 = RG_rl_158 ;
	7'h21 :
		rl_a58_t8 = RG_rl_158 ;
	7'h22 :
		rl_a58_t8 = RG_rl_158 ;
	7'h23 :
		rl_a58_t8 = RG_rl_158 ;
	7'h24 :
		rl_a58_t8 = RG_rl_158 ;
	7'h25 :
		rl_a58_t8 = RG_rl_158 ;
	7'h26 :
		rl_a58_t8 = RG_rl_158 ;
	7'h27 :
		rl_a58_t8 = RG_rl_158 ;
	7'h28 :
		rl_a58_t8 = RG_rl_158 ;
	7'h29 :
		rl_a58_t8 = RG_rl_158 ;
	7'h2a :
		rl_a58_t8 = RG_rl_158 ;
	7'h2b :
		rl_a58_t8 = RG_rl_158 ;
	7'h2c :
		rl_a58_t8 = RG_rl_158 ;
	7'h2d :
		rl_a58_t8 = RG_rl_158 ;
	7'h2e :
		rl_a58_t8 = RG_rl_158 ;
	7'h2f :
		rl_a58_t8 = RG_rl_158 ;
	7'h30 :
		rl_a58_t8 = RG_rl_158 ;
	7'h31 :
		rl_a58_t8 = RG_rl_158 ;
	7'h32 :
		rl_a58_t8 = RG_rl_158 ;
	7'h33 :
		rl_a58_t8 = RG_rl_158 ;
	7'h34 :
		rl_a58_t8 = RG_rl_158 ;
	7'h35 :
		rl_a58_t8 = RG_rl_158 ;
	7'h36 :
		rl_a58_t8 = RG_rl_158 ;
	7'h37 :
		rl_a58_t8 = RG_rl_158 ;
	7'h38 :
		rl_a58_t8 = RG_rl_158 ;
	7'h39 :
		rl_a58_t8 = RG_rl_158 ;
	7'h3a :
		rl_a58_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h3b :
		rl_a58_t8 = RG_rl_158 ;
	7'h3c :
		rl_a58_t8 = RG_rl_158 ;
	7'h3d :
		rl_a58_t8 = RG_rl_158 ;
	7'h3e :
		rl_a58_t8 = RG_rl_158 ;
	7'h3f :
		rl_a58_t8 = RG_rl_158 ;
	7'h40 :
		rl_a58_t8 = RG_rl_158 ;
	7'h41 :
		rl_a58_t8 = RG_rl_158 ;
	7'h42 :
		rl_a58_t8 = RG_rl_158 ;
	7'h43 :
		rl_a58_t8 = RG_rl_158 ;
	7'h44 :
		rl_a58_t8 = RG_rl_158 ;
	7'h45 :
		rl_a58_t8 = RG_rl_158 ;
	7'h46 :
		rl_a58_t8 = RG_rl_158 ;
	7'h47 :
		rl_a58_t8 = RG_rl_158 ;
	7'h48 :
		rl_a58_t8 = RG_rl_158 ;
	7'h49 :
		rl_a58_t8 = RG_rl_158 ;
	7'h4a :
		rl_a58_t8 = RG_rl_158 ;
	7'h4b :
		rl_a58_t8 = RG_rl_158 ;
	7'h4c :
		rl_a58_t8 = RG_rl_158 ;
	7'h4d :
		rl_a58_t8 = RG_rl_158 ;
	7'h4e :
		rl_a58_t8 = RG_rl_158 ;
	7'h4f :
		rl_a58_t8 = RG_rl_158 ;
	7'h50 :
		rl_a58_t8 = RG_rl_158 ;
	7'h51 :
		rl_a58_t8 = RG_rl_158 ;
	7'h52 :
		rl_a58_t8 = RG_rl_158 ;
	7'h53 :
		rl_a58_t8 = RG_rl_158 ;
	7'h54 :
		rl_a58_t8 = RG_rl_158 ;
	7'h55 :
		rl_a58_t8 = RG_rl_158 ;
	7'h56 :
		rl_a58_t8 = RG_rl_158 ;
	7'h57 :
		rl_a58_t8 = RG_rl_158 ;
	7'h58 :
		rl_a58_t8 = RG_rl_158 ;
	7'h59 :
		rl_a58_t8 = RG_rl_158 ;
	7'h5a :
		rl_a58_t8 = RG_rl_158 ;
	7'h5b :
		rl_a58_t8 = RG_rl_158 ;
	7'h5c :
		rl_a58_t8 = RG_rl_158 ;
	7'h5d :
		rl_a58_t8 = RG_rl_158 ;
	7'h5e :
		rl_a58_t8 = RG_rl_158 ;
	7'h5f :
		rl_a58_t8 = RG_rl_158 ;
	7'h60 :
		rl_a58_t8 = RG_rl_158 ;
	7'h61 :
		rl_a58_t8 = RG_rl_158 ;
	7'h62 :
		rl_a58_t8 = RG_rl_158 ;
	7'h63 :
		rl_a58_t8 = RG_rl_158 ;
	7'h64 :
		rl_a58_t8 = RG_rl_158 ;
	7'h65 :
		rl_a58_t8 = RG_rl_158 ;
	7'h66 :
		rl_a58_t8 = RG_rl_158 ;
	7'h67 :
		rl_a58_t8 = RG_rl_158 ;
	7'h68 :
		rl_a58_t8 = RG_rl_158 ;
	7'h69 :
		rl_a58_t8 = RG_rl_158 ;
	7'h6a :
		rl_a58_t8 = RG_rl_158 ;
	7'h6b :
		rl_a58_t8 = RG_rl_158 ;
	7'h6c :
		rl_a58_t8 = RG_rl_158 ;
	7'h6d :
		rl_a58_t8 = RG_rl_158 ;
	7'h6e :
		rl_a58_t8 = RG_rl_158 ;
	7'h6f :
		rl_a58_t8 = RG_rl_158 ;
	7'h70 :
		rl_a58_t8 = RG_rl_158 ;
	7'h71 :
		rl_a58_t8 = RG_rl_158 ;
	7'h72 :
		rl_a58_t8 = RG_rl_158 ;
	7'h73 :
		rl_a58_t8 = RG_rl_158 ;
	7'h74 :
		rl_a58_t8 = RG_rl_158 ;
	7'h75 :
		rl_a58_t8 = RG_rl_158 ;
	7'h76 :
		rl_a58_t8 = RG_rl_158 ;
	7'h77 :
		rl_a58_t8 = RG_rl_158 ;
	7'h78 :
		rl_a58_t8 = RG_rl_158 ;
	7'h79 :
		rl_a58_t8 = RG_rl_158 ;
	7'h7a :
		rl_a58_t8 = RG_rl_158 ;
	7'h7b :
		rl_a58_t8 = RG_rl_158 ;
	7'h7c :
		rl_a58_t8 = RG_rl_158 ;
	7'h7d :
		rl_a58_t8 = RG_rl_158 ;
	7'h7e :
		rl_a58_t8 = RG_rl_158 ;
	7'h7f :
		rl_a58_t8 = RG_rl_158 ;
	default :
		rl_a58_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_27 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h01 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h02 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h03 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h04 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h05 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h06 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h07 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h08 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h09 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h0a :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h0b :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h0c :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h0d :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h0e :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h0f :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h10 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h11 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h12 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h13 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h14 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h15 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h16 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h17 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h18 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h19 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h1a :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h1b :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h1c :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h1d :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h1e :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h1f :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h20 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h21 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h22 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h23 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h24 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h25 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h26 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h27 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h28 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h29 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h2a :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h2b :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h2c :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h2d :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h2e :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h2f :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h30 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h31 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h32 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h33 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h34 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h35 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h36 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h37 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h38 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h39 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h3a :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h3b :
		rl_a59_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h3c :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h3d :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h3e :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h3f :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h40 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h41 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h42 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h43 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h44 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h45 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h46 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h47 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h48 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h49 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h4a :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h4b :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h4c :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h4d :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h4e :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h4f :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h50 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h51 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h52 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h53 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h54 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h55 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h56 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h57 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h58 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h59 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h5a :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h5b :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h5c :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h5d :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h5e :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h5f :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h60 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h61 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h62 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h63 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h64 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h65 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h66 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h67 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h68 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h69 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h6a :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h6b :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h6c :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h6d :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h6e :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h6f :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h70 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h71 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h72 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h73 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h74 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h75 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h76 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h77 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h78 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h79 :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h7a :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h7b :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h7c :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h7d :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h7e :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	7'h7f :
		rl_a59_t8 = RG_quantized_block_rl_27 ;
	default :
		rl_a59_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_159 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a60_t8 = RG_rl_159 ;
	7'h01 :
		rl_a60_t8 = RG_rl_159 ;
	7'h02 :
		rl_a60_t8 = RG_rl_159 ;
	7'h03 :
		rl_a60_t8 = RG_rl_159 ;
	7'h04 :
		rl_a60_t8 = RG_rl_159 ;
	7'h05 :
		rl_a60_t8 = RG_rl_159 ;
	7'h06 :
		rl_a60_t8 = RG_rl_159 ;
	7'h07 :
		rl_a60_t8 = RG_rl_159 ;
	7'h08 :
		rl_a60_t8 = RG_rl_159 ;
	7'h09 :
		rl_a60_t8 = RG_rl_159 ;
	7'h0a :
		rl_a60_t8 = RG_rl_159 ;
	7'h0b :
		rl_a60_t8 = RG_rl_159 ;
	7'h0c :
		rl_a60_t8 = RG_rl_159 ;
	7'h0d :
		rl_a60_t8 = RG_rl_159 ;
	7'h0e :
		rl_a60_t8 = RG_rl_159 ;
	7'h0f :
		rl_a60_t8 = RG_rl_159 ;
	7'h10 :
		rl_a60_t8 = RG_rl_159 ;
	7'h11 :
		rl_a60_t8 = RG_rl_159 ;
	7'h12 :
		rl_a60_t8 = RG_rl_159 ;
	7'h13 :
		rl_a60_t8 = RG_rl_159 ;
	7'h14 :
		rl_a60_t8 = RG_rl_159 ;
	7'h15 :
		rl_a60_t8 = RG_rl_159 ;
	7'h16 :
		rl_a60_t8 = RG_rl_159 ;
	7'h17 :
		rl_a60_t8 = RG_rl_159 ;
	7'h18 :
		rl_a60_t8 = RG_rl_159 ;
	7'h19 :
		rl_a60_t8 = RG_rl_159 ;
	7'h1a :
		rl_a60_t8 = RG_rl_159 ;
	7'h1b :
		rl_a60_t8 = RG_rl_159 ;
	7'h1c :
		rl_a60_t8 = RG_rl_159 ;
	7'h1d :
		rl_a60_t8 = RG_rl_159 ;
	7'h1e :
		rl_a60_t8 = RG_rl_159 ;
	7'h1f :
		rl_a60_t8 = RG_rl_159 ;
	7'h20 :
		rl_a60_t8 = RG_rl_159 ;
	7'h21 :
		rl_a60_t8 = RG_rl_159 ;
	7'h22 :
		rl_a60_t8 = RG_rl_159 ;
	7'h23 :
		rl_a60_t8 = RG_rl_159 ;
	7'h24 :
		rl_a60_t8 = RG_rl_159 ;
	7'h25 :
		rl_a60_t8 = RG_rl_159 ;
	7'h26 :
		rl_a60_t8 = RG_rl_159 ;
	7'h27 :
		rl_a60_t8 = RG_rl_159 ;
	7'h28 :
		rl_a60_t8 = RG_rl_159 ;
	7'h29 :
		rl_a60_t8 = RG_rl_159 ;
	7'h2a :
		rl_a60_t8 = RG_rl_159 ;
	7'h2b :
		rl_a60_t8 = RG_rl_159 ;
	7'h2c :
		rl_a60_t8 = RG_rl_159 ;
	7'h2d :
		rl_a60_t8 = RG_rl_159 ;
	7'h2e :
		rl_a60_t8 = RG_rl_159 ;
	7'h2f :
		rl_a60_t8 = RG_rl_159 ;
	7'h30 :
		rl_a60_t8 = RG_rl_159 ;
	7'h31 :
		rl_a60_t8 = RG_rl_159 ;
	7'h32 :
		rl_a60_t8 = RG_rl_159 ;
	7'h33 :
		rl_a60_t8 = RG_rl_159 ;
	7'h34 :
		rl_a60_t8 = RG_rl_159 ;
	7'h35 :
		rl_a60_t8 = RG_rl_159 ;
	7'h36 :
		rl_a60_t8 = RG_rl_159 ;
	7'h37 :
		rl_a60_t8 = RG_rl_159 ;
	7'h38 :
		rl_a60_t8 = RG_rl_159 ;
	7'h39 :
		rl_a60_t8 = RG_rl_159 ;
	7'h3a :
		rl_a60_t8 = RG_rl_159 ;
	7'h3b :
		rl_a60_t8 = RG_rl_159 ;
	7'h3c :
		rl_a60_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h3d :
		rl_a60_t8 = RG_rl_159 ;
	7'h3e :
		rl_a60_t8 = RG_rl_159 ;
	7'h3f :
		rl_a60_t8 = RG_rl_159 ;
	7'h40 :
		rl_a60_t8 = RG_rl_159 ;
	7'h41 :
		rl_a60_t8 = RG_rl_159 ;
	7'h42 :
		rl_a60_t8 = RG_rl_159 ;
	7'h43 :
		rl_a60_t8 = RG_rl_159 ;
	7'h44 :
		rl_a60_t8 = RG_rl_159 ;
	7'h45 :
		rl_a60_t8 = RG_rl_159 ;
	7'h46 :
		rl_a60_t8 = RG_rl_159 ;
	7'h47 :
		rl_a60_t8 = RG_rl_159 ;
	7'h48 :
		rl_a60_t8 = RG_rl_159 ;
	7'h49 :
		rl_a60_t8 = RG_rl_159 ;
	7'h4a :
		rl_a60_t8 = RG_rl_159 ;
	7'h4b :
		rl_a60_t8 = RG_rl_159 ;
	7'h4c :
		rl_a60_t8 = RG_rl_159 ;
	7'h4d :
		rl_a60_t8 = RG_rl_159 ;
	7'h4e :
		rl_a60_t8 = RG_rl_159 ;
	7'h4f :
		rl_a60_t8 = RG_rl_159 ;
	7'h50 :
		rl_a60_t8 = RG_rl_159 ;
	7'h51 :
		rl_a60_t8 = RG_rl_159 ;
	7'h52 :
		rl_a60_t8 = RG_rl_159 ;
	7'h53 :
		rl_a60_t8 = RG_rl_159 ;
	7'h54 :
		rl_a60_t8 = RG_rl_159 ;
	7'h55 :
		rl_a60_t8 = RG_rl_159 ;
	7'h56 :
		rl_a60_t8 = RG_rl_159 ;
	7'h57 :
		rl_a60_t8 = RG_rl_159 ;
	7'h58 :
		rl_a60_t8 = RG_rl_159 ;
	7'h59 :
		rl_a60_t8 = RG_rl_159 ;
	7'h5a :
		rl_a60_t8 = RG_rl_159 ;
	7'h5b :
		rl_a60_t8 = RG_rl_159 ;
	7'h5c :
		rl_a60_t8 = RG_rl_159 ;
	7'h5d :
		rl_a60_t8 = RG_rl_159 ;
	7'h5e :
		rl_a60_t8 = RG_rl_159 ;
	7'h5f :
		rl_a60_t8 = RG_rl_159 ;
	7'h60 :
		rl_a60_t8 = RG_rl_159 ;
	7'h61 :
		rl_a60_t8 = RG_rl_159 ;
	7'h62 :
		rl_a60_t8 = RG_rl_159 ;
	7'h63 :
		rl_a60_t8 = RG_rl_159 ;
	7'h64 :
		rl_a60_t8 = RG_rl_159 ;
	7'h65 :
		rl_a60_t8 = RG_rl_159 ;
	7'h66 :
		rl_a60_t8 = RG_rl_159 ;
	7'h67 :
		rl_a60_t8 = RG_rl_159 ;
	7'h68 :
		rl_a60_t8 = RG_rl_159 ;
	7'h69 :
		rl_a60_t8 = RG_rl_159 ;
	7'h6a :
		rl_a60_t8 = RG_rl_159 ;
	7'h6b :
		rl_a60_t8 = RG_rl_159 ;
	7'h6c :
		rl_a60_t8 = RG_rl_159 ;
	7'h6d :
		rl_a60_t8 = RG_rl_159 ;
	7'h6e :
		rl_a60_t8 = RG_rl_159 ;
	7'h6f :
		rl_a60_t8 = RG_rl_159 ;
	7'h70 :
		rl_a60_t8 = RG_rl_159 ;
	7'h71 :
		rl_a60_t8 = RG_rl_159 ;
	7'h72 :
		rl_a60_t8 = RG_rl_159 ;
	7'h73 :
		rl_a60_t8 = RG_rl_159 ;
	7'h74 :
		rl_a60_t8 = RG_rl_159 ;
	7'h75 :
		rl_a60_t8 = RG_rl_159 ;
	7'h76 :
		rl_a60_t8 = RG_rl_159 ;
	7'h77 :
		rl_a60_t8 = RG_rl_159 ;
	7'h78 :
		rl_a60_t8 = RG_rl_159 ;
	7'h79 :
		rl_a60_t8 = RG_rl_159 ;
	7'h7a :
		rl_a60_t8 = RG_rl_159 ;
	7'h7b :
		rl_a60_t8 = RG_rl_159 ;
	7'h7c :
		rl_a60_t8 = RG_rl_159 ;
	7'h7d :
		rl_a60_t8 = RG_rl_159 ;
	7'h7e :
		rl_a60_t8 = RG_rl_159 ;
	7'h7f :
		rl_a60_t8 = RG_rl_159 ;
	default :
		rl_a60_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_28 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h01 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h02 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h03 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h04 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h05 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h06 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h07 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h08 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h09 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h0a :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h0b :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h0c :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h0d :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h0e :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h0f :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h10 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h11 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h12 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h13 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h14 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h15 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h16 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h17 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h18 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h19 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h1a :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h1b :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h1c :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h1d :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h1e :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h1f :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h20 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h21 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h22 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h23 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h24 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h25 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h26 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h27 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h28 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h29 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h2a :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h2b :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h2c :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h2d :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h2e :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h2f :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h30 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h31 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h32 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h33 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h34 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h35 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h36 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h37 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h38 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h39 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h3a :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h3b :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h3c :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h3d :
		rl_a61_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h3e :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h3f :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h40 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h41 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h42 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h43 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h44 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h45 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h46 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h47 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h48 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h49 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h4a :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h4b :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h4c :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h4d :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h4e :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h4f :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h50 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h51 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h52 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h53 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h54 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h55 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h56 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h57 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h58 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h59 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h5a :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h5b :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h5c :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h5d :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h5e :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h5f :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h60 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h61 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h62 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h63 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h64 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h65 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h66 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h67 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h68 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h69 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h6a :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h6b :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h6c :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h6d :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h6e :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h6f :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h70 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h71 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h72 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h73 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h74 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h75 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h76 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h77 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h78 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h79 :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h7a :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h7b :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h7c :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h7d :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h7e :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	7'h7f :
		rl_a61_t8 = RG_quantized_block_rl_28 ;
	default :
		rl_a61_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_160 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a62_t8 = RG_rl_160 ;
	7'h01 :
		rl_a62_t8 = RG_rl_160 ;
	7'h02 :
		rl_a62_t8 = RG_rl_160 ;
	7'h03 :
		rl_a62_t8 = RG_rl_160 ;
	7'h04 :
		rl_a62_t8 = RG_rl_160 ;
	7'h05 :
		rl_a62_t8 = RG_rl_160 ;
	7'h06 :
		rl_a62_t8 = RG_rl_160 ;
	7'h07 :
		rl_a62_t8 = RG_rl_160 ;
	7'h08 :
		rl_a62_t8 = RG_rl_160 ;
	7'h09 :
		rl_a62_t8 = RG_rl_160 ;
	7'h0a :
		rl_a62_t8 = RG_rl_160 ;
	7'h0b :
		rl_a62_t8 = RG_rl_160 ;
	7'h0c :
		rl_a62_t8 = RG_rl_160 ;
	7'h0d :
		rl_a62_t8 = RG_rl_160 ;
	7'h0e :
		rl_a62_t8 = RG_rl_160 ;
	7'h0f :
		rl_a62_t8 = RG_rl_160 ;
	7'h10 :
		rl_a62_t8 = RG_rl_160 ;
	7'h11 :
		rl_a62_t8 = RG_rl_160 ;
	7'h12 :
		rl_a62_t8 = RG_rl_160 ;
	7'h13 :
		rl_a62_t8 = RG_rl_160 ;
	7'h14 :
		rl_a62_t8 = RG_rl_160 ;
	7'h15 :
		rl_a62_t8 = RG_rl_160 ;
	7'h16 :
		rl_a62_t8 = RG_rl_160 ;
	7'h17 :
		rl_a62_t8 = RG_rl_160 ;
	7'h18 :
		rl_a62_t8 = RG_rl_160 ;
	7'h19 :
		rl_a62_t8 = RG_rl_160 ;
	7'h1a :
		rl_a62_t8 = RG_rl_160 ;
	7'h1b :
		rl_a62_t8 = RG_rl_160 ;
	7'h1c :
		rl_a62_t8 = RG_rl_160 ;
	7'h1d :
		rl_a62_t8 = RG_rl_160 ;
	7'h1e :
		rl_a62_t8 = RG_rl_160 ;
	7'h1f :
		rl_a62_t8 = RG_rl_160 ;
	7'h20 :
		rl_a62_t8 = RG_rl_160 ;
	7'h21 :
		rl_a62_t8 = RG_rl_160 ;
	7'h22 :
		rl_a62_t8 = RG_rl_160 ;
	7'h23 :
		rl_a62_t8 = RG_rl_160 ;
	7'h24 :
		rl_a62_t8 = RG_rl_160 ;
	7'h25 :
		rl_a62_t8 = RG_rl_160 ;
	7'h26 :
		rl_a62_t8 = RG_rl_160 ;
	7'h27 :
		rl_a62_t8 = RG_rl_160 ;
	7'h28 :
		rl_a62_t8 = RG_rl_160 ;
	7'h29 :
		rl_a62_t8 = RG_rl_160 ;
	7'h2a :
		rl_a62_t8 = RG_rl_160 ;
	7'h2b :
		rl_a62_t8 = RG_rl_160 ;
	7'h2c :
		rl_a62_t8 = RG_rl_160 ;
	7'h2d :
		rl_a62_t8 = RG_rl_160 ;
	7'h2e :
		rl_a62_t8 = RG_rl_160 ;
	7'h2f :
		rl_a62_t8 = RG_rl_160 ;
	7'h30 :
		rl_a62_t8 = RG_rl_160 ;
	7'h31 :
		rl_a62_t8 = RG_rl_160 ;
	7'h32 :
		rl_a62_t8 = RG_rl_160 ;
	7'h33 :
		rl_a62_t8 = RG_rl_160 ;
	7'h34 :
		rl_a62_t8 = RG_rl_160 ;
	7'h35 :
		rl_a62_t8 = RG_rl_160 ;
	7'h36 :
		rl_a62_t8 = RG_rl_160 ;
	7'h37 :
		rl_a62_t8 = RG_rl_160 ;
	7'h38 :
		rl_a62_t8 = RG_rl_160 ;
	7'h39 :
		rl_a62_t8 = RG_rl_160 ;
	7'h3a :
		rl_a62_t8 = RG_rl_160 ;
	7'h3b :
		rl_a62_t8 = RG_rl_160 ;
	7'h3c :
		rl_a62_t8 = RG_rl_160 ;
	7'h3d :
		rl_a62_t8 = RG_rl_160 ;
	7'h3e :
		rl_a62_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h3f :
		rl_a62_t8 = RG_rl_160 ;
	7'h40 :
		rl_a62_t8 = RG_rl_160 ;
	7'h41 :
		rl_a62_t8 = RG_rl_160 ;
	7'h42 :
		rl_a62_t8 = RG_rl_160 ;
	7'h43 :
		rl_a62_t8 = RG_rl_160 ;
	7'h44 :
		rl_a62_t8 = RG_rl_160 ;
	7'h45 :
		rl_a62_t8 = RG_rl_160 ;
	7'h46 :
		rl_a62_t8 = RG_rl_160 ;
	7'h47 :
		rl_a62_t8 = RG_rl_160 ;
	7'h48 :
		rl_a62_t8 = RG_rl_160 ;
	7'h49 :
		rl_a62_t8 = RG_rl_160 ;
	7'h4a :
		rl_a62_t8 = RG_rl_160 ;
	7'h4b :
		rl_a62_t8 = RG_rl_160 ;
	7'h4c :
		rl_a62_t8 = RG_rl_160 ;
	7'h4d :
		rl_a62_t8 = RG_rl_160 ;
	7'h4e :
		rl_a62_t8 = RG_rl_160 ;
	7'h4f :
		rl_a62_t8 = RG_rl_160 ;
	7'h50 :
		rl_a62_t8 = RG_rl_160 ;
	7'h51 :
		rl_a62_t8 = RG_rl_160 ;
	7'h52 :
		rl_a62_t8 = RG_rl_160 ;
	7'h53 :
		rl_a62_t8 = RG_rl_160 ;
	7'h54 :
		rl_a62_t8 = RG_rl_160 ;
	7'h55 :
		rl_a62_t8 = RG_rl_160 ;
	7'h56 :
		rl_a62_t8 = RG_rl_160 ;
	7'h57 :
		rl_a62_t8 = RG_rl_160 ;
	7'h58 :
		rl_a62_t8 = RG_rl_160 ;
	7'h59 :
		rl_a62_t8 = RG_rl_160 ;
	7'h5a :
		rl_a62_t8 = RG_rl_160 ;
	7'h5b :
		rl_a62_t8 = RG_rl_160 ;
	7'h5c :
		rl_a62_t8 = RG_rl_160 ;
	7'h5d :
		rl_a62_t8 = RG_rl_160 ;
	7'h5e :
		rl_a62_t8 = RG_rl_160 ;
	7'h5f :
		rl_a62_t8 = RG_rl_160 ;
	7'h60 :
		rl_a62_t8 = RG_rl_160 ;
	7'h61 :
		rl_a62_t8 = RG_rl_160 ;
	7'h62 :
		rl_a62_t8 = RG_rl_160 ;
	7'h63 :
		rl_a62_t8 = RG_rl_160 ;
	7'h64 :
		rl_a62_t8 = RG_rl_160 ;
	7'h65 :
		rl_a62_t8 = RG_rl_160 ;
	7'h66 :
		rl_a62_t8 = RG_rl_160 ;
	7'h67 :
		rl_a62_t8 = RG_rl_160 ;
	7'h68 :
		rl_a62_t8 = RG_rl_160 ;
	7'h69 :
		rl_a62_t8 = RG_rl_160 ;
	7'h6a :
		rl_a62_t8 = RG_rl_160 ;
	7'h6b :
		rl_a62_t8 = RG_rl_160 ;
	7'h6c :
		rl_a62_t8 = RG_rl_160 ;
	7'h6d :
		rl_a62_t8 = RG_rl_160 ;
	7'h6e :
		rl_a62_t8 = RG_rl_160 ;
	7'h6f :
		rl_a62_t8 = RG_rl_160 ;
	7'h70 :
		rl_a62_t8 = RG_rl_160 ;
	7'h71 :
		rl_a62_t8 = RG_rl_160 ;
	7'h72 :
		rl_a62_t8 = RG_rl_160 ;
	7'h73 :
		rl_a62_t8 = RG_rl_160 ;
	7'h74 :
		rl_a62_t8 = RG_rl_160 ;
	7'h75 :
		rl_a62_t8 = RG_rl_160 ;
	7'h76 :
		rl_a62_t8 = RG_rl_160 ;
	7'h77 :
		rl_a62_t8 = RG_rl_160 ;
	7'h78 :
		rl_a62_t8 = RG_rl_160 ;
	7'h79 :
		rl_a62_t8 = RG_rl_160 ;
	7'h7a :
		rl_a62_t8 = RG_rl_160 ;
	7'h7b :
		rl_a62_t8 = RG_rl_160 ;
	7'h7c :
		rl_a62_t8 = RG_rl_160 ;
	7'h7d :
		rl_a62_t8 = RG_rl_160 ;
	7'h7e :
		rl_a62_t8 = RG_rl_160 ;
	7'h7f :
		rl_a62_t8 = RG_rl_160 ;
	default :
		rl_a62_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_29 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h01 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h02 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h03 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h04 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h05 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h06 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h07 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h08 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h09 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h0a :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h0b :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h0c :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h0d :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h0e :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h0f :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h10 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h11 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h12 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h13 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h14 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h15 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h16 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h17 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h18 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h19 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h1a :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h1b :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h1c :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h1d :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h1e :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h1f :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h20 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h21 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h22 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h23 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h24 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h25 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h26 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h27 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h28 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h29 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h2a :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h2b :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h2c :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h2d :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h2e :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h2f :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h30 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h31 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h32 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h33 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h34 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h35 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h36 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h37 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h38 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h39 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h3a :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h3b :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h3c :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h3d :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h3e :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h3f :
		rl_a63_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h40 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h41 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h42 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h43 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h44 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h45 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h46 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h47 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h48 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h49 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h4a :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h4b :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h4c :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h4d :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h4e :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h4f :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h50 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h51 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h52 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h53 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h54 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h55 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h56 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h57 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h58 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h59 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h5a :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h5b :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h5c :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h5d :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h5e :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h5f :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h60 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h61 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h62 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h63 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h64 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h65 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h66 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h67 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h68 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h69 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h6a :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h6b :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h6c :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h6d :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h6e :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h6f :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h70 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h71 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h72 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h73 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h74 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h75 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h76 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h77 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h78 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h79 :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h7a :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h7b :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h7c :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h7d :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h7e :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	7'h7f :
		rl_a63_t8 = RG_quantized_block_rl_29 ;
	default :
		rl_a63_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_161 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a64_t8 = RG_rl_161 ;
	7'h01 :
		rl_a64_t8 = RG_rl_161 ;
	7'h02 :
		rl_a64_t8 = RG_rl_161 ;
	7'h03 :
		rl_a64_t8 = RG_rl_161 ;
	7'h04 :
		rl_a64_t8 = RG_rl_161 ;
	7'h05 :
		rl_a64_t8 = RG_rl_161 ;
	7'h06 :
		rl_a64_t8 = RG_rl_161 ;
	7'h07 :
		rl_a64_t8 = RG_rl_161 ;
	7'h08 :
		rl_a64_t8 = RG_rl_161 ;
	7'h09 :
		rl_a64_t8 = RG_rl_161 ;
	7'h0a :
		rl_a64_t8 = RG_rl_161 ;
	7'h0b :
		rl_a64_t8 = RG_rl_161 ;
	7'h0c :
		rl_a64_t8 = RG_rl_161 ;
	7'h0d :
		rl_a64_t8 = RG_rl_161 ;
	7'h0e :
		rl_a64_t8 = RG_rl_161 ;
	7'h0f :
		rl_a64_t8 = RG_rl_161 ;
	7'h10 :
		rl_a64_t8 = RG_rl_161 ;
	7'h11 :
		rl_a64_t8 = RG_rl_161 ;
	7'h12 :
		rl_a64_t8 = RG_rl_161 ;
	7'h13 :
		rl_a64_t8 = RG_rl_161 ;
	7'h14 :
		rl_a64_t8 = RG_rl_161 ;
	7'h15 :
		rl_a64_t8 = RG_rl_161 ;
	7'h16 :
		rl_a64_t8 = RG_rl_161 ;
	7'h17 :
		rl_a64_t8 = RG_rl_161 ;
	7'h18 :
		rl_a64_t8 = RG_rl_161 ;
	7'h19 :
		rl_a64_t8 = RG_rl_161 ;
	7'h1a :
		rl_a64_t8 = RG_rl_161 ;
	7'h1b :
		rl_a64_t8 = RG_rl_161 ;
	7'h1c :
		rl_a64_t8 = RG_rl_161 ;
	7'h1d :
		rl_a64_t8 = RG_rl_161 ;
	7'h1e :
		rl_a64_t8 = RG_rl_161 ;
	7'h1f :
		rl_a64_t8 = RG_rl_161 ;
	7'h20 :
		rl_a64_t8 = RG_rl_161 ;
	7'h21 :
		rl_a64_t8 = RG_rl_161 ;
	7'h22 :
		rl_a64_t8 = RG_rl_161 ;
	7'h23 :
		rl_a64_t8 = RG_rl_161 ;
	7'h24 :
		rl_a64_t8 = RG_rl_161 ;
	7'h25 :
		rl_a64_t8 = RG_rl_161 ;
	7'h26 :
		rl_a64_t8 = RG_rl_161 ;
	7'h27 :
		rl_a64_t8 = RG_rl_161 ;
	7'h28 :
		rl_a64_t8 = RG_rl_161 ;
	7'h29 :
		rl_a64_t8 = RG_rl_161 ;
	7'h2a :
		rl_a64_t8 = RG_rl_161 ;
	7'h2b :
		rl_a64_t8 = RG_rl_161 ;
	7'h2c :
		rl_a64_t8 = RG_rl_161 ;
	7'h2d :
		rl_a64_t8 = RG_rl_161 ;
	7'h2e :
		rl_a64_t8 = RG_rl_161 ;
	7'h2f :
		rl_a64_t8 = RG_rl_161 ;
	7'h30 :
		rl_a64_t8 = RG_rl_161 ;
	7'h31 :
		rl_a64_t8 = RG_rl_161 ;
	7'h32 :
		rl_a64_t8 = RG_rl_161 ;
	7'h33 :
		rl_a64_t8 = RG_rl_161 ;
	7'h34 :
		rl_a64_t8 = RG_rl_161 ;
	7'h35 :
		rl_a64_t8 = RG_rl_161 ;
	7'h36 :
		rl_a64_t8 = RG_rl_161 ;
	7'h37 :
		rl_a64_t8 = RG_rl_161 ;
	7'h38 :
		rl_a64_t8 = RG_rl_161 ;
	7'h39 :
		rl_a64_t8 = RG_rl_161 ;
	7'h3a :
		rl_a64_t8 = RG_rl_161 ;
	7'h3b :
		rl_a64_t8 = RG_rl_161 ;
	7'h3c :
		rl_a64_t8 = RG_rl_161 ;
	7'h3d :
		rl_a64_t8 = RG_rl_161 ;
	7'h3e :
		rl_a64_t8 = RG_rl_161 ;
	7'h3f :
		rl_a64_t8 = RG_rl_161 ;
	7'h40 :
		rl_a64_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h41 :
		rl_a64_t8 = RG_rl_161 ;
	7'h42 :
		rl_a64_t8 = RG_rl_161 ;
	7'h43 :
		rl_a64_t8 = RG_rl_161 ;
	7'h44 :
		rl_a64_t8 = RG_rl_161 ;
	7'h45 :
		rl_a64_t8 = RG_rl_161 ;
	7'h46 :
		rl_a64_t8 = RG_rl_161 ;
	7'h47 :
		rl_a64_t8 = RG_rl_161 ;
	7'h48 :
		rl_a64_t8 = RG_rl_161 ;
	7'h49 :
		rl_a64_t8 = RG_rl_161 ;
	7'h4a :
		rl_a64_t8 = RG_rl_161 ;
	7'h4b :
		rl_a64_t8 = RG_rl_161 ;
	7'h4c :
		rl_a64_t8 = RG_rl_161 ;
	7'h4d :
		rl_a64_t8 = RG_rl_161 ;
	7'h4e :
		rl_a64_t8 = RG_rl_161 ;
	7'h4f :
		rl_a64_t8 = RG_rl_161 ;
	7'h50 :
		rl_a64_t8 = RG_rl_161 ;
	7'h51 :
		rl_a64_t8 = RG_rl_161 ;
	7'h52 :
		rl_a64_t8 = RG_rl_161 ;
	7'h53 :
		rl_a64_t8 = RG_rl_161 ;
	7'h54 :
		rl_a64_t8 = RG_rl_161 ;
	7'h55 :
		rl_a64_t8 = RG_rl_161 ;
	7'h56 :
		rl_a64_t8 = RG_rl_161 ;
	7'h57 :
		rl_a64_t8 = RG_rl_161 ;
	7'h58 :
		rl_a64_t8 = RG_rl_161 ;
	7'h59 :
		rl_a64_t8 = RG_rl_161 ;
	7'h5a :
		rl_a64_t8 = RG_rl_161 ;
	7'h5b :
		rl_a64_t8 = RG_rl_161 ;
	7'h5c :
		rl_a64_t8 = RG_rl_161 ;
	7'h5d :
		rl_a64_t8 = RG_rl_161 ;
	7'h5e :
		rl_a64_t8 = RG_rl_161 ;
	7'h5f :
		rl_a64_t8 = RG_rl_161 ;
	7'h60 :
		rl_a64_t8 = RG_rl_161 ;
	7'h61 :
		rl_a64_t8 = RG_rl_161 ;
	7'h62 :
		rl_a64_t8 = RG_rl_161 ;
	7'h63 :
		rl_a64_t8 = RG_rl_161 ;
	7'h64 :
		rl_a64_t8 = RG_rl_161 ;
	7'h65 :
		rl_a64_t8 = RG_rl_161 ;
	7'h66 :
		rl_a64_t8 = RG_rl_161 ;
	7'h67 :
		rl_a64_t8 = RG_rl_161 ;
	7'h68 :
		rl_a64_t8 = RG_rl_161 ;
	7'h69 :
		rl_a64_t8 = RG_rl_161 ;
	7'h6a :
		rl_a64_t8 = RG_rl_161 ;
	7'h6b :
		rl_a64_t8 = RG_rl_161 ;
	7'h6c :
		rl_a64_t8 = RG_rl_161 ;
	7'h6d :
		rl_a64_t8 = RG_rl_161 ;
	7'h6e :
		rl_a64_t8 = RG_rl_161 ;
	7'h6f :
		rl_a64_t8 = RG_rl_161 ;
	7'h70 :
		rl_a64_t8 = RG_rl_161 ;
	7'h71 :
		rl_a64_t8 = RG_rl_161 ;
	7'h72 :
		rl_a64_t8 = RG_rl_161 ;
	7'h73 :
		rl_a64_t8 = RG_rl_161 ;
	7'h74 :
		rl_a64_t8 = RG_rl_161 ;
	7'h75 :
		rl_a64_t8 = RG_rl_161 ;
	7'h76 :
		rl_a64_t8 = RG_rl_161 ;
	7'h77 :
		rl_a64_t8 = RG_rl_161 ;
	7'h78 :
		rl_a64_t8 = RG_rl_161 ;
	7'h79 :
		rl_a64_t8 = RG_rl_161 ;
	7'h7a :
		rl_a64_t8 = RG_rl_161 ;
	7'h7b :
		rl_a64_t8 = RG_rl_161 ;
	7'h7c :
		rl_a64_t8 = RG_rl_161 ;
	7'h7d :
		rl_a64_t8 = RG_rl_161 ;
	7'h7e :
		rl_a64_t8 = RG_rl_161 ;
	7'h7f :
		rl_a64_t8 = RG_rl_161 ;
	default :
		rl_a64_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_30 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h01 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h02 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h03 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h04 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h05 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h06 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h07 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h08 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h09 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h0a :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h0b :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h0c :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h0d :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h0e :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h0f :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h10 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h11 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h12 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h13 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h14 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h15 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h16 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h17 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h18 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h19 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h1a :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h1b :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h1c :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h1d :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h1e :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h1f :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h20 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h21 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h22 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h23 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h24 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h25 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h26 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h27 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h28 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h29 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h2a :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h2b :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h2c :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h2d :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h2e :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h2f :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h30 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h31 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h32 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h33 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h34 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h35 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h36 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h37 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h38 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h39 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h3a :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h3b :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h3c :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h3d :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h3e :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h3f :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h40 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h41 :
		rl_a65_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h42 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h43 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h44 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h45 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h46 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h47 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h48 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h49 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h4a :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h4b :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h4c :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h4d :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h4e :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h4f :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h50 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h51 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h52 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h53 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h54 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h55 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h56 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h57 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h58 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h59 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h5a :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h5b :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h5c :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h5d :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h5e :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h5f :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h60 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h61 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h62 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h63 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h64 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h65 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h66 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h67 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h68 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h69 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h6a :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h6b :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h6c :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h6d :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h6e :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h6f :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h70 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h71 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h72 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h73 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h74 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h75 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h76 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h77 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h78 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h79 :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h7a :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h7b :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h7c :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h7d :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h7e :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	7'h7f :
		rl_a65_t8 = RG_quantized_block_rl_30 ;
	default :
		rl_a65_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_162 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a66_t8 = RG_rl_162 ;
	7'h01 :
		rl_a66_t8 = RG_rl_162 ;
	7'h02 :
		rl_a66_t8 = RG_rl_162 ;
	7'h03 :
		rl_a66_t8 = RG_rl_162 ;
	7'h04 :
		rl_a66_t8 = RG_rl_162 ;
	7'h05 :
		rl_a66_t8 = RG_rl_162 ;
	7'h06 :
		rl_a66_t8 = RG_rl_162 ;
	7'h07 :
		rl_a66_t8 = RG_rl_162 ;
	7'h08 :
		rl_a66_t8 = RG_rl_162 ;
	7'h09 :
		rl_a66_t8 = RG_rl_162 ;
	7'h0a :
		rl_a66_t8 = RG_rl_162 ;
	7'h0b :
		rl_a66_t8 = RG_rl_162 ;
	7'h0c :
		rl_a66_t8 = RG_rl_162 ;
	7'h0d :
		rl_a66_t8 = RG_rl_162 ;
	7'h0e :
		rl_a66_t8 = RG_rl_162 ;
	7'h0f :
		rl_a66_t8 = RG_rl_162 ;
	7'h10 :
		rl_a66_t8 = RG_rl_162 ;
	7'h11 :
		rl_a66_t8 = RG_rl_162 ;
	7'h12 :
		rl_a66_t8 = RG_rl_162 ;
	7'h13 :
		rl_a66_t8 = RG_rl_162 ;
	7'h14 :
		rl_a66_t8 = RG_rl_162 ;
	7'h15 :
		rl_a66_t8 = RG_rl_162 ;
	7'h16 :
		rl_a66_t8 = RG_rl_162 ;
	7'h17 :
		rl_a66_t8 = RG_rl_162 ;
	7'h18 :
		rl_a66_t8 = RG_rl_162 ;
	7'h19 :
		rl_a66_t8 = RG_rl_162 ;
	7'h1a :
		rl_a66_t8 = RG_rl_162 ;
	7'h1b :
		rl_a66_t8 = RG_rl_162 ;
	7'h1c :
		rl_a66_t8 = RG_rl_162 ;
	7'h1d :
		rl_a66_t8 = RG_rl_162 ;
	7'h1e :
		rl_a66_t8 = RG_rl_162 ;
	7'h1f :
		rl_a66_t8 = RG_rl_162 ;
	7'h20 :
		rl_a66_t8 = RG_rl_162 ;
	7'h21 :
		rl_a66_t8 = RG_rl_162 ;
	7'h22 :
		rl_a66_t8 = RG_rl_162 ;
	7'h23 :
		rl_a66_t8 = RG_rl_162 ;
	7'h24 :
		rl_a66_t8 = RG_rl_162 ;
	7'h25 :
		rl_a66_t8 = RG_rl_162 ;
	7'h26 :
		rl_a66_t8 = RG_rl_162 ;
	7'h27 :
		rl_a66_t8 = RG_rl_162 ;
	7'h28 :
		rl_a66_t8 = RG_rl_162 ;
	7'h29 :
		rl_a66_t8 = RG_rl_162 ;
	7'h2a :
		rl_a66_t8 = RG_rl_162 ;
	7'h2b :
		rl_a66_t8 = RG_rl_162 ;
	7'h2c :
		rl_a66_t8 = RG_rl_162 ;
	7'h2d :
		rl_a66_t8 = RG_rl_162 ;
	7'h2e :
		rl_a66_t8 = RG_rl_162 ;
	7'h2f :
		rl_a66_t8 = RG_rl_162 ;
	7'h30 :
		rl_a66_t8 = RG_rl_162 ;
	7'h31 :
		rl_a66_t8 = RG_rl_162 ;
	7'h32 :
		rl_a66_t8 = RG_rl_162 ;
	7'h33 :
		rl_a66_t8 = RG_rl_162 ;
	7'h34 :
		rl_a66_t8 = RG_rl_162 ;
	7'h35 :
		rl_a66_t8 = RG_rl_162 ;
	7'h36 :
		rl_a66_t8 = RG_rl_162 ;
	7'h37 :
		rl_a66_t8 = RG_rl_162 ;
	7'h38 :
		rl_a66_t8 = RG_rl_162 ;
	7'h39 :
		rl_a66_t8 = RG_rl_162 ;
	7'h3a :
		rl_a66_t8 = RG_rl_162 ;
	7'h3b :
		rl_a66_t8 = RG_rl_162 ;
	7'h3c :
		rl_a66_t8 = RG_rl_162 ;
	7'h3d :
		rl_a66_t8 = RG_rl_162 ;
	7'h3e :
		rl_a66_t8 = RG_rl_162 ;
	7'h3f :
		rl_a66_t8 = RG_rl_162 ;
	7'h40 :
		rl_a66_t8 = RG_rl_162 ;
	7'h41 :
		rl_a66_t8 = RG_rl_162 ;
	7'h42 :
		rl_a66_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h43 :
		rl_a66_t8 = RG_rl_162 ;
	7'h44 :
		rl_a66_t8 = RG_rl_162 ;
	7'h45 :
		rl_a66_t8 = RG_rl_162 ;
	7'h46 :
		rl_a66_t8 = RG_rl_162 ;
	7'h47 :
		rl_a66_t8 = RG_rl_162 ;
	7'h48 :
		rl_a66_t8 = RG_rl_162 ;
	7'h49 :
		rl_a66_t8 = RG_rl_162 ;
	7'h4a :
		rl_a66_t8 = RG_rl_162 ;
	7'h4b :
		rl_a66_t8 = RG_rl_162 ;
	7'h4c :
		rl_a66_t8 = RG_rl_162 ;
	7'h4d :
		rl_a66_t8 = RG_rl_162 ;
	7'h4e :
		rl_a66_t8 = RG_rl_162 ;
	7'h4f :
		rl_a66_t8 = RG_rl_162 ;
	7'h50 :
		rl_a66_t8 = RG_rl_162 ;
	7'h51 :
		rl_a66_t8 = RG_rl_162 ;
	7'h52 :
		rl_a66_t8 = RG_rl_162 ;
	7'h53 :
		rl_a66_t8 = RG_rl_162 ;
	7'h54 :
		rl_a66_t8 = RG_rl_162 ;
	7'h55 :
		rl_a66_t8 = RG_rl_162 ;
	7'h56 :
		rl_a66_t8 = RG_rl_162 ;
	7'h57 :
		rl_a66_t8 = RG_rl_162 ;
	7'h58 :
		rl_a66_t8 = RG_rl_162 ;
	7'h59 :
		rl_a66_t8 = RG_rl_162 ;
	7'h5a :
		rl_a66_t8 = RG_rl_162 ;
	7'h5b :
		rl_a66_t8 = RG_rl_162 ;
	7'h5c :
		rl_a66_t8 = RG_rl_162 ;
	7'h5d :
		rl_a66_t8 = RG_rl_162 ;
	7'h5e :
		rl_a66_t8 = RG_rl_162 ;
	7'h5f :
		rl_a66_t8 = RG_rl_162 ;
	7'h60 :
		rl_a66_t8 = RG_rl_162 ;
	7'h61 :
		rl_a66_t8 = RG_rl_162 ;
	7'h62 :
		rl_a66_t8 = RG_rl_162 ;
	7'h63 :
		rl_a66_t8 = RG_rl_162 ;
	7'h64 :
		rl_a66_t8 = RG_rl_162 ;
	7'h65 :
		rl_a66_t8 = RG_rl_162 ;
	7'h66 :
		rl_a66_t8 = RG_rl_162 ;
	7'h67 :
		rl_a66_t8 = RG_rl_162 ;
	7'h68 :
		rl_a66_t8 = RG_rl_162 ;
	7'h69 :
		rl_a66_t8 = RG_rl_162 ;
	7'h6a :
		rl_a66_t8 = RG_rl_162 ;
	7'h6b :
		rl_a66_t8 = RG_rl_162 ;
	7'h6c :
		rl_a66_t8 = RG_rl_162 ;
	7'h6d :
		rl_a66_t8 = RG_rl_162 ;
	7'h6e :
		rl_a66_t8 = RG_rl_162 ;
	7'h6f :
		rl_a66_t8 = RG_rl_162 ;
	7'h70 :
		rl_a66_t8 = RG_rl_162 ;
	7'h71 :
		rl_a66_t8 = RG_rl_162 ;
	7'h72 :
		rl_a66_t8 = RG_rl_162 ;
	7'h73 :
		rl_a66_t8 = RG_rl_162 ;
	7'h74 :
		rl_a66_t8 = RG_rl_162 ;
	7'h75 :
		rl_a66_t8 = RG_rl_162 ;
	7'h76 :
		rl_a66_t8 = RG_rl_162 ;
	7'h77 :
		rl_a66_t8 = RG_rl_162 ;
	7'h78 :
		rl_a66_t8 = RG_rl_162 ;
	7'h79 :
		rl_a66_t8 = RG_rl_162 ;
	7'h7a :
		rl_a66_t8 = RG_rl_162 ;
	7'h7b :
		rl_a66_t8 = RG_rl_162 ;
	7'h7c :
		rl_a66_t8 = RG_rl_162 ;
	7'h7d :
		rl_a66_t8 = RG_rl_162 ;
	7'h7e :
		rl_a66_t8 = RG_rl_162 ;
	7'h7f :
		rl_a66_t8 = RG_rl_162 ;
	default :
		rl_a66_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_31 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h01 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h02 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h03 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h04 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h05 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h06 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h07 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h08 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h09 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h0a :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h0b :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h0c :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h0d :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h0e :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h0f :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h10 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h11 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h12 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h13 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h14 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h15 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h16 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h17 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h18 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h19 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h1a :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h1b :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h1c :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h1d :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h1e :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h1f :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h20 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h21 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h22 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h23 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h24 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h25 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h26 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h27 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h28 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h29 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h2a :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h2b :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h2c :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h2d :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h2e :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h2f :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h30 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h31 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h32 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h33 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h34 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h35 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h36 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h37 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h38 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h39 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h3a :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h3b :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h3c :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h3d :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h3e :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h3f :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h40 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h41 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h42 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h43 :
		rl_a67_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h44 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h45 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h46 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h47 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h48 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h49 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h4a :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h4b :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h4c :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h4d :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h4e :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h4f :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h50 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h51 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h52 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h53 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h54 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h55 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h56 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h57 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h58 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h59 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h5a :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h5b :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h5c :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h5d :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h5e :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h5f :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h60 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h61 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h62 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h63 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h64 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h65 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h66 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h67 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h68 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h69 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h6a :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h6b :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h6c :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h6d :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h6e :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h6f :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h70 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h71 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h72 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h73 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h74 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h75 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h76 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h77 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h78 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h79 :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h7a :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h7b :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h7c :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h7d :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h7e :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	7'h7f :
		rl_a67_t8 = RG_quantized_block_rl_31 ;
	default :
		rl_a67_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_163 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a68_t8 = RG_rl_163 ;
	7'h01 :
		rl_a68_t8 = RG_rl_163 ;
	7'h02 :
		rl_a68_t8 = RG_rl_163 ;
	7'h03 :
		rl_a68_t8 = RG_rl_163 ;
	7'h04 :
		rl_a68_t8 = RG_rl_163 ;
	7'h05 :
		rl_a68_t8 = RG_rl_163 ;
	7'h06 :
		rl_a68_t8 = RG_rl_163 ;
	7'h07 :
		rl_a68_t8 = RG_rl_163 ;
	7'h08 :
		rl_a68_t8 = RG_rl_163 ;
	7'h09 :
		rl_a68_t8 = RG_rl_163 ;
	7'h0a :
		rl_a68_t8 = RG_rl_163 ;
	7'h0b :
		rl_a68_t8 = RG_rl_163 ;
	7'h0c :
		rl_a68_t8 = RG_rl_163 ;
	7'h0d :
		rl_a68_t8 = RG_rl_163 ;
	7'h0e :
		rl_a68_t8 = RG_rl_163 ;
	7'h0f :
		rl_a68_t8 = RG_rl_163 ;
	7'h10 :
		rl_a68_t8 = RG_rl_163 ;
	7'h11 :
		rl_a68_t8 = RG_rl_163 ;
	7'h12 :
		rl_a68_t8 = RG_rl_163 ;
	7'h13 :
		rl_a68_t8 = RG_rl_163 ;
	7'h14 :
		rl_a68_t8 = RG_rl_163 ;
	7'h15 :
		rl_a68_t8 = RG_rl_163 ;
	7'h16 :
		rl_a68_t8 = RG_rl_163 ;
	7'h17 :
		rl_a68_t8 = RG_rl_163 ;
	7'h18 :
		rl_a68_t8 = RG_rl_163 ;
	7'h19 :
		rl_a68_t8 = RG_rl_163 ;
	7'h1a :
		rl_a68_t8 = RG_rl_163 ;
	7'h1b :
		rl_a68_t8 = RG_rl_163 ;
	7'h1c :
		rl_a68_t8 = RG_rl_163 ;
	7'h1d :
		rl_a68_t8 = RG_rl_163 ;
	7'h1e :
		rl_a68_t8 = RG_rl_163 ;
	7'h1f :
		rl_a68_t8 = RG_rl_163 ;
	7'h20 :
		rl_a68_t8 = RG_rl_163 ;
	7'h21 :
		rl_a68_t8 = RG_rl_163 ;
	7'h22 :
		rl_a68_t8 = RG_rl_163 ;
	7'h23 :
		rl_a68_t8 = RG_rl_163 ;
	7'h24 :
		rl_a68_t8 = RG_rl_163 ;
	7'h25 :
		rl_a68_t8 = RG_rl_163 ;
	7'h26 :
		rl_a68_t8 = RG_rl_163 ;
	7'h27 :
		rl_a68_t8 = RG_rl_163 ;
	7'h28 :
		rl_a68_t8 = RG_rl_163 ;
	7'h29 :
		rl_a68_t8 = RG_rl_163 ;
	7'h2a :
		rl_a68_t8 = RG_rl_163 ;
	7'h2b :
		rl_a68_t8 = RG_rl_163 ;
	7'h2c :
		rl_a68_t8 = RG_rl_163 ;
	7'h2d :
		rl_a68_t8 = RG_rl_163 ;
	7'h2e :
		rl_a68_t8 = RG_rl_163 ;
	7'h2f :
		rl_a68_t8 = RG_rl_163 ;
	7'h30 :
		rl_a68_t8 = RG_rl_163 ;
	7'h31 :
		rl_a68_t8 = RG_rl_163 ;
	7'h32 :
		rl_a68_t8 = RG_rl_163 ;
	7'h33 :
		rl_a68_t8 = RG_rl_163 ;
	7'h34 :
		rl_a68_t8 = RG_rl_163 ;
	7'h35 :
		rl_a68_t8 = RG_rl_163 ;
	7'h36 :
		rl_a68_t8 = RG_rl_163 ;
	7'h37 :
		rl_a68_t8 = RG_rl_163 ;
	7'h38 :
		rl_a68_t8 = RG_rl_163 ;
	7'h39 :
		rl_a68_t8 = RG_rl_163 ;
	7'h3a :
		rl_a68_t8 = RG_rl_163 ;
	7'h3b :
		rl_a68_t8 = RG_rl_163 ;
	7'h3c :
		rl_a68_t8 = RG_rl_163 ;
	7'h3d :
		rl_a68_t8 = RG_rl_163 ;
	7'h3e :
		rl_a68_t8 = RG_rl_163 ;
	7'h3f :
		rl_a68_t8 = RG_rl_163 ;
	7'h40 :
		rl_a68_t8 = RG_rl_163 ;
	7'h41 :
		rl_a68_t8 = RG_rl_163 ;
	7'h42 :
		rl_a68_t8 = RG_rl_163 ;
	7'h43 :
		rl_a68_t8 = RG_rl_163 ;
	7'h44 :
		rl_a68_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h45 :
		rl_a68_t8 = RG_rl_163 ;
	7'h46 :
		rl_a68_t8 = RG_rl_163 ;
	7'h47 :
		rl_a68_t8 = RG_rl_163 ;
	7'h48 :
		rl_a68_t8 = RG_rl_163 ;
	7'h49 :
		rl_a68_t8 = RG_rl_163 ;
	7'h4a :
		rl_a68_t8 = RG_rl_163 ;
	7'h4b :
		rl_a68_t8 = RG_rl_163 ;
	7'h4c :
		rl_a68_t8 = RG_rl_163 ;
	7'h4d :
		rl_a68_t8 = RG_rl_163 ;
	7'h4e :
		rl_a68_t8 = RG_rl_163 ;
	7'h4f :
		rl_a68_t8 = RG_rl_163 ;
	7'h50 :
		rl_a68_t8 = RG_rl_163 ;
	7'h51 :
		rl_a68_t8 = RG_rl_163 ;
	7'h52 :
		rl_a68_t8 = RG_rl_163 ;
	7'h53 :
		rl_a68_t8 = RG_rl_163 ;
	7'h54 :
		rl_a68_t8 = RG_rl_163 ;
	7'h55 :
		rl_a68_t8 = RG_rl_163 ;
	7'h56 :
		rl_a68_t8 = RG_rl_163 ;
	7'h57 :
		rl_a68_t8 = RG_rl_163 ;
	7'h58 :
		rl_a68_t8 = RG_rl_163 ;
	7'h59 :
		rl_a68_t8 = RG_rl_163 ;
	7'h5a :
		rl_a68_t8 = RG_rl_163 ;
	7'h5b :
		rl_a68_t8 = RG_rl_163 ;
	7'h5c :
		rl_a68_t8 = RG_rl_163 ;
	7'h5d :
		rl_a68_t8 = RG_rl_163 ;
	7'h5e :
		rl_a68_t8 = RG_rl_163 ;
	7'h5f :
		rl_a68_t8 = RG_rl_163 ;
	7'h60 :
		rl_a68_t8 = RG_rl_163 ;
	7'h61 :
		rl_a68_t8 = RG_rl_163 ;
	7'h62 :
		rl_a68_t8 = RG_rl_163 ;
	7'h63 :
		rl_a68_t8 = RG_rl_163 ;
	7'h64 :
		rl_a68_t8 = RG_rl_163 ;
	7'h65 :
		rl_a68_t8 = RG_rl_163 ;
	7'h66 :
		rl_a68_t8 = RG_rl_163 ;
	7'h67 :
		rl_a68_t8 = RG_rl_163 ;
	7'h68 :
		rl_a68_t8 = RG_rl_163 ;
	7'h69 :
		rl_a68_t8 = RG_rl_163 ;
	7'h6a :
		rl_a68_t8 = RG_rl_163 ;
	7'h6b :
		rl_a68_t8 = RG_rl_163 ;
	7'h6c :
		rl_a68_t8 = RG_rl_163 ;
	7'h6d :
		rl_a68_t8 = RG_rl_163 ;
	7'h6e :
		rl_a68_t8 = RG_rl_163 ;
	7'h6f :
		rl_a68_t8 = RG_rl_163 ;
	7'h70 :
		rl_a68_t8 = RG_rl_163 ;
	7'h71 :
		rl_a68_t8 = RG_rl_163 ;
	7'h72 :
		rl_a68_t8 = RG_rl_163 ;
	7'h73 :
		rl_a68_t8 = RG_rl_163 ;
	7'h74 :
		rl_a68_t8 = RG_rl_163 ;
	7'h75 :
		rl_a68_t8 = RG_rl_163 ;
	7'h76 :
		rl_a68_t8 = RG_rl_163 ;
	7'h77 :
		rl_a68_t8 = RG_rl_163 ;
	7'h78 :
		rl_a68_t8 = RG_rl_163 ;
	7'h79 :
		rl_a68_t8 = RG_rl_163 ;
	7'h7a :
		rl_a68_t8 = RG_rl_163 ;
	7'h7b :
		rl_a68_t8 = RG_rl_163 ;
	7'h7c :
		rl_a68_t8 = RG_rl_163 ;
	7'h7d :
		rl_a68_t8 = RG_rl_163 ;
	7'h7e :
		rl_a68_t8 = RG_rl_163 ;
	7'h7f :
		rl_a68_t8 = RG_rl_163 ;
	default :
		rl_a68_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_32 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h01 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h02 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h03 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h04 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h05 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h06 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h07 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h08 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h09 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h0a :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h0b :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h0c :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h0d :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h0e :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h0f :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h10 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h11 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h12 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h13 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h14 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h15 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h16 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h17 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h18 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h19 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h1a :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h1b :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h1c :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h1d :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h1e :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h1f :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h20 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h21 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h22 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h23 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h24 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h25 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h26 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h27 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h28 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h29 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h2a :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h2b :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h2c :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h2d :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h2e :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h2f :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h30 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h31 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h32 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h33 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h34 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h35 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h36 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h37 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h38 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h39 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h3a :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h3b :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h3c :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h3d :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h3e :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h3f :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h40 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h41 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h42 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h43 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h44 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h45 :
		rl_a69_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h46 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h47 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h48 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h49 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h4a :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h4b :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h4c :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h4d :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h4e :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h4f :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h50 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h51 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h52 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h53 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h54 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h55 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h56 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h57 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h58 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h59 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h5a :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h5b :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h5c :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h5d :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h5e :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h5f :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h60 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h61 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h62 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h63 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h64 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h65 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h66 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h67 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h68 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h69 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h6a :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h6b :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h6c :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h6d :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h6e :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h6f :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h70 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h71 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h72 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h73 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h74 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h75 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h76 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h77 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h78 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h79 :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h7a :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h7b :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h7c :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h7d :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h7e :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	7'h7f :
		rl_a69_t8 = RG_quantized_block_rl_32 ;
	default :
		rl_a69_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_164 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a70_t8 = RG_rl_164 ;
	7'h01 :
		rl_a70_t8 = RG_rl_164 ;
	7'h02 :
		rl_a70_t8 = RG_rl_164 ;
	7'h03 :
		rl_a70_t8 = RG_rl_164 ;
	7'h04 :
		rl_a70_t8 = RG_rl_164 ;
	7'h05 :
		rl_a70_t8 = RG_rl_164 ;
	7'h06 :
		rl_a70_t8 = RG_rl_164 ;
	7'h07 :
		rl_a70_t8 = RG_rl_164 ;
	7'h08 :
		rl_a70_t8 = RG_rl_164 ;
	7'h09 :
		rl_a70_t8 = RG_rl_164 ;
	7'h0a :
		rl_a70_t8 = RG_rl_164 ;
	7'h0b :
		rl_a70_t8 = RG_rl_164 ;
	7'h0c :
		rl_a70_t8 = RG_rl_164 ;
	7'h0d :
		rl_a70_t8 = RG_rl_164 ;
	7'h0e :
		rl_a70_t8 = RG_rl_164 ;
	7'h0f :
		rl_a70_t8 = RG_rl_164 ;
	7'h10 :
		rl_a70_t8 = RG_rl_164 ;
	7'h11 :
		rl_a70_t8 = RG_rl_164 ;
	7'h12 :
		rl_a70_t8 = RG_rl_164 ;
	7'h13 :
		rl_a70_t8 = RG_rl_164 ;
	7'h14 :
		rl_a70_t8 = RG_rl_164 ;
	7'h15 :
		rl_a70_t8 = RG_rl_164 ;
	7'h16 :
		rl_a70_t8 = RG_rl_164 ;
	7'h17 :
		rl_a70_t8 = RG_rl_164 ;
	7'h18 :
		rl_a70_t8 = RG_rl_164 ;
	7'h19 :
		rl_a70_t8 = RG_rl_164 ;
	7'h1a :
		rl_a70_t8 = RG_rl_164 ;
	7'h1b :
		rl_a70_t8 = RG_rl_164 ;
	7'h1c :
		rl_a70_t8 = RG_rl_164 ;
	7'h1d :
		rl_a70_t8 = RG_rl_164 ;
	7'h1e :
		rl_a70_t8 = RG_rl_164 ;
	7'h1f :
		rl_a70_t8 = RG_rl_164 ;
	7'h20 :
		rl_a70_t8 = RG_rl_164 ;
	7'h21 :
		rl_a70_t8 = RG_rl_164 ;
	7'h22 :
		rl_a70_t8 = RG_rl_164 ;
	7'h23 :
		rl_a70_t8 = RG_rl_164 ;
	7'h24 :
		rl_a70_t8 = RG_rl_164 ;
	7'h25 :
		rl_a70_t8 = RG_rl_164 ;
	7'h26 :
		rl_a70_t8 = RG_rl_164 ;
	7'h27 :
		rl_a70_t8 = RG_rl_164 ;
	7'h28 :
		rl_a70_t8 = RG_rl_164 ;
	7'h29 :
		rl_a70_t8 = RG_rl_164 ;
	7'h2a :
		rl_a70_t8 = RG_rl_164 ;
	7'h2b :
		rl_a70_t8 = RG_rl_164 ;
	7'h2c :
		rl_a70_t8 = RG_rl_164 ;
	7'h2d :
		rl_a70_t8 = RG_rl_164 ;
	7'h2e :
		rl_a70_t8 = RG_rl_164 ;
	7'h2f :
		rl_a70_t8 = RG_rl_164 ;
	7'h30 :
		rl_a70_t8 = RG_rl_164 ;
	7'h31 :
		rl_a70_t8 = RG_rl_164 ;
	7'h32 :
		rl_a70_t8 = RG_rl_164 ;
	7'h33 :
		rl_a70_t8 = RG_rl_164 ;
	7'h34 :
		rl_a70_t8 = RG_rl_164 ;
	7'h35 :
		rl_a70_t8 = RG_rl_164 ;
	7'h36 :
		rl_a70_t8 = RG_rl_164 ;
	7'h37 :
		rl_a70_t8 = RG_rl_164 ;
	7'h38 :
		rl_a70_t8 = RG_rl_164 ;
	7'h39 :
		rl_a70_t8 = RG_rl_164 ;
	7'h3a :
		rl_a70_t8 = RG_rl_164 ;
	7'h3b :
		rl_a70_t8 = RG_rl_164 ;
	7'h3c :
		rl_a70_t8 = RG_rl_164 ;
	7'h3d :
		rl_a70_t8 = RG_rl_164 ;
	7'h3e :
		rl_a70_t8 = RG_rl_164 ;
	7'h3f :
		rl_a70_t8 = RG_rl_164 ;
	7'h40 :
		rl_a70_t8 = RG_rl_164 ;
	7'h41 :
		rl_a70_t8 = RG_rl_164 ;
	7'h42 :
		rl_a70_t8 = RG_rl_164 ;
	7'h43 :
		rl_a70_t8 = RG_rl_164 ;
	7'h44 :
		rl_a70_t8 = RG_rl_164 ;
	7'h45 :
		rl_a70_t8 = RG_rl_164 ;
	7'h46 :
		rl_a70_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h47 :
		rl_a70_t8 = RG_rl_164 ;
	7'h48 :
		rl_a70_t8 = RG_rl_164 ;
	7'h49 :
		rl_a70_t8 = RG_rl_164 ;
	7'h4a :
		rl_a70_t8 = RG_rl_164 ;
	7'h4b :
		rl_a70_t8 = RG_rl_164 ;
	7'h4c :
		rl_a70_t8 = RG_rl_164 ;
	7'h4d :
		rl_a70_t8 = RG_rl_164 ;
	7'h4e :
		rl_a70_t8 = RG_rl_164 ;
	7'h4f :
		rl_a70_t8 = RG_rl_164 ;
	7'h50 :
		rl_a70_t8 = RG_rl_164 ;
	7'h51 :
		rl_a70_t8 = RG_rl_164 ;
	7'h52 :
		rl_a70_t8 = RG_rl_164 ;
	7'h53 :
		rl_a70_t8 = RG_rl_164 ;
	7'h54 :
		rl_a70_t8 = RG_rl_164 ;
	7'h55 :
		rl_a70_t8 = RG_rl_164 ;
	7'h56 :
		rl_a70_t8 = RG_rl_164 ;
	7'h57 :
		rl_a70_t8 = RG_rl_164 ;
	7'h58 :
		rl_a70_t8 = RG_rl_164 ;
	7'h59 :
		rl_a70_t8 = RG_rl_164 ;
	7'h5a :
		rl_a70_t8 = RG_rl_164 ;
	7'h5b :
		rl_a70_t8 = RG_rl_164 ;
	7'h5c :
		rl_a70_t8 = RG_rl_164 ;
	7'h5d :
		rl_a70_t8 = RG_rl_164 ;
	7'h5e :
		rl_a70_t8 = RG_rl_164 ;
	7'h5f :
		rl_a70_t8 = RG_rl_164 ;
	7'h60 :
		rl_a70_t8 = RG_rl_164 ;
	7'h61 :
		rl_a70_t8 = RG_rl_164 ;
	7'h62 :
		rl_a70_t8 = RG_rl_164 ;
	7'h63 :
		rl_a70_t8 = RG_rl_164 ;
	7'h64 :
		rl_a70_t8 = RG_rl_164 ;
	7'h65 :
		rl_a70_t8 = RG_rl_164 ;
	7'h66 :
		rl_a70_t8 = RG_rl_164 ;
	7'h67 :
		rl_a70_t8 = RG_rl_164 ;
	7'h68 :
		rl_a70_t8 = RG_rl_164 ;
	7'h69 :
		rl_a70_t8 = RG_rl_164 ;
	7'h6a :
		rl_a70_t8 = RG_rl_164 ;
	7'h6b :
		rl_a70_t8 = RG_rl_164 ;
	7'h6c :
		rl_a70_t8 = RG_rl_164 ;
	7'h6d :
		rl_a70_t8 = RG_rl_164 ;
	7'h6e :
		rl_a70_t8 = RG_rl_164 ;
	7'h6f :
		rl_a70_t8 = RG_rl_164 ;
	7'h70 :
		rl_a70_t8 = RG_rl_164 ;
	7'h71 :
		rl_a70_t8 = RG_rl_164 ;
	7'h72 :
		rl_a70_t8 = RG_rl_164 ;
	7'h73 :
		rl_a70_t8 = RG_rl_164 ;
	7'h74 :
		rl_a70_t8 = RG_rl_164 ;
	7'h75 :
		rl_a70_t8 = RG_rl_164 ;
	7'h76 :
		rl_a70_t8 = RG_rl_164 ;
	7'h77 :
		rl_a70_t8 = RG_rl_164 ;
	7'h78 :
		rl_a70_t8 = RG_rl_164 ;
	7'h79 :
		rl_a70_t8 = RG_rl_164 ;
	7'h7a :
		rl_a70_t8 = RG_rl_164 ;
	7'h7b :
		rl_a70_t8 = RG_rl_164 ;
	7'h7c :
		rl_a70_t8 = RG_rl_164 ;
	7'h7d :
		rl_a70_t8 = RG_rl_164 ;
	7'h7e :
		rl_a70_t8 = RG_rl_164 ;
	7'h7f :
		rl_a70_t8 = RG_rl_164 ;
	default :
		rl_a70_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_33 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h01 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h02 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h03 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h04 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h05 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h06 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h07 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h08 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h09 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h0a :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h0b :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h0c :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h0d :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h0e :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h0f :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h10 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h11 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h12 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h13 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h14 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h15 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h16 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h17 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h18 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h19 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h1a :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h1b :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h1c :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h1d :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h1e :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h1f :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h20 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h21 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h22 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h23 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h24 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h25 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h26 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h27 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h28 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h29 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h2a :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h2b :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h2c :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h2d :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h2e :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h2f :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h30 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h31 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h32 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h33 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h34 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h35 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h36 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h37 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h38 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h39 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h3a :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h3b :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h3c :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h3d :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h3e :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h3f :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h40 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h41 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h42 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h43 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h44 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h45 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h46 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h47 :
		rl_a71_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h48 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h49 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h4a :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h4b :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h4c :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h4d :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h4e :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h4f :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h50 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h51 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h52 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h53 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h54 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h55 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h56 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h57 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h58 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h59 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h5a :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h5b :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h5c :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h5d :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h5e :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h5f :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h60 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h61 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h62 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h63 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h64 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h65 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h66 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h67 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h68 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h69 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h6a :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h6b :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h6c :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h6d :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h6e :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h6f :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h70 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h71 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h72 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h73 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h74 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h75 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h76 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h77 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h78 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h79 :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h7a :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h7b :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h7c :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h7d :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h7e :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	7'h7f :
		rl_a71_t8 = RG_quantized_block_rl_33 ;
	default :
		rl_a71_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_165 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a72_t8 = RG_rl_165 ;
	7'h01 :
		rl_a72_t8 = RG_rl_165 ;
	7'h02 :
		rl_a72_t8 = RG_rl_165 ;
	7'h03 :
		rl_a72_t8 = RG_rl_165 ;
	7'h04 :
		rl_a72_t8 = RG_rl_165 ;
	7'h05 :
		rl_a72_t8 = RG_rl_165 ;
	7'h06 :
		rl_a72_t8 = RG_rl_165 ;
	7'h07 :
		rl_a72_t8 = RG_rl_165 ;
	7'h08 :
		rl_a72_t8 = RG_rl_165 ;
	7'h09 :
		rl_a72_t8 = RG_rl_165 ;
	7'h0a :
		rl_a72_t8 = RG_rl_165 ;
	7'h0b :
		rl_a72_t8 = RG_rl_165 ;
	7'h0c :
		rl_a72_t8 = RG_rl_165 ;
	7'h0d :
		rl_a72_t8 = RG_rl_165 ;
	7'h0e :
		rl_a72_t8 = RG_rl_165 ;
	7'h0f :
		rl_a72_t8 = RG_rl_165 ;
	7'h10 :
		rl_a72_t8 = RG_rl_165 ;
	7'h11 :
		rl_a72_t8 = RG_rl_165 ;
	7'h12 :
		rl_a72_t8 = RG_rl_165 ;
	7'h13 :
		rl_a72_t8 = RG_rl_165 ;
	7'h14 :
		rl_a72_t8 = RG_rl_165 ;
	7'h15 :
		rl_a72_t8 = RG_rl_165 ;
	7'h16 :
		rl_a72_t8 = RG_rl_165 ;
	7'h17 :
		rl_a72_t8 = RG_rl_165 ;
	7'h18 :
		rl_a72_t8 = RG_rl_165 ;
	7'h19 :
		rl_a72_t8 = RG_rl_165 ;
	7'h1a :
		rl_a72_t8 = RG_rl_165 ;
	7'h1b :
		rl_a72_t8 = RG_rl_165 ;
	7'h1c :
		rl_a72_t8 = RG_rl_165 ;
	7'h1d :
		rl_a72_t8 = RG_rl_165 ;
	7'h1e :
		rl_a72_t8 = RG_rl_165 ;
	7'h1f :
		rl_a72_t8 = RG_rl_165 ;
	7'h20 :
		rl_a72_t8 = RG_rl_165 ;
	7'h21 :
		rl_a72_t8 = RG_rl_165 ;
	7'h22 :
		rl_a72_t8 = RG_rl_165 ;
	7'h23 :
		rl_a72_t8 = RG_rl_165 ;
	7'h24 :
		rl_a72_t8 = RG_rl_165 ;
	7'h25 :
		rl_a72_t8 = RG_rl_165 ;
	7'h26 :
		rl_a72_t8 = RG_rl_165 ;
	7'h27 :
		rl_a72_t8 = RG_rl_165 ;
	7'h28 :
		rl_a72_t8 = RG_rl_165 ;
	7'h29 :
		rl_a72_t8 = RG_rl_165 ;
	7'h2a :
		rl_a72_t8 = RG_rl_165 ;
	7'h2b :
		rl_a72_t8 = RG_rl_165 ;
	7'h2c :
		rl_a72_t8 = RG_rl_165 ;
	7'h2d :
		rl_a72_t8 = RG_rl_165 ;
	7'h2e :
		rl_a72_t8 = RG_rl_165 ;
	7'h2f :
		rl_a72_t8 = RG_rl_165 ;
	7'h30 :
		rl_a72_t8 = RG_rl_165 ;
	7'h31 :
		rl_a72_t8 = RG_rl_165 ;
	7'h32 :
		rl_a72_t8 = RG_rl_165 ;
	7'h33 :
		rl_a72_t8 = RG_rl_165 ;
	7'h34 :
		rl_a72_t8 = RG_rl_165 ;
	7'h35 :
		rl_a72_t8 = RG_rl_165 ;
	7'h36 :
		rl_a72_t8 = RG_rl_165 ;
	7'h37 :
		rl_a72_t8 = RG_rl_165 ;
	7'h38 :
		rl_a72_t8 = RG_rl_165 ;
	7'h39 :
		rl_a72_t8 = RG_rl_165 ;
	7'h3a :
		rl_a72_t8 = RG_rl_165 ;
	7'h3b :
		rl_a72_t8 = RG_rl_165 ;
	7'h3c :
		rl_a72_t8 = RG_rl_165 ;
	7'h3d :
		rl_a72_t8 = RG_rl_165 ;
	7'h3e :
		rl_a72_t8 = RG_rl_165 ;
	7'h3f :
		rl_a72_t8 = RG_rl_165 ;
	7'h40 :
		rl_a72_t8 = RG_rl_165 ;
	7'h41 :
		rl_a72_t8 = RG_rl_165 ;
	7'h42 :
		rl_a72_t8 = RG_rl_165 ;
	7'h43 :
		rl_a72_t8 = RG_rl_165 ;
	7'h44 :
		rl_a72_t8 = RG_rl_165 ;
	7'h45 :
		rl_a72_t8 = RG_rl_165 ;
	7'h46 :
		rl_a72_t8 = RG_rl_165 ;
	7'h47 :
		rl_a72_t8 = RG_rl_165 ;
	7'h48 :
		rl_a72_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h49 :
		rl_a72_t8 = RG_rl_165 ;
	7'h4a :
		rl_a72_t8 = RG_rl_165 ;
	7'h4b :
		rl_a72_t8 = RG_rl_165 ;
	7'h4c :
		rl_a72_t8 = RG_rl_165 ;
	7'h4d :
		rl_a72_t8 = RG_rl_165 ;
	7'h4e :
		rl_a72_t8 = RG_rl_165 ;
	7'h4f :
		rl_a72_t8 = RG_rl_165 ;
	7'h50 :
		rl_a72_t8 = RG_rl_165 ;
	7'h51 :
		rl_a72_t8 = RG_rl_165 ;
	7'h52 :
		rl_a72_t8 = RG_rl_165 ;
	7'h53 :
		rl_a72_t8 = RG_rl_165 ;
	7'h54 :
		rl_a72_t8 = RG_rl_165 ;
	7'h55 :
		rl_a72_t8 = RG_rl_165 ;
	7'h56 :
		rl_a72_t8 = RG_rl_165 ;
	7'h57 :
		rl_a72_t8 = RG_rl_165 ;
	7'h58 :
		rl_a72_t8 = RG_rl_165 ;
	7'h59 :
		rl_a72_t8 = RG_rl_165 ;
	7'h5a :
		rl_a72_t8 = RG_rl_165 ;
	7'h5b :
		rl_a72_t8 = RG_rl_165 ;
	7'h5c :
		rl_a72_t8 = RG_rl_165 ;
	7'h5d :
		rl_a72_t8 = RG_rl_165 ;
	7'h5e :
		rl_a72_t8 = RG_rl_165 ;
	7'h5f :
		rl_a72_t8 = RG_rl_165 ;
	7'h60 :
		rl_a72_t8 = RG_rl_165 ;
	7'h61 :
		rl_a72_t8 = RG_rl_165 ;
	7'h62 :
		rl_a72_t8 = RG_rl_165 ;
	7'h63 :
		rl_a72_t8 = RG_rl_165 ;
	7'h64 :
		rl_a72_t8 = RG_rl_165 ;
	7'h65 :
		rl_a72_t8 = RG_rl_165 ;
	7'h66 :
		rl_a72_t8 = RG_rl_165 ;
	7'h67 :
		rl_a72_t8 = RG_rl_165 ;
	7'h68 :
		rl_a72_t8 = RG_rl_165 ;
	7'h69 :
		rl_a72_t8 = RG_rl_165 ;
	7'h6a :
		rl_a72_t8 = RG_rl_165 ;
	7'h6b :
		rl_a72_t8 = RG_rl_165 ;
	7'h6c :
		rl_a72_t8 = RG_rl_165 ;
	7'h6d :
		rl_a72_t8 = RG_rl_165 ;
	7'h6e :
		rl_a72_t8 = RG_rl_165 ;
	7'h6f :
		rl_a72_t8 = RG_rl_165 ;
	7'h70 :
		rl_a72_t8 = RG_rl_165 ;
	7'h71 :
		rl_a72_t8 = RG_rl_165 ;
	7'h72 :
		rl_a72_t8 = RG_rl_165 ;
	7'h73 :
		rl_a72_t8 = RG_rl_165 ;
	7'h74 :
		rl_a72_t8 = RG_rl_165 ;
	7'h75 :
		rl_a72_t8 = RG_rl_165 ;
	7'h76 :
		rl_a72_t8 = RG_rl_165 ;
	7'h77 :
		rl_a72_t8 = RG_rl_165 ;
	7'h78 :
		rl_a72_t8 = RG_rl_165 ;
	7'h79 :
		rl_a72_t8 = RG_rl_165 ;
	7'h7a :
		rl_a72_t8 = RG_rl_165 ;
	7'h7b :
		rl_a72_t8 = RG_rl_165 ;
	7'h7c :
		rl_a72_t8 = RG_rl_165 ;
	7'h7d :
		rl_a72_t8 = RG_rl_165 ;
	7'h7e :
		rl_a72_t8 = RG_rl_165 ;
	7'h7f :
		rl_a72_t8 = RG_rl_165 ;
	default :
		rl_a72_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_34 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h01 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h02 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h03 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h04 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h05 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h06 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h07 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h08 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h09 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h0a :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h0b :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h0c :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h0d :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h0e :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h0f :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h10 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h11 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h12 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h13 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h14 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h15 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h16 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h17 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h18 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h19 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h1a :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h1b :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h1c :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h1d :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h1e :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h1f :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h20 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h21 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h22 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h23 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h24 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h25 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h26 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h27 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h28 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h29 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h2a :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h2b :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h2c :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h2d :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h2e :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h2f :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h30 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h31 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h32 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h33 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h34 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h35 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h36 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h37 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h38 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h39 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h3a :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h3b :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h3c :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h3d :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h3e :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h3f :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h40 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h41 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h42 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h43 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h44 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h45 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h46 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h47 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h48 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h49 :
		rl_a73_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h4a :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h4b :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h4c :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h4d :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h4e :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h4f :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h50 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h51 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h52 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h53 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h54 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h55 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h56 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h57 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h58 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h59 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h5a :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h5b :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h5c :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h5d :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h5e :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h5f :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h60 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h61 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h62 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h63 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h64 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h65 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h66 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h67 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h68 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h69 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h6a :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h6b :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h6c :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h6d :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h6e :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h6f :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h70 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h71 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h72 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h73 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h74 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h75 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h76 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h77 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h78 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h79 :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h7a :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h7b :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h7c :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h7d :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h7e :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	7'h7f :
		rl_a73_t8 = RG_quantized_block_rl_34 ;
	default :
		rl_a73_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_166 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a74_t8 = RG_rl_166 ;
	7'h01 :
		rl_a74_t8 = RG_rl_166 ;
	7'h02 :
		rl_a74_t8 = RG_rl_166 ;
	7'h03 :
		rl_a74_t8 = RG_rl_166 ;
	7'h04 :
		rl_a74_t8 = RG_rl_166 ;
	7'h05 :
		rl_a74_t8 = RG_rl_166 ;
	7'h06 :
		rl_a74_t8 = RG_rl_166 ;
	7'h07 :
		rl_a74_t8 = RG_rl_166 ;
	7'h08 :
		rl_a74_t8 = RG_rl_166 ;
	7'h09 :
		rl_a74_t8 = RG_rl_166 ;
	7'h0a :
		rl_a74_t8 = RG_rl_166 ;
	7'h0b :
		rl_a74_t8 = RG_rl_166 ;
	7'h0c :
		rl_a74_t8 = RG_rl_166 ;
	7'h0d :
		rl_a74_t8 = RG_rl_166 ;
	7'h0e :
		rl_a74_t8 = RG_rl_166 ;
	7'h0f :
		rl_a74_t8 = RG_rl_166 ;
	7'h10 :
		rl_a74_t8 = RG_rl_166 ;
	7'h11 :
		rl_a74_t8 = RG_rl_166 ;
	7'h12 :
		rl_a74_t8 = RG_rl_166 ;
	7'h13 :
		rl_a74_t8 = RG_rl_166 ;
	7'h14 :
		rl_a74_t8 = RG_rl_166 ;
	7'h15 :
		rl_a74_t8 = RG_rl_166 ;
	7'h16 :
		rl_a74_t8 = RG_rl_166 ;
	7'h17 :
		rl_a74_t8 = RG_rl_166 ;
	7'h18 :
		rl_a74_t8 = RG_rl_166 ;
	7'h19 :
		rl_a74_t8 = RG_rl_166 ;
	7'h1a :
		rl_a74_t8 = RG_rl_166 ;
	7'h1b :
		rl_a74_t8 = RG_rl_166 ;
	7'h1c :
		rl_a74_t8 = RG_rl_166 ;
	7'h1d :
		rl_a74_t8 = RG_rl_166 ;
	7'h1e :
		rl_a74_t8 = RG_rl_166 ;
	7'h1f :
		rl_a74_t8 = RG_rl_166 ;
	7'h20 :
		rl_a74_t8 = RG_rl_166 ;
	7'h21 :
		rl_a74_t8 = RG_rl_166 ;
	7'h22 :
		rl_a74_t8 = RG_rl_166 ;
	7'h23 :
		rl_a74_t8 = RG_rl_166 ;
	7'h24 :
		rl_a74_t8 = RG_rl_166 ;
	7'h25 :
		rl_a74_t8 = RG_rl_166 ;
	7'h26 :
		rl_a74_t8 = RG_rl_166 ;
	7'h27 :
		rl_a74_t8 = RG_rl_166 ;
	7'h28 :
		rl_a74_t8 = RG_rl_166 ;
	7'h29 :
		rl_a74_t8 = RG_rl_166 ;
	7'h2a :
		rl_a74_t8 = RG_rl_166 ;
	7'h2b :
		rl_a74_t8 = RG_rl_166 ;
	7'h2c :
		rl_a74_t8 = RG_rl_166 ;
	7'h2d :
		rl_a74_t8 = RG_rl_166 ;
	7'h2e :
		rl_a74_t8 = RG_rl_166 ;
	7'h2f :
		rl_a74_t8 = RG_rl_166 ;
	7'h30 :
		rl_a74_t8 = RG_rl_166 ;
	7'h31 :
		rl_a74_t8 = RG_rl_166 ;
	7'h32 :
		rl_a74_t8 = RG_rl_166 ;
	7'h33 :
		rl_a74_t8 = RG_rl_166 ;
	7'h34 :
		rl_a74_t8 = RG_rl_166 ;
	7'h35 :
		rl_a74_t8 = RG_rl_166 ;
	7'h36 :
		rl_a74_t8 = RG_rl_166 ;
	7'h37 :
		rl_a74_t8 = RG_rl_166 ;
	7'h38 :
		rl_a74_t8 = RG_rl_166 ;
	7'h39 :
		rl_a74_t8 = RG_rl_166 ;
	7'h3a :
		rl_a74_t8 = RG_rl_166 ;
	7'h3b :
		rl_a74_t8 = RG_rl_166 ;
	7'h3c :
		rl_a74_t8 = RG_rl_166 ;
	7'h3d :
		rl_a74_t8 = RG_rl_166 ;
	7'h3e :
		rl_a74_t8 = RG_rl_166 ;
	7'h3f :
		rl_a74_t8 = RG_rl_166 ;
	7'h40 :
		rl_a74_t8 = RG_rl_166 ;
	7'h41 :
		rl_a74_t8 = RG_rl_166 ;
	7'h42 :
		rl_a74_t8 = RG_rl_166 ;
	7'h43 :
		rl_a74_t8 = RG_rl_166 ;
	7'h44 :
		rl_a74_t8 = RG_rl_166 ;
	7'h45 :
		rl_a74_t8 = RG_rl_166 ;
	7'h46 :
		rl_a74_t8 = RG_rl_166 ;
	7'h47 :
		rl_a74_t8 = RG_rl_166 ;
	7'h48 :
		rl_a74_t8 = RG_rl_166 ;
	7'h49 :
		rl_a74_t8 = RG_rl_166 ;
	7'h4a :
		rl_a74_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h4b :
		rl_a74_t8 = RG_rl_166 ;
	7'h4c :
		rl_a74_t8 = RG_rl_166 ;
	7'h4d :
		rl_a74_t8 = RG_rl_166 ;
	7'h4e :
		rl_a74_t8 = RG_rl_166 ;
	7'h4f :
		rl_a74_t8 = RG_rl_166 ;
	7'h50 :
		rl_a74_t8 = RG_rl_166 ;
	7'h51 :
		rl_a74_t8 = RG_rl_166 ;
	7'h52 :
		rl_a74_t8 = RG_rl_166 ;
	7'h53 :
		rl_a74_t8 = RG_rl_166 ;
	7'h54 :
		rl_a74_t8 = RG_rl_166 ;
	7'h55 :
		rl_a74_t8 = RG_rl_166 ;
	7'h56 :
		rl_a74_t8 = RG_rl_166 ;
	7'h57 :
		rl_a74_t8 = RG_rl_166 ;
	7'h58 :
		rl_a74_t8 = RG_rl_166 ;
	7'h59 :
		rl_a74_t8 = RG_rl_166 ;
	7'h5a :
		rl_a74_t8 = RG_rl_166 ;
	7'h5b :
		rl_a74_t8 = RG_rl_166 ;
	7'h5c :
		rl_a74_t8 = RG_rl_166 ;
	7'h5d :
		rl_a74_t8 = RG_rl_166 ;
	7'h5e :
		rl_a74_t8 = RG_rl_166 ;
	7'h5f :
		rl_a74_t8 = RG_rl_166 ;
	7'h60 :
		rl_a74_t8 = RG_rl_166 ;
	7'h61 :
		rl_a74_t8 = RG_rl_166 ;
	7'h62 :
		rl_a74_t8 = RG_rl_166 ;
	7'h63 :
		rl_a74_t8 = RG_rl_166 ;
	7'h64 :
		rl_a74_t8 = RG_rl_166 ;
	7'h65 :
		rl_a74_t8 = RG_rl_166 ;
	7'h66 :
		rl_a74_t8 = RG_rl_166 ;
	7'h67 :
		rl_a74_t8 = RG_rl_166 ;
	7'h68 :
		rl_a74_t8 = RG_rl_166 ;
	7'h69 :
		rl_a74_t8 = RG_rl_166 ;
	7'h6a :
		rl_a74_t8 = RG_rl_166 ;
	7'h6b :
		rl_a74_t8 = RG_rl_166 ;
	7'h6c :
		rl_a74_t8 = RG_rl_166 ;
	7'h6d :
		rl_a74_t8 = RG_rl_166 ;
	7'h6e :
		rl_a74_t8 = RG_rl_166 ;
	7'h6f :
		rl_a74_t8 = RG_rl_166 ;
	7'h70 :
		rl_a74_t8 = RG_rl_166 ;
	7'h71 :
		rl_a74_t8 = RG_rl_166 ;
	7'h72 :
		rl_a74_t8 = RG_rl_166 ;
	7'h73 :
		rl_a74_t8 = RG_rl_166 ;
	7'h74 :
		rl_a74_t8 = RG_rl_166 ;
	7'h75 :
		rl_a74_t8 = RG_rl_166 ;
	7'h76 :
		rl_a74_t8 = RG_rl_166 ;
	7'h77 :
		rl_a74_t8 = RG_rl_166 ;
	7'h78 :
		rl_a74_t8 = RG_rl_166 ;
	7'h79 :
		rl_a74_t8 = RG_rl_166 ;
	7'h7a :
		rl_a74_t8 = RG_rl_166 ;
	7'h7b :
		rl_a74_t8 = RG_rl_166 ;
	7'h7c :
		rl_a74_t8 = RG_rl_166 ;
	7'h7d :
		rl_a74_t8 = RG_rl_166 ;
	7'h7e :
		rl_a74_t8 = RG_rl_166 ;
	7'h7f :
		rl_a74_t8 = RG_rl_166 ;
	default :
		rl_a74_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_35 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h01 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h02 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h03 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h04 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h05 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h06 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h07 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h08 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h09 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h0a :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h0b :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h0c :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h0d :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h0e :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h0f :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h10 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h11 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h12 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h13 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h14 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h15 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h16 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h17 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h18 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h19 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h1a :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h1b :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h1c :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h1d :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h1e :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h1f :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h20 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h21 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h22 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h23 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h24 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h25 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h26 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h27 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h28 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h29 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h2a :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h2b :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h2c :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h2d :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h2e :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h2f :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h30 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h31 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h32 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h33 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h34 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h35 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h36 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h37 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h38 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h39 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h3a :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h3b :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h3c :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h3d :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h3e :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h3f :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h40 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h41 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h42 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h43 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h44 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h45 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h46 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h47 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h48 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h49 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h4a :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h4b :
		rl_a75_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h4c :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h4d :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h4e :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h4f :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h50 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h51 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h52 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h53 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h54 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h55 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h56 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h57 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h58 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h59 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h5a :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h5b :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h5c :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h5d :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h5e :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h5f :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h60 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h61 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h62 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h63 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h64 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h65 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h66 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h67 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h68 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h69 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h6a :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h6b :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h6c :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h6d :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h6e :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h6f :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h70 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h71 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h72 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h73 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h74 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h75 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h76 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h77 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h78 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h79 :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h7a :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h7b :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h7c :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h7d :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h7e :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	7'h7f :
		rl_a75_t8 = RG_quantized_block_rl_35 ;
	default :
		rl_a75_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_167 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a76_t8 = RG_rl_167 ;
	7'h01 :
		rl_a76_t8 = RG_rl_167 ;
	7'h02 :
		rl_a76_t8 = RG_rl_167 ;
	7'h03 :
		rl_a76_t8 = RG_rl_167 ;
	7'h04 :
		rl_a76_t8 = RG_rl_167 ;
	7'h05 :
		rl_a76_t8 = RG_rl_167 ;
	7'h06 :
		rl_a76_t8 = RG_rl_167 ;
	7'h07 :
		rl_a76_t8 = RG_rl_167 ;
	7'h08 :
		rl_a76_t8 = RG_rl_167 ;
	7'h09 :
		rl_a76_t8 = RG_rl_167 ;
	7'h0a :
		rl_a76_t8 = RG_rl_167 ;
	7'h0b :
		rl_a76_t8 = RG_rl_167 ;
	7'h0c :
		rl_a76_t8 = RG_rl_167 ;
	7'h0d :
		rl_a76_t8 = RG_rl_167 ;
	7'h0e :
		rl_a76_t8 = RG_rl_167 ;
	7'h0f :
		rl_a76_t8 = RG_rl_167 ;
	7'h10 :
		rl_a76_t8 = RG_rl_167 ;
	7'h11 :
		rl_a76_t8 = RG_rl_167 ;
	7'h12 :
		rl_a76_t8 = RG_rl_167 ;
	7'h13 :
		rl_a76_t8 = RG_rl_167 ;
	7'h14 :
		rl_a76_t8 = RG_rl_167 ;
	7'h15 :
		rl_a76_t8 = RG_rl_167 ;
	7'h16 :
		rl_a76_t8 = RG_rl_167 ;
	7'h17 :
		rl_a76_t8 = RG_rl_167 ;
	7'h18 :
		rl_a76_t8 = RG_rl_167 ;
	7'h19 :
		rl_a76_t8 = RG_rl_167 ;
	7'h1a :
		rl_a76_t8 = RG_rl_167 ;
	7'h1b :
		rl_a76_t8 = RG_rl_167 ;
	7'h1c :
		rl_a76_t8 = RG_rl_167 ;
	7'h1d :
		rl_a76_t8 = RG_rl_167 ;
	7'h1e :
		rl_a76_t8 = RG_rl_167 ;
	7'h1f :
		rl_a76_t8 = RG_rl_167 ;
	7'h20 :
		rl_a76_t8 = RG_rl_167 ;
	7'h21 :
		rl_a76_t8 = RG_rl_167 ;
	7'h22 :
		rl_a76_t8 = RG_rl_167 ;
	7'h23 :
		rl_a76_t8 = RG_rl_167 ;
	7'h24 :
		rl_a76_t8 = RG_rl_167 ;
	7'h25 :
		rl_a76_t8 = RG_rl_167 ;
	7'h26 :
		rl_a76_t8 = RG_rl_167 ;
	7'h27 :
		rl_a76_t8 = RG_rl_167 ;
	7'h28 :
		rl_a76_t8 = RG_rl_167 ;
	7'h29 :
		rl_a76_t8 = RG_rl_167 ;
	7'h2a :
		rl_a76_t8 = RG_rl_167 ;
	7'h2b :
		rl_a76_t8 = RG_rl_167 ;
	7'h2c :
		rl_a76_t8 = RG_rl_167 ;
	7'h2d :
		rl_a76_t8 = RG_rl_167 ;
	7'h2e :
		rl_a76_t8 = RG_rl_167 ;
	7'h2f :
		rl_a76_t8 = RG_rl_167 ;
	7'h30 :
		rl_a76_t8 = RG_rl_167 ;
	7'h31 :
		rl_a76_t8 = RG_rl_167 ;
	7'h32 :
		rl_a76_t8 = RG_rl_167 ;
	7'h33 :
		rl_a76_t8 = RG_rl_167 ;
	7'h34 :
		rl_a76_t8 = RG_rl_167 ;
	7'h35 :
		rl_a76_t8 = RG_rl_167 ;
	7'h36 :
		rl_a76_t8 = RG_rl_167 ;
	7'h37 :
		rl_a76_t8 = RG_rl_167 ;
	7'h38 :
		rl_a76_t8 = RG_rl_167 ;
	7'h39 :
		rl_a76_t8 = RG_rl_167 ;
	7'h3a :
		rl_a76_t8 = RG_rl_167 ;
	7'h3b :
		rl_a76_t8 = RG_rl_167 ;
	7'h3c :
		rl_a76_t8 = RG_rl_167 ;
	7'h3d :
		rl_a76_t8 = RG_rl_167 ;
	7'h3e :
		rl_a76_t8 = RG_rl_167 ;
	7'h3f :
		rl_a76_t8 = RG_rl_167 ;
	7'h40 :
		rl_a76_t8 = RG_rl_167 ;
	7'h41 :
		rl_a76_t8 = RG_rl_167 ;
	7'h42 :
		rl_a76_t8 = RG_rl_167 ;
	7'h43 :
		rl_a76_t8 = RG_rl_167 ;
	7'h44 :
		rl_a76_t8 = RG_rl_167 ;
	7'h45 :
		rl_a76_t8 = RG_rl_167 ;
	7'h46 :
		rl_a76_t8 = RG_rl_167 ;
	7'h47 :
		rl_a76_t8 = RG_rl_167 ;
	7'h48 :
		rl_a76_t8 = RG_rl_167 ;
	7'h49 :
		rl_a76_t8 = RG_rl_167 ;
	7'h4a :
		rl_a76_t8 = RG_rl_167 ;
	7'h4b :
		rl_a76_t8 = RG_rl_167 ;
	7'h4c :
		rl_a76_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h4d :
		rl_a76_t8 = RG_rl_167 ;
	7'h4e :
		rl_a76_t8 = RG_rl_167 ;
	7'h4f :
		rl_a76_t8 = RG_rl_167 ;
	7'h50 :
		rl_a76_t8 = RG_rl_167 ;
	7'h51 :
		rl_a76_t8 = RG_rl_167 ;
	7'h52 :
		rl_a76_t8 = RG_rl_167 ;
	7'h53 :
		rl_a76_t8 = RG_rl_167 ;
	7'h54 :
		rl_a76_t8 = RG_rl_167 ;
	7'h55 :
		rl_a76_t8 = RG_rl_167 ;
	7'h56 :
		rl_a76_t8 = RG_rl_167 ;
	7'h57 :
		rl_a76_t8 = RG_rl_167 ;
	7'h58 :
		rl_a76_t8 = RG_rl_167 ;
	7'h59 :
		rl_a76_t8 = RG_rl_167 ;
	7'h5a :
		rl_a76_t8 = RG_rl_167 ;
	7'h5b :
		rl_a76_t8 = RG_rl_167 ;
	7'h5c :
		rl_a76_t8 = RG_rl_167 ;
	7'h5d :
		rl_a76_t8 = RG_rl_167 ;
	7'h5e :
		rl_a76_t8 = RG_rl_167 ;
	7'h5f :
		rl_a76_t8 = RG_rl_167 ;
	7'h60 :
		rl_a76_t8 = RG_rl_167 ;
	7'h61 :
		rl_a76_t8 = RG_rl_167 ;
	7'h62 :
		rl_a76_t8 = RG_rl_167 ;
	7'h63 :
		rl_a76_t8 = RG_rl_167 ;
	7'h64 :
		rl_a76_t8 = RG_rl_167 ;
	7'h65 :
		rl_a76_t8 = RG_rl_167 ;
	7'h66 :
		rl_a76_t8 = RG_rl_167 ;
	7'h67 :
		rl_a76_t8 = RG_rl_167 ;
	7'h68 :
		rl_a76_t8 = RG_rl_167 ;
	7'h69 :
		rl_a76_t8 = RG_rl_167 ;
	7'h6a :
		rl_a76_t8 = RG_rl_167 ;
	7'h6b :
		rl_a76_t8 = RG_rl_167 ;
	7'h6c :
		rl_a76_t8 = RG_rl_167 ;
	7'h6d :
		rl_a76_t8 = RG_rl_167 ;
	7'h6e :
		rl_a76_t8 = RG_rl_167 ;
	7'h6f :
		rl_a76_t8 = RG_rl_167 ;
	7'h70 :
		rl_a76_t8 = RG_rl_167 ;
	7'h71 :
		rl_a76_t8 = RG_rl_167 ;
	7'h72 :
		rl_a76_t8 = RG_rl_167 ;
	7'h73 :
		rl_a76_t8 = RG_rl_167 ;
	7'h74 :
		rl_a76_t8 = RG_rl_167 ;
	7'h75 :
		rl_a76_t8 = RG_rl_167 ;
	7'h76 :
		rl_a76_t8 = RG_rl_167 ;
	7'h77 :
		rl_a76_t8 = RG_rl_167 ;
	7'h78 :
		rl_a76_t8 = RG_rl_167 ;
	7'h79 :
		rl_a76_t8 = RG_rl_167 ;
	7'h7a :
		rl_a76_t8 = RG_rl_167 ;
	7'h7b :
		rl_a76_t8 = RG_rl_167 ;
	7'h7c :
		rl_a76_t8 = RG_rl_167 ;
	7'h7d :
		rl_a76_t8 = RG_rl_167 ;
	7'h7e :
		rl_a76_t8 = RG_rl_167 ;
	7'h7f :
		rl_a76_t8 = RG_rl_167 ;
	default :
		rl_a76_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_36 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h01 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h02 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h03 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h04 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h05 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h06 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h07 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h08 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h09 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h0a :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h0b :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h0c :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h0d :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h0e :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h0f :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h10 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h11 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h12 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h13 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h14 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h15 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h16 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h17 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h18 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h19 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h1a :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h1b :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h1c :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h1d :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h1e :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h1f :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h20 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h21 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h22 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h23 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h24 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h25 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h26 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h27 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h28 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h29 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h2a :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h2b :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h2c :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h2d :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h2e :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h2f :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h30 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h31 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h32 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h33 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h34 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h35 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h36 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h37 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h38 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h39 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h3a :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h3b :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h3c :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h3d :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h3e :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h3f :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h40 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h41 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h42 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h43 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h44 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h45 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h46 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h47 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h48 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h49 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h4a :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h4b :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h4c :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h4d :
		rl_a77_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h4e :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h4f :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h50 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h51 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h52 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h53 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h54 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h55 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h56 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h57 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h58 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h59 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h5a :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h5b :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h5c :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h5d :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h5e :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h5f :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h60 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h61 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h62 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h63 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h64 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h65 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h66 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h67 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h68 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h69 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h6a :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h6b :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h6c :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h6d :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h6e :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h6f :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h70 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h71 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h72 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h73 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h74 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h75 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h76 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h77 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h78 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h79 :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h7a :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h7b :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h7c :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h7d :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h7e :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	7'h7f :
		rl_a77_t8 = RG_quantized_block_rl_36 ;
	default :
		rl_a77_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_168 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a78_t8 = RG_rl_168 ;
	7'h01 :
		rl_a78_t8 = RG_rl_168 ;
	7'h02 :
		rl_a78_t8 = RG_rl_168 ;
	7'h03 :
		rl_a78_t8 = RG_rl_168 ;
	7'h04 :
		rl_a78_t8 = RG_rl_168 ;
	7'h05 :
		rl_a78_t8 = RG_rl_168 ;
	7'h06 :
		rl_a78_t8 = RG_rl_168 ;
	7'h07 :
		rl_a78_t8 = RG_rl_168 ;
	7'h08 :
		rl_a78_t8 = RG_rl_168 ;
	7'h09 :
		rl_a78_t8 = RG_rl_168 ;
	7'h0a :
		rl_a78_t8 = RG_rl_168 ;
	7'h0b :
		rl_a78_t8 = RG_rl_168 ;
	7'h0c :
		rl_a78_t8 = RG_rl_168 ;
	7'h0d :
		rl_a78_t8 = RG_rl_168 ;
	7'h0e :
		rl_a78_t8 = RG_rl_168 ;
	7'h0f :
		rl_a78_t8 = RG_rl_168 ;
	7'h10 :
		rl_a78_t8 = RG_rl_168 ;
	7'h11 :
		rl_a78_t8 = RG_rl_168 ;
	7'h12 :
		rl_a78_t8 = RG_rl_168 ;
	7'h13 :
		rl_a78_t8 = RG_rl_168 ;
	7'h14 :
		rl_a78_t8 = RG_rl_168 ;
	7'h15 :
		rl_a78_t8 = RG_rl_168 ;
	7'h16 :
		rl_a78_t8 = RG_rl_168 ;
	7'h17 :
		rl_a78_t8 = RG_rl_168 ;
	7'h18 :
		rl_a78_t8 = RG_rl_168 ;
	7'h19 :
		rl_a78_t8 = RG_rl_168 ;
	7'h1a :
		rl_a78_t8 = RG_rl_168 ;
	7'h1b :
		rl_a78_t8 = RG_rl_168 ;
	7'h1c :
		rl_a78_t8 = RG_rl_168 ;
	7'h1d :
		rl_a78_t8 = RG_rl_168 ;
	7'h1e :
		rl_a78_t8 = RG_rl_168 ;
	7'h1f :
		rl_a78_t8 = RG_rl_168 ;
	7'h20 :
		rl_a78_t8 = RG_rl_168 ;
	7'h21 :
		rl_a78_t8 = RG_rl_168 ;
	7'h22 :
		rl_a78_t8 = RG_rl_168 ;
	7'h23 :
		rl_a78_t8 = RG_rl_168 ;
	7'h24 :
		rl_a78_t8 = RG_rl_168 ;
	7'h25 :
		rl_a78_t8 = RG_rl_168 ;
	7'h26 :
		rl_a78_t8 = RG_rl_168 ;
	7'h27 :
		rl_a78_t8 = RG_rl_168 ;
	7'h28 :
		rl_a78_t8 = RG_rl_168 ;
	7'h29 :
		rl_a78_t8 = RG_rl_168 ;
	7'h2a :
		rl_a78_t8 = RG_rl_168 ;
	7'h2b :
		rl_a78_t8 = RG_rl_168 ;
	7'h2c :
		rl_a78_t8 = RG_rl_168 ;
	7'h2d :
		rl_a78_t8 = RG_rl_168 ;
	7'h2e :
		rl_a78_t8 = RG_rl_168 ;
	7'h2f :
		rl_a78_t8 = RG_rl_168 ;
	7'h30 :
		rl_a78_t8 = RG_rl_168 ;
	7'h31 :
		rl_a78_t8 = RG_rl_168 ;
	7'h32 :
		rl_a78_t8 = RG_rl_168 ;
	7'h33 :
		rl_a78_t8 = RG_rl_168 ;
	7'h34 :
		rl_a78_t8 = RG_rl_168 ;
	7'h35 :
		rl_a78_t8 = RG_rl_168 ;
	7'h36 :
		rl_a78_t8 = RG_rl_168 ;
	7'h37 :
		rl_a78_t8 = RG_rl_168 ;
	7'h38 :
		rl_a78_t8 = RG_rl_168 ;
	7'h39 :
		rl_a78_t8 = RG_rl_168 ;
	7'h3a :
		rl_a78_t8 = RG_rl_168 ;
	7'h3b :
		rl_a78_t8 = RG_rl_168 ;
	7'h3c :
		rl_a78_t8 = RG_rl_168 ;
	7'h3d :
		rl_a78_t8 = RG_rl_168 ;
	7'h3e :
		rl_a78_t8 = RG_rl_168 ;
	7'h3f :
		rl_a78_t8 = RG_rl_168 ;
	7'h40 :
		rl_a78_t8 = RG_rl_168 ;
	7'h41 :
		rl_a78_t8 = RG_rl_168 ;
	7'h42 :
		rl_a78_t8 = RG_rl_168 ;
	7'h43 :
		rl_a78_t8 = RG_rl_168 ;
	7'h44 :
		rl_a78_t8 = RG_rl_168 ;
	7'h45 :
		rl_a78_t8 = RG_rl_168 ;
	7'h46 :
		rl_a78_t8 = RG_rl_168 ;
	7'h47 :
		rl_a78_t8 = RG_rl_168 ;
	7'h48 :
		rl_a78_t8 = RG_rl_168 ;
	7'h49 :
		rl_a78_t8 = RG_rl_168 ;
	7'h4a :
		rl_a78_t8 = RG_rl_168 ;
	7'h4b :
		rl_a78_t8 = RG_rl_168 ;
	7'h4c :
		rl_a78_t8 = RG_rl_168 ;
	7'h4d :
		rl_a78_t8 = RG_rl_168 ;
	7'h4e :
		rl_a78_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h4f :
		rl_a78_t8 = RG_rl_168 ;
	7'h50 :
		rl_a78_t8 = RG_rl_168 ;
	7'h51 :
		rl_a78_t8 = RG_rl_168 ;
	7'h52 :
		rl_a78_t8 = RG_rl_168 ;
	7'h53 :
		rl_a78_t8 = RG_rl_168 ;
	7'h54 :
		rl_a78_t8 = RG_rl_168 ;
	7'h55 :
		rl_a78_t8 = RG_rl_168 ;
	7'h56 :
		rl_a78_t8 = RG_rl_168 ;
	7'h57 :
		rl_a78_t8 = RG_rl_168 ;
	7'h58 :
		rl_a78_t8 = RG_rl_168 ;
	7'h59 :
		rl_a78_t8 = RG_rl_168 ;
	7'h5a :
		rl_a78_t8 = RG_rl_168 ;
	7'h5b :
		rl_a78_t8 = RG_rl_168 ;
	7'h5c :
		rl_a78_t8 = RG_rl_168 ;
	7'h5d :
		rl_a78_t8 = RG_rl_168 ;
	7'h5e :
		rl_a78_t8 = RG_rl_168 ;
	7'h5f :
		rl_a78_t8 = RG_rl_168 ;
	7'h60 :
		rl_a78_t8 = RG_rl_168 ;
	7'h61 :
		rl_a78_t8 = RG_rl_168 ;
	7'h62 :
		rl_a78_t8 = RG_rl_168 ;
	7'h63 :
		rl_a78_t8 = RG_rl_168 ;
	7'h64 :
		rl_a78_t8 = RG_rl_168 ;
	7'h65 :
		rl_a78_t8 = RG_rl_168 ;
	7'h66 :
		rl_a78_t8 = RG_rl_168 ;
	7'h67 :
		rl_a78_t8 = RG_rl_168 ;
	7'h68 :
		rl_a78_t8 = RG_rl_168 ;
	7'h69 :
		rl_a78_t8 = RG_rl_168 ;
	7'h6a :
		rl_a78_t8 = RG_rl_168 ;
	7'h6b :
		rl_a78_t8 = RG_rl_168 ;
	7'h6c :
		rl_a78_t8 = RG_rl_168 ;
	7'h6d :
		rl_a78_t8 = RG_rl_168 ;
	7'h6e :
		rl_a78_t8 = RG_rl_168 ;
	7'h6f :
		rl_a78_t8 = RG_rl_168 ;
	7'h70 :
		rl_a78_t8 = RG_rl_168 ;
	7'h71 :
		rl_a78_t8 = RG_rl_168 ;
	7'h72 :
		rl_a78_t8 = RG_rl_168 ;
	7'h73 :
		rl_a78_t8 = RG_rl_168 ;
	7'h74 :
		rl_a78_t8 = RG_rl_168 ;
	7'h75 :
		rl_a78_t8 = RG_rl_168 ;
	7'h76 :
		rl_a78_t8 = RG_rl_168 ;
	7'h77 :
		rl_a78_t8 = RG_rl_168 ;
	7'h78 :
		rl_a78_t8 = RG_rl_168 ;
	7'h79 :
		rl_a78_t8 = RG_rl_168 ;
	7'h7a :
		rl_a78_t8 = RG_rl_168 ;
	7'h7b :
		rl_a78_t8 = RG_rl_168 ;
	7'h7c :
		rl_a78_t8 = RG_rl_168 ;
	7'h7d :
		rl_a78_t8 = RG_rl_168 ;
	7'h7e :
		rl_a78_t8 = RG_rl_168 ;
	7'h7f :
		rl_a78_t8 = RG_rl_168 ;
	default :
		rl_a78_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_37 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h01 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h02 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h03 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h04 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h05 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h06 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h07 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h08 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h09 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h0a :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h0b :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h0c :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h0d :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h0e :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h0f :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h10 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h11 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h12 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h13 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h14 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h15 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h16 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h17 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h18 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h19 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h1a :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h1b :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h1c :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h1d :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h1e :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h1f :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h20 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h21 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h22 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h23 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h24 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h25 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h26 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h27 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h28 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h29 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h2a :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h2b :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h2c :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h2d :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h2e :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h2f :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h30 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h31 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h32 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h33 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h34 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h35 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h36 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h37 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h38 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h39 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h3a :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h3b :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h3c :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h3d :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h3e :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h3f :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h40 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h41 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h42 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h43 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h44 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h45 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h46 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h47 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h48 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h49 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h4a :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h4b :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h4c :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h4d :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h4e :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h4f :
		rl_a79_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h50 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h51 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h52 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h53 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h54 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h55 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h56 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h57 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h58 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h59 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h5a :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h5b :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h5c :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h5d :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h5e :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h5f :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h60 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h61 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h62 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h63 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h64 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h65 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h66 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h67 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h68 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h69 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h6a :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h6b :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h6c :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h6d :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h6e :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h6f :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h70 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h71 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h72 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h73 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h74 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h75 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h76 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h77 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h78 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h79 :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h7a :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h7b :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h7c :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h7d :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h7e :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	7'h7f :
		rl_a79_t8 = RG_quantized_block_rl_37 ;
	default :
		rl_a79_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_169 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a80_t8 = RG_rl_169 ;
	7'h01 :
		rl_a80_t8 = RG_rl_169 ;
	7'h02 :
		rl_a80_t8 = RG_rl_169 ;
	7'h03 :
		rl_a80_t8 = RG_rl_169 ;
	7'h04 :
		rl_a80_t8 = RG_rl_169 ;
	7'h05 :
		rl_a80_t8 = RG_rl_169 ;
	7'h06 :
		rl_a80_t8 = RG_rl_169 ;
	7'h07 :
		rl_a80_t8 = RG_rl_169 ;
	7'h08 :
		rl_a80_t8 = RG_rl_169 ;
	7'h09 :
		rl_a80_t8 = RG_rl_169 ;
	7'h0a :
		rl_a80_t8 = RG_rl_169 ;
	7'h0b :
		rl_a80_t8 = RG_rl_169 ;
	7'h0c :
		rl_a80_t8 = RG_rl_169 ;
	7'h0d :
		rl_a80_t8 = RG_rl_169 ;
	7'h0e :
		rl_a80_t8 = RG_rl_169 ;
	7'h0f :
		rl_a80_t8 = RG_rl_169 ;
	7'h10 :
		rl_a80_t8 = RG_rl_169 ;
	7'h11 :
		rl_a80_t8 = RG_rl_169 ;
	7'h12 :
		rl_a80_t8 = RG_rl_169 ;
	7'h13 :
		rl_a80_t8 = RG_rl_169 ;
	7'h14 :
		rl_a80_t8 = RG_rl_169 ;
	7'h15 :
		rl_a80_t8 = RG_rl_169 ;
	7'h16 :
		rl_a80_t8 = RG_rl_169 ;
	7'h17 :
		rl_a80_t8 = RG_rl_169 ;
	7'h18 :
		rl_a80_t8 = RG_rl_169 ;
	7'h19 :
		rl_a80_t8 = RG_rl_169 ;
	7'h1a :
		rl_a80_t8 = RG_rl_169 ;
	7'h1b :
		rl_a80_t8 = RG_rl_169 ;
	7'h1c :
		rl_a80_t8 = RG_rl_169 ;
	7'h1d :
		rl_a80_t8 = RG_rl_169 ;
	7'h1e :
		rl_a80_t8 = RG_rl_169 ;
	7'h1f :
		rl_a80_t8 = RG_rl_169 ;
	7'h20 :
		rl_a80_t8 = RG_rl_169 ;
	7'h21 :
		rl_a80_t8 = RG_rl_169 ;
	7'h22 :
		rl_a80_t8 = RG_rl_169 ;
	7'h23 :
		rl_a80_t8 = RG_rl_169 ;
	7'h24 :
		rl_a80_t8 = RG_rl_169 ;
	7'h25 :
		rl_a80_t8 = RG_rl_169 ;
	7'h26 :
		rl_a80_t8 = RG_rl_169 ;
	7'h27 :
		rl_a80_t8 = RG_rl_169 ;
	7'h28 :
		rl_a80_t8 = RG_rl_169 ;
	7'h29 :
		rl_a80_t8 = RG_rl_169 ;
	7'h2a :
		rl_a80_t8 = RG_rl_169 ;
	7'h2b :
		rl_a80_t8 = RG_rl_169 ;
	7'h2c :
		rl_a80_t8 = RG_rl_169 ;
	7'h2d :
		rl_a80_t8 = RG_rl_169 ;
	7'h2e :
		rl_a80_t8 = RG_rl_169 ;
	7'h2f :
		rl_a80_t8 = RG_rl_169 ;
	7'h30 :
		rl_a80_t8 = RG_rl_169 ;
	7'h31 :
		rl_a80_t8 = RG_rl_169 ;
	7'h32 :
		rl_a80_t8 = RG_rl_169 ;
	7'h33 :
		rl_a80_t8 = RG_rl_169 ;
	7'h34 :
		rl_a80_t8 = RG_rl_169 ;
	7'h35 :
		rl_a80_t8 = RG_rl_169 ;
	7'h36 :
		rl_a80_t8 = RG_rl_169 ;
	7'h37 :
		rl_a80_t8 = RG_rl_169 ;
	7'h38 :
		rl_a80_t8 = RG_rl_169 ;
	7'h39 :
		rl_a80_t8 = RG_rl_169 ;
	7'h3a :
		rl_a80_t8 = RG_rl_169 ;
	7'h3b :
		rl_a80_t8 = RG_rl_169 ;
	7'h3c :
		rl_a80_t8 = RG_rl_169 ;
	7'h3d :
		rl_a80_t8 = RG_rl_169 ;
	7'h3e :
		rl_a80_t8 = RG_rl_169 ;
	7'h3f :
		rl_a80_t8 = RG_rl_169 ;
	7'h40 :
		rl_a80_t8 = RG_rl_169 ;
	7'h41 :
		rl_a80_t8 = RG_rl_169 ;
	7'h42 :
		rl_a80_t8 = RG_rl_169 ;
	7'h43 :
		rl_a80_t8 = RG_rl_169 ;
	7'h44 :
		rl_a80_t8 = RG_rl_169 ;
	7'h45 :
		rl_a80_t8 = RG_rl_169 ;
	7'h46 :
		rl_a80_t8 = RG_rl_169 ;
	7'h47 :
		rl_a80_t8 = RG_rl_169 ;
	7'h48 :
		rl_a80_t8 = RG_rl_169 ;
	7'h49 :
		rl_a80_t8 = RG_rl_169 ;
	7'h4a :
		rl_a80_t8 = RG_rl_169 ;
	7'h4b :
		rl_a80_t8 = RG_rl_169 ;
	7'h4c :
		rl_a80_t8 = RG_rl_169 ;
	7'h4d :
		rl_a80_t8 = RG_rl_169 ;
	7'h4e :
		rl_a80_t8 = RG_rl_169 ;
	7'h4f :
		rl_a80_t8 = RG_rl_169 ;
	7'h50 :
		rl_a80_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h51 :
		rl_a80_t8 = RG_rl_169 ;
	7'h52 :
		rl_a80_t8 = RG_rl_169 ;
	7'h53 :
		rl_a80_t8 = RG_rl_169 ;
	7'h54 :
		rl_a80_t8 = RG_rl_169 ;
	7'h55 :
		rl_a80_t8 = RG_rl_169 ;
	7'h56 :
		rl_a80_t8 = RG_rl_169 ;
	7'h57 :
		rl_a80_t8 = RG_rl_169 ;
	7'h58 :
		rl_a80_t8 = RG_rl_169 ;
	7'h59 :
		rl_a80_t8 = RG_rl_169 ;
	7'h5a :
		rl_a80_t8 = RG_rl_169 ;
	7'h5b :
		rl_a80_t8 = RG_rl_169 ;
	7'h5c :
		rl_a80_t8 = RG_rl_169 ;
	7'h5d :
		rl_a80_t8 = RG_rl_169 ;
	7'h5e :
		rl_a80_t8 = RG_rl_169 ;
	7'h5f :
		rl_a80_t8 = RG_rl_169 ;
	7'h60 :
		rl_a80_t8 = RG_rl_169 ;
	7'h61 :
		rl_a80_t8 = RG_rl_169 ;
	7'h62 :
		rl_a80_t8 = RG_rl_169 ;
	7'h63 :
		rl_a80_t8 = RG_rl_169 ;
	7'h64 :
		rl_a80_t8 = RG_rl_169 ;
	7'h65 :
		rl_a80_t8 = RG_rl_169 ;
	7'h66 :
		rl_a80_t8 = RG_rl_169 ;
	7'h67 :
		rl_a80_t8 = RG_rl_169 ;
	7'h68 :
		rl_a80_t8 = RG_rl_169 ;
	7'h69 :
		rl_a80_t8 = RG_rl_169 ;
	7'h6a :
		rl_a80_t8 = RG_rl_169 ;
	7'h6b :
		rl_a80_t8 = RG_rl_169 ;
	7'h6c :
		rl_a80_t8 = RG_rl_169 ;
	7'h6d :
		rl_a80_t8 = RG_rl_169 ;
	7'h6e :
		rl_a80_t8 = RG_rl_169 ;
	7'h6f :
		rl_a80_t8 = RG_rl_169 ;
	7'h70 :
		rl_a80_t8 = RG_rl_169 ;
	7'h71 :
		rl_a80_t8 = RG_rl_169 ;
	7'h72 :
		rl_a80_t8 = RG_rl_169 ;
	7'h73 :
		rl_a80_t8 = RG_rl_169 ;
	7'h74 :
		rl_a80_t8 = RG_rl_169 ;
	7'h75 :
		rl_a80_t8 = RG_rl_169 ;
	7'h76 :
		rl_a80_t8 = RG_rl_169 ;
	7'h77 :
		rl_a80_t8 = RG_rl_169 ;
	7'h78 :
		rl_a80_t8 = RG_rl_169 ;
	7'h79 :
		rl_a80_t8 = RG_rl_169 ;
	7'h7a :
		rl_a80_t8 = RG_rl_169 ;
	7'h7b :
		rl_a80_t8 = RG_rl_169 ;
	7'h7c :
		rl_a80_t8 = RG_rl_169 ;
	7'h7d :
		rl_a80_t8 = RG_rl_169 ;
	7'h7e :
		rl_a80_t8 = RG_rl_169 ;
	7'h7f :
		rl_a80_t8 = RG_rl_169 ;
	default :
		rl_a80_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_38 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h01 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h02 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h03 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h04 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h05 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h06 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h07 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h08 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h09 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h0a :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h0b :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h0c :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h0d :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h0e :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h0f :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h10 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h11 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h12 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h13 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h14 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h15 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h16 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h17 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h18 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h19 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h1a :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h1b :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h1c :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h1d :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h1e :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h1f :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h20 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h21 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h22 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h23 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h24 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h25 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h26 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h27 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h28 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h29 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h2a :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h2b :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h2c :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h2d :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h2e :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h2f :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h30 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h31 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h32 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h33 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h34 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h35 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h36 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h37 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h38 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h39 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h3a :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h3b :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h3c :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h3d :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h3e :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h3f :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h40 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h41 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h42 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h43 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h44 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h45 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h46 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h47 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h48 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h49 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h4a :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h4b :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h4c :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h4d :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h4e :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h4f :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h50 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h51 :
		rl_a81_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h52 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h53 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h54 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h55 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h56 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h57 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h58 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h59 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h5a :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h5b :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h5c :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h5d :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h5e :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h5f :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h60 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h61 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h62 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h63 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h64 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h65 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h66 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h67 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h68 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h69 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h6a :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h6b :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h6c :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h6d :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h6e :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h6f :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h70 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h71 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h72 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h73 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h74 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h75 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h76 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h77 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h78 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h79 :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h7a :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h7b :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h7c :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h7d :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h7e :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	7'h7f :
		rl_a81_t8 = RG_quantized_block_rl_38 ;
	default :
		rl_a81_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_170 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a82_t8 = RG_rl_170 ;
	7'h01 :
		rl_a82_t8 = RG_rl_170 ;
	7'h02 :
		rl_a82_t8 = RG_rl_170 ;
	7'h03 :
		rl_a82_t8 = RG_rl_170 ;
	7'h04 :
		rl_a82_t8 = RG_rl_170 ;
	7'h05 :
		rl_a82_t8 = RG_rl_170 ;
	7'h06 :
		rl_a82_t8 = RG_rl_170 ;
	7'h07 :
		rl_a82_t8 = RG_rl_170 ;
	7'h08 :
		rl_a82_t8 = RG_rl_170 ;
	7'h09 :
		rl_a82_t8 = RG_rl_170 ;
	7'h0a :
		rl_a82_t8 = RG_rl_170 ;
	7'h0b :
		rl_a82_t8 = RG_rl_170 ;
	7'h0c :
		rl_a82_t8 = RG_rl_170 ;
	7'h0d :
		rl_a82_t8 = RG_rl_170 ;
	7'h0e :
		rl_a82_t8 = RG_rl_170 ;
	7'h0f :
		rl_a82_t8 = RG_rl_170 ;
	7'h10 :
		rl_a82_t8 = RG_rl_170 ;
	7'h11 :
		rl_a82_t8 = RG_rl_170 ;
	7'h12 :
		rl_a82_t8 = RG_rl_170 ;
	7'h13 :
		rl_a82_t8 = RG_rl_170 ;
	7'h14 :
		rl_a82_t8 = RG_rl_170 ;
	7'h15 :
		rl_a82_t8 = RG_rl_170 ;
	7'h16 :
		rl_a82_t8 = RG_rl_170 ;
	7'h17 :
		rl_a82_t8 = RG_rl_170 ;
	7'h18 :
		rl_a82_t8 = RG_rl_170 ;
	7'h19 :
		rl_a82_t8 = RG_rl_170 ;
	7'h1a :
		rl_a82_t8 = RG_rl_170 ;
	7'h1b :
		rl_a82_t8 = RG_rl_170 ;
	7'h1c :
		rl_a82_t8 = RG_rl_170 ;
	7'h1d :
		rl_a82_t8 = RG_rl_170 ;
	7'h1e :
		rl_a82_t8 = RG_rl_170 ;
	7'h1f :
		rl_a82_t8 = RG_rl_170 ;
	7'h20 :
		rl_a82_t8 = RG_rl_170 ;
	7'h21 :
		rl_a82_t8 = RG_rl_170 ;
	7'h22 :
		rl_a82_t8 = RG_rl_170 ;
	7'h23 :
		rl_a82_t8 = RG_rl_170 ;
	7'h24 :
		rl_a82_t8 = RG_rl_170 ;
	7'h25 :
		rl_a82_t8 = RG_rl_170 ;
	7'h26 :
		rl_a82_t8 = RG_rl_170 ;
	7'h27 :
		rl_a82_t8 = RG_rl_170 ;
	7'h28 :
		rl_a82_t8 = RG_rl_170 ;
	7'h29 :
		rl_a82_t8 = RG_rl_170 ;
	7'h2a :
		rl_a82_t8 = RG_rl_170 ;
	7'h2b :
		rl_a82_t8 = RG_rl_170 ;
	7'h2c :
		rl_a82_t8 = RG_rl_170 ;
	7'h2d :
		rl_a82_t8 = RG_rl_170 ;
	7'h2e :
		rl_a82_t8 = RG_rl_170 ;
	7'h2f :
		rl_a82_t8 = RG_rl_170 ;
	7'h30 :
		rl_a82_t8 = RG_rl_170 ;
	7'h31 :
		rl_a82_t8 = RG_rl_170 ;
	7'h32 :
		rl_a82_t8 = RG_rl_170 ;
	7'h33 :
		rl_a82_t8 = RG_rl_170 ;
	7'h34 :
		rl_a82_t8 = RG_rl_170 ;
	7'h35 :
		rl_a82_t8 = RG_rl_170 ;
	7'h36 :
		rl_a82_t8 = RG_rl_170 ;
	7'h37 :
		rl_a82_t8 = RG_rl_170 ;
	7'h38 :
		rl_a82_t8 = RG_rl_170 ;
	7'h39 :
		rl_a82_t8 = RG_rl_170 ;
	7'h3a :
		rl_a82_t8 = RG_rl_170 ;
	7'h3b :
		rl_a82_t8 = RG_rl_170 ;
	7'h3c :
		rl_a82_t8 = RG_rl_170 ;
	7'h3d :
		rl_a82_t8 = RG_rl_170 ;
	7'h3e :
		rl_a82_t8 = RG_rl_170 ;
	7'h3f :
		rl_a82_t8 = RG_rl_170 ;
	7'h40 :
		rl_a82_t8 = RG_rl_170 ;
	7'h41 :
		rl_a82_t8 = RG_rl_170 ;
	7'h42 :
		rl_a82_t8 = RG_rl_170 ;
	7'h43 :
		rl_a82_t8 = RG_rl_170 ;
	7'h44 :
		rl_a82_t8 = RG_rl_170 ;
	7'h45 :
		rl_a82_t8 = RG_rl_170 ;
	7'h46 :
		rl_a82_t8 = RG_rl_170 ;
	7'h47 :
		rl_a82_t8 = RG_rl_170 ;
	7'h48 :
		rl_a82_t8 = RG_rl_170 ;
	7'h49 :
		rl_a82_t8 = RG_rl_170 ;
	7'h4a :
		rl_a82_t8 = RG_rl_170 ;
	7'h4b :
		rl_a82_t8 = RG_rl_170 ;
	7'h4c :
		rl_a82_t8 = RG_rl_170 ;
	7'h4d :
		rl_a82_t8 = RG_rl_170 ;
	7'h4e :
		rl_a82_t8 = RG_rl_170 ;
	7'h4f :
		rl_a82_t8 = RG_rl_170 ;
	7'h50 :
		rl_a82_t8 = RG_rl_170 ;
	7'h51 :
		rl_a82_t8 = RG_rl_170 ;
	7'h52 :
		rl_a82_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h53 :
		rl_a82_t8 = RG_rl_170 ;
	7'h54 :
		rl_a82_t8 = RG_rl_170 ;
	7'h55 :
		rl_a82_t8 = RG_rl_170 ;
	7'h56 :
		rl_a82_t8 = RG_rl_170 ;
	7'h57 :
		rl_a82_t8 = RG_rl_170 ;
	7'h58 :
		rl_a82_t8 = RG_rl_170 ;
	7'h59 :
		rl_a82_t8 = RG_rl_170 ;
	7'h5a :
		rl_a82_t8 = RG_rl_170 ;
	7'h5b :
		rl_a82_t8 = RG_rl_170 ;
	7'h5c :
		rl_a82_t8 = RG_rl_170 ;
	7'h5d :
		rl_a82_t8 = RG_rl_170 ;
	7'h5e :
		rl_a82_t8 = RG_rl_170 ;
	7'h5f :
		rl_a82_t8 = RG_rl_170 ;
	7'h60 :
		rl_a82_t8 = RG_rl_170 ;
	7'h61 :
		rl_a82_t8 = RG_rl_170 ;
	7'h62 :
		rl_a82_t8 = RG_rl_170 ;
	7'h63 :
		rl_a82_t8 = RG_rl_170 ;
	7'h64 :
		rl_a82_t8 = RG_rl_170 ;
	7'h65 :
		rl_a82_t8 = RG_rl_170 ;
	7'h66 :
		rl_a82_t8 = RG_rl_170 ;
	7'h67 :
		rl_a82_t8 = RG_rl_170 ;
	7'h68 :
		rl_a82_t8 = RG_rl_170 ;
	7'h69 :
		rl_a82_t8 = RG_rl_170 ;
	7'h6a :
		rl_a82_t8 = RG_rl_170 ;
	7'h6b :
		rl_a82_t8 = RG_rl_170 ;
	7'h6c :
		rl_a82_t8 = RG_rl_170 ;
	7'h6d :
		rl_a82_t8 = RG_rl_170 ;
	7'h6e :
		rl_a82_t8 = RG_rl_170 ;
	7'h6f :
		rl_a82_t8 = RG_rl_170 ;
	7'h70 :
		rl_a82_t8 = RG_rl_170 ;
	7'h71 :
		rl_a82_t8 = RG_rl_170 ;
	7'h72 :
		rl_a82_t8 = RG_rl_170 ;
	7'h73 :
		rl_a82_t8 = RG_rl_170 ;
	7'h74 :
		rl_a82_t8 = RG_rl_170 ;
	7'h75 :
		rl_a82_t8 = RG_rl_170 ;
	7'h76 :
		rl_a82_t8 = RG_rl_170 ;
	7'h77 :
		rl_a82_t8 = RG_rl_170 ;
	7'h78 :
		rl_a82_t8 = RG_rl_170 ;
	7'h79 :
		rl_a82_t8 = RG_rl_170 ;
	7'h7a :
		rl_a82_t8 = RG_rl_170 ;
	7'h7b :
		rl_a82_t8 = RG_rl_170 ;
	7'h7c :
		rl_a82_t8 = RG_rl_170 ;
	7'h7d :
		rl_a82_t8 = RG_rl_170 ;
	7'h7e :
		rl_a82_t8 = RG_rl_170 ;
	7'h7f :
		rl_a82_t8 = RG_rl_170 ;
	default :
		rl_a82_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_39 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h01 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h02 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h03 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h04 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h05 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h06 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h07 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h08 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h09 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h0a :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h0b :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h0c :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h0d :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h0e :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h0f :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h10 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h11 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h12 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h13 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h14 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h15 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h16 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h17 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h18 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h19 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h1a :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h1b :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h1c :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h1d :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h1e :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h1f :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h20 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h21 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h22 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h23 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h24 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h25 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h26 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h27 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h28 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h29 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h2a :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h2b :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h2c :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h2d :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h2e :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h2f :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h30 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h31 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h32 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h33 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h34 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h35 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h36 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h37 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h38 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h39 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h3a :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h3b :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h3c :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h3d :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h3e :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h3f :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h40 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h41 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h42 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h43 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h44 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h45 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h46 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h47 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h48 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h49 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h4a :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h4b :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h4c :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h4d :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h4e :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h4f :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h50 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h51 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h52 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h53 :
		rl_a83_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h54 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h55 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h56 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h57 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h58 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h59 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h5a :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h5b :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h5c :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h5d :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h5e :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h5f :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h60 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h61 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h62 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h63 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h64 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h65 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h66 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h67 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h68 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h69 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h6a :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h6b :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h6c :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h6d :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h6e :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h6f :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h70 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h71 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h72 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h73 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h74 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h75 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h76 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h77 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h78 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h79 :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h7a :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h7b :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h7c :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h7d :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h7e :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	7'h7f :
		rl_a83_t8 = RG_quantized_block_rl_39 ;
	default :
		rl_a83_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_171 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a84_t8 = RG_rl_171 ;
	7'h01 :
		rl_a84_t8 = RG_rl_171 ;
	7'h02 :
		rl_a84_t8 = RG_rl_171 ;
	7'h03 :
		rl_a84_t8 = RG_rl_171 ;
	7'h04 :
		rl_a84_t8 = RG_rl_171 ;
	7'h05 :
		rl_a84_t8 = RG_rl_171 ;
	7'h06 :
		rl_a84_t8 = RG_rl_171 ;
	7'h07 :
		rl_a84_t8 = RG_rl_171 ;
	7'h08 :
		rl_a84_t8 = RG_rl_171 ;
	7'h09 :
		rl_a84_t8 = RG_rl_171 ;
	7'h0a :
		rl_a84_t8 = RG_rl_171 ;
	7'h0b :
		rl_a84_t8 = RG_rl_171 ;
	7'h0c :
		rl_a84_t8 = RG_rl_171 ;
	7'h0d :
		rl_a84_t8 = RG_rl_171 ;
	7'h0e :
		rl_a84_t8 = RG_rl_171 ;
	7'h0f :
		rl_a84_t8 = RG_rl_171 ;
	7'h10 :
		rl_a84_t8 = RG_rl_171 ;
	7'h11 :
		rl_a84_t8 = RG_rl_171 ;
	7'h12 :
		rl_a84_t8 = RG_rl_171 ;
	7'h13 :
		rl_a84_t8 = RG_rl_171 ;
	7'h14 :
		rl_a84_t8 = RG_rl_171 ;
	7'h15 :
		rl_a84_t8 = RG_rl_171 ;
	7'h16 :
		rl_a84_t8 = RG_rl_171 ;
	7'h17 :
		rl_a84_t8 = RG_rl_171 ;
	7'h18 :
		rl_a84_t8 = RG_rl_171 ;
	7'h19 :
		rl_a84_t8 = RG_rl_171 ;
	7'h1a :
		rl_a84_t8 = RG_rl_171 ;
	7'h1b :
		rl_a84_t8 = RG_rl_171 ;
	7'h1c :
		rl_a84_t8 = RG_rl_171 ;
	7'h1d :
		rl_a84_t8 = RG_rl_171 ;
	7'h1e :
		rl_a84_t8 = RG_rl_171 ;
	7'h1f :
		rl_a84_t8 = RG_rl_171 ;
	7'h20 :
		rl_a84_t8 = RG_rl_171 ;
	7'h21 :
		rl_a84_t8 = RG_rl_171 ;
	7'h22 :
		rl_a84_t8 = RG_rl_171 ;
	7'h23 :
		rl_a84_t8 = RG_rl_171 ;
	7'h24 :
		rl_a84_t8 = RG_rl_171 ;
	7'h25 :
		rl_a84_t8 = RG_rl_171 ;
	7'h26 :
		rl_a84_t8 = RG_rl_171 ;
	7'h27 :
		rl_a84_t8 = RG_rl_171 ;
	7'h28 :
		rl_a84_t8 = RG_rl_171 ;
	7'h29 :
		rl_a84_t8 = RG_rl_171 ;
	7'h2a :
		rl_a84_t8 = RG_rl_171 ;
	7'h2b :
		rl_a84_t8 = RG_rl_171 ;
	7'h2c :
		rl_a84_t8 = RG_rl_171 ;
	7'h2d :
		rl_a84_t8 = RG_rl_171 ;
	7'h2e :
		rl_a84_t8 = RG_rl_171 ;
	7'h2f :
		rl_a84_t8 = RG_rl_171 ;
	7'h30 :
		rl_a84_t8 = RG_rl_171 ;
	7'h31 :
		rl_a84_t8 = RG_rl_171 ;
	7'h32 :
		rl_a84_t8 = RG_rl_171 ;
	7'h33 :
		rl_a84_t8 = RG_rl_171 ;
	7'h34 :
		rl_a84_t8 = RG_rl_171 ;
	7'h35 :
		rl_a84_t8 = RG_rl_171 ;
	7'h36 :
		rl_a84_t8 = RG_rl_171 ;
	7'h37 :
		rl_a84_t8 = RG_rl_171 ;
	7'h38 :
		rl_a84_t8 = RG_rl_171 ;
	7'h39 :
		rl_a84_t8 = RG_rl_171 ;
	7'h3a :
		rl_a84_t8 = RG_rl_171 ;
	7'h3b :
		rl_a84_t8 = RG_rl_171 ;
	7'h3c :
		rl_a84_t8 = RG_rl_171 ;
	7'h3d :
		rl_a84_t8 = RG_rl_171 ;
	7'h3e :
		rl_a84_t8 = RG_rl_171 ;
	7'h3f :
		rl_a84_t8 = RG_rl_171 ;
	7'h40 :
		rl_a84_t8 = RG_rl_171 ;
	7'h41 :
		rl_a84_t8 = RG_rl_171 ;
	7'h42 :
		rl_a84_t8 = RG_rl_171 ;
	7'h43 :
		rl_a84_t8 = RG_rl_171 ;
	7'h44 :
		rl_a84_t8 = RG_rl_171 ;
	7'h45 :
		rl_a84_t8 = RG_rl_171 ;
	7'h46 :
		rl_a84_t8 = RG_rl_171 ;
	7'h47 :
		rl_a84_t8 = RG_rl_171 ;
	7'h48 :
		rl_a84_t8 = RG_rl_171 ;
	7'h49 :
		rl_a84_t8 = RG_rl_171 ;
	7'h4a :
		rl_a84_t8 = RG_rl_171 ;
	7'h4b :
		rl_a84_t8 = RG_rl_171 ;
	7'h4c :
		rl_a84_t8 = RG_rl_171 ;
	7'h4d :
		rl_a84_t8 = RG_rl_171 ;
	7'h4e :
		rl_a84_t8 = RG_rl_171 ;
	7'h4f :
		rl_a84_t8 = RG_rl_171 ;
	7'h50 :
		rl_a84_t8 = RG_rl_171 ;
	7'h51 :
		rl_a84_t8 = RG_rl_171 ;
	7'h52 :
		rl_a84_t8 = RG_rl_171 ;
	7'h53 :
		rl_a84_t8 = RG_rl_171 ;
	7'h54 :
		rl_a84_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h55 :
		rl_a84_t8 = RG_rl_171 ;
	7'h56 :
		rl_a84_t8 = RG_rl_171 ;
	7'h57 :
		rl_a84_t8 = RG_rl_171 ;
	7'h58 :
		rl_a84_t8 = RG_rl_171 ;
	7'h59 :
		rl_a84_t8 = RG_rl_171 ;
	7'h5a :
		rl_a84_t8 = RG_rl_171 ;
	7'h5b :
		rl_a84_t8 = RG_rl_171 ;
	7'h5c :
		rl_a84_t8 = RG_rl_171 ;
	7'h5d :
		rl_a84_t8 = RG_rl_171 ;
	7'h5e :
		rl_a84_t8 = RG_rl_171 ;
	7'h5f :
		rl_a84_t8 = RG_rl_171 ;
	7'h60 :
		rl_a84_t8 = RG_rl_171 ;
	7'h61 :
		rl_a84_t8 = RG_rl_171 ;
	7'h62 :
		rl_a84_t8 = RG_rl_171 ;
	7'h63 :
		rl_a84_t8 = RG_rl_171 ;
	7'h64 :
		rl_a84_t8 = RG_rl_171 ;
	7'h65 :
		rl_a84_t8 = RG_rl_171 ;
	7'h66 :
		rl_a84_t8 = RG_rl_171 ;
	7'h67 :
		rl_a84_t8 = RG_rl_171 ;
	7'h68 :
		rl_a84_t8 = RG_rl_171 ;
	7'h69 :
		rl_a84_t8 = RG_rl_171 ;
	7'h6a :
		rl_a84_t8 = RG_rl_171 ;
	7'h6b :
		rl_a84_t8 = RG_rl_171 ;
	7'h6c :
		rl_a84_t8 = RG_rl_171 ;
	7'h6d :
		rl_a84_t8 = RG_rl_171 ;
	7'h6e :
		rl_a84_t8 = RG_rl_171 ;
	7'h6f :
		rl_a84_t8 = RG_rl_171 ;
	7'h70 :
		rl_a84_t8 = RG_rl_171 ;
	7'h71 :
		rl_a84_t8 = RG_rl_171 ;
	7'h72 :
		rl_a84_t8 = RG_rl_171 ;
	7'h73 :
		rl_a84_t8 = RG_rl_171 ;
	7'h74 :
		rl_a84_t8 = RG_rl_171 ;
	7'h75 :
		rl_a84_t8 = RG_rl_171 ;
	7'h76 :
		rl_a84_t8 = RG_rl_171 ;
	7'h77 :
		rl_a84_t8 = RG_rl_171 ;
	7'h78 :
		rl_a84_t8 = RG_rl_171 ;
	7'h79 :
		rl_a84_t8 = RG_rl_171 ;
	7'h7a :
		rl_a84_t8 = RG_rl_171 ;
	7'h7b :
		rl_a84_t8 = RG_rl_171 ;
	7'h7c :
		rl_a84_t8 = RG_rl_171 ;
	7'h7d :
		rl_a84_t8 = RG_rl_171 ;
	7'h7e :
		rl_a84_t8 = RG_rl_171 ;
	7'h7f :
		rl_a84_t8 = RG_rl_171 ;
	default :
		rl_a84_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_40 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h01 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h02 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h03 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h04 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h05 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h06 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h07 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h08 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h09 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h0a :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h0b :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h0c :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h0d :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h0e :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h0f :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h10 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h11 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h12 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h13 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h14 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h15 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h16 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h17 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h18 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h19 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h1a :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h1b :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h1c :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h1d :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h1e :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h1f :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h20 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h21 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h22 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h23 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h24 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h25 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h26 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h27 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h28 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h29 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h2a :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h2b :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h2c :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h2d :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h2e :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h2f :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h30 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h31 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h32 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h33 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h34 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h35 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h36 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h37 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h38 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h39 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h3a :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h3b :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h3c :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h3d :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h3e :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h3f :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h40 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h41 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h42 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h43 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h44 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h45 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h46 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h47 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h48 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h49 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h4a :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h4b :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h4c :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h4d :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h4e :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h4f :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h50 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h51 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h52 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h53 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h54 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h55 :
		rl_a85_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h56 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h57 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h58 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h59 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h5a :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h5b :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h5c :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h5d :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h5e :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h5f :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h60 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h61 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h62 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h63 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h64 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h65 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h66 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h67 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h68 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h69 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h6a :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h6b :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h6c :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h6d :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h6e :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h6f :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h70 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h71 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h72 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h73 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h74 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h75 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h76 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h77 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h78 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h79 :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h7a :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h7b :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h7c :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h7d :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h7e :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	7'h7f :
		rl_a85_t8 = RG_quantized_block_rl_40 ;
	default :
		rl_a85_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_172 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a86_t8 = RG_rl_172 ;
	7'h01 :
		rl_a86_t8 = RG_rl_172 ;
	7'h02 :
		rl_a86_t8 = RG_rl_172 ;
	7'h03 :
		rl_a86_t8 = RG_rl_172 ;
	7'h04 :
		rl_a86_t8 = RG_rl_172 ;
	7'h05 :
		rl_a86_t8 = RG_rl_172 ;
	7'h06 :
		rl_a86_t8 = RG_rl_172 ;
	7'h07 :
		rl_a86_t8 = RG_rl_172 ;
	7'h08 :
		rl_a86_t8 = RG_rl_172 ;
	7'h09 :
		rl_a86_t8 = RG_rl_172 ;
	7'h0a :
		rl_a86_t8 = RG_rl_172 ;
	7'h0b :
		rl_a86_t8 = RG_rl_172 ;
	7'h0c :
		rl_a86_t8 = RG_rl_172 ;
	7'h0d :
		rl_a86_t8 = RG_rl_172 ;
	7'h0e :
		rl_a86_t8 = RG_rl_172 ;
	7'h0f :
		rl_a86_t8 = RG_rl_172 ;
	7'h10 :
		rl_a86_t8 = RG_rl_172 ;
	7'h11 :
		rl_a86_t8 = RG_rl_172 ;
	7'h12 :
		rl_a86_t8 = RG_rl_172 ;
	7'h13 :
		rl_a86_t8 = RG_rl_172 ;
	7'h14 :
		rl_a86_t8 = RG_rl_172 ;
	7'h15 :
		rl_a86_t8 = RG_rl_172 ;
	7'h16 :
		rl_a86_t8 = RG_rl_172 ;
	7'h17 :
		rl_a86_t8 = RG_rl_172 ;
	7'h18 :
		rl_a86_t8 = RG_rl_172 ;
	7'h19 :
		rl_a86_t8 = RG_rl_172 ;
	7'h1a :
		rl_a86_t8 = RG_rl_172 ;
	7'h1b :
		rl_a86_t8 = RG_rl_172 ;
	7'h1c :
		rl_a86_t8 = RG_rl_172 ;
	7'h1d :
		rl_a86_t8 = RG_rl_172 ;
	7'h1e :
		rl_a86_t8 = RG_rl_172 ;
	7'h1f :
		rl_a86_t8 = RG_rl_172 ;
	7'h20 :
		rl_a86_t8 = RG_rl_172 ;
	7'h21 :
		rl_a86_t8 = RG_rl_172 ;
	7'h22 :
		rl_a86_t8 = RG_rl_172 ;
	7'h23 :
		rl_a86_t8 = RG_rl_172 ;
	7'h24 :
		rl_a86_t8 = RG_rl_172 ;
	7'h25 :
		rl_a86_t8 = RG_rl_172 ;
	7'h26 :
		rl_a86_t8 = RG_rl_172 ;
	7'h27 :
		rl_a86_t8 = RG_rl_172 ;
	7'h28 :
		rl_a86_t8 = RG_rl_172 ;
	7'h29 :
		rl_a86_t8 = RG_rl_172 ;
	7'h2a :
		rl_a86_t8 = RG_rl_172 ;
	7'h2b :
		rl_a86_t8 = RG_rl_172 ;
	7'h2c :
		rl_a86_t8 = RG_rl_172 ;
	7'h2d :
		rl_a86_t8 = RG_rl_172 ;
	7'h2e :
		rl_a86_t8 = RG_rl_172 ;
	7'h2f :
		rl_a86_t8 = RG_rl_172 ;
	7'h30 :
		rl_a86_t8 = RG_rl_172 ;
	7'h31 :
		rl_a86_t8 = RG_rl_172 ;
	7'h32 :
		rl_a86_t8 = RG_rl_172 ;
	7'h33 :
		rl_a86_t8 = RG_rl_172 ;
	7'h34 :
		rl_a86_t8 = RG_rl_172 ;
	7'h35 :
		rl_a86_t8 = RG_rl_172 ;
	7'h36 :
		rl_a86_t8 = RG_rl_172 ;
	7'h37 :
		rl_a86_t8 = RG_rl_172 ;
	7'h38 :
		rl_a86_t8 = RG_rl_172 ;
	7'h39 :
		rl_a86_t8 = RG_rl_172 ;
	7'h3a :
		rl_a86_t8 = RG_rl_172 ;
	7'h3b :
		rl_a86_t8 = RG_rl_172 ;
	7'h3c :
		rl_a86_t8 = RG_rl_172 ;
	7'h3d :
		rl_a86_t8 = RG_rl_172 ;
	7'h3e :
		rl_a86_t8 = RG_rl_172 ;
	7'h3f :
		rl_a86_t8 = RG_rl_172 ;
	7'h40 :
		rl_a86_t8 = RG_rl_172 ;
	7'h41 :
		rl_a86_t8 = RG_rl_172 ;
	7'h42 :
		rl_a86_t8 = RG_rl_172 ;
	7'h43 :
		rl_a86_t8 = RG_rl_172 ;
	7'h44 :
		rl_a86_t8 = RG_rl_172 ;
	7'h45 :
		rl_a86_t8 = RG_rl_172 ;
	7'h46 :
		rl_a86_t8 = RG_rl_172 ;
	7'h47 :
		rl_a86_t8 = RG_rl_172 ;
	7'h48 :
		rl_a86_t8 = RG_rl_172 ;
	7'h49 :
		rl_a86_t8 = RG_rl_172 ;
	7'h4a :
		rl_a86_t8 = RG_rl_172 ;
	7'h4b :
		rl_a86_t8 = RG_rl_172 ;
	7'h4c :
		rl_a86_t8 = RG_rl_172 ;
	7'h4d :
		rl_a86_t8 = RG_rl_172 ;
	7'h4e :
		rl_a86_t8 = RG_rl_172 ;
	7'h4f :
		rl_a86_t8 = RG_rl_172 ;
	7'h50 :
		rl_a86_t8 = RG_rl_172 ;
	7'h51 :
		rl_a86_t8 = RG_rl_172 ;
	7'h52 :
		rl_a86_t8 = RG_rl_172 ;
	7'h53 :
		rl_a86_t8 = RG_rl_172 ;
	7'h54 :
		rl_a86_t8 = RG_rl_172 ;
	7'h55 :
		rl_a86_t8 = RG_rl_172 ;
	7'h56 :
		rl_a86_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h57 :
		rl_a86_t8 = RG_rl_172 ;
	7'h58 :
		rl_a86_t8 = RG_rl_172 ;
	7'h59 :
		rl_a86_t8 = RG_rl_172 ;
	7'h5a :
		rl_a86_t8 = RG_rl_172 ;
	7'h5b :
		rl_a86_t8 = RG_rl_172 ;
	7'h5c :
		rl_a86_t8 = RG_rl_172 ;
	7'h5d :
		rl_a86_t8 = RG_rl_172 ;
	7'h5e :
		rl_a86_t8 = RG_rl_172 ;
	7'h5f :
		rl_a86_t8 = RG_rl_172 ;
	7'h60 :
		rl_a86_t8 = RG_rl_172 ;
	7'h61 :
		rl_a86_t8 = RG_rl_172 ;
	7'h62 :
		rl_a86_t8 = RG_rl_172 ;
	7'h63 :
		rl_a86_t8 = RG_rl_172 ;
	7'h64 :
		rl_a86_t8 = RG_rl_172 ;
	7'h65 :
		rl_a86_t8 = RG_rl_172 ;
	7'h66 :
		rl_a86_t8 = RG_rl_172 ;
	7'h67 :
		rl_a86_t8 = RG_rl_172 ;
	7'h68 :
		rl_a86_t8 = RG_rl_172 ;
	7'h69 :
		rl_a86_t8 = RG_rl_172 ;
	7'h6a :
		rl_a86_t8 = RG_rl_172 ;
	7'h6b :
		rl_a86_t8 = RG_rl_172 ;
	7'h6c :
		rl_a86_t8 = RG_rl_172 ;
	7'h6d :
		rl_a86_t8 = RG_rl_172 ;
	7'h6e :
		rl_a86_t8 = RG_rl_172 ;
	7'h6f :
		rl_a86_t8 = RG_rl_172 ;
	7'h70 :
		rl_a86_t8 = RG_rl_172 ;
	7'h71 :
		rl_a86_t8 = RG_rl_172 ;
	7'h72 :
		rl_a86_t8 = RG_rl_172 ;
	7'h73 :
		rl_a86_t8 = RG_rl_172 ;
	7'h74 :
		rl_a86_t8 = RG_rl_172 ;
	7'h75 :
		rl_a86_t8 = RG_rl_172 ;
	7'h76 :
		rl_a86_t8 = RG_rl_172 ;
	7'h77 :
		rl_a86_t8 = RG_rl_172 ;
	7'h78 :
		rl_a86_t8 = RG_rl_172 ;
	7'h79 :
		rl_a86_t8 = RG_rl_172 ;
	7'h7a :
		rl_a86_t8 = RG_rl_172 ;
	7'h7b :
		rl_a86_t8 = RG_rl_172 ;
	7'h7c :
		rl_a86_t8 = RG_rl_172 ;
	7'h7d :
		rl_a86_t8 = RG_rl_172 ;
	7'h7e :
		rl_a86_t8 = RG_rl_172 ;
	7'h7f :
		rl_a86_t8 = RG_rl_172 ;
	default :
		rl_a86_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_41 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h01 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h02 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h03 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h04 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h05 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h06 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h07 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h08 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h09 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h0a :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h0b :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h0c :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h0d :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h0e :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h0f :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h10 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h11 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h12 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h13 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h14 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h15 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h16 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h17 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h18 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h19 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h1a :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h1b :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h1c :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h1d :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h1e :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h1f :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h20 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h21 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h22 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h23 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h24 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h25 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h26 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h27 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h28 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h29 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h2a :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h2b :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h2c :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h2d :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h2e :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h2f :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h30 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h31 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h32 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h33 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h34 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h35 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h36 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h37 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h38 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h39 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h3a :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h3b :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h3c :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h3d :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h3e :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h3f :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h40 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h41 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h42 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h43 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h44 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h45 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h46 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h47 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h48 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h49 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h4a :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h4b :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h4c :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h4d :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h4e :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h4f :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h50 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h51 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h52 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h53 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h54 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h55 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h56 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h57 :
		rl_a87_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h58 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h59 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h5a :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h5b :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h5c :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h5d :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h5e :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h5f :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h60 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h61 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h62 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h63 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h64 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h65 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h66 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h67 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h68 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h69 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h6a :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h6b :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h6c :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h6d :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h6e :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h6f :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h70 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h71 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h72 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h73 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h74 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h75 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h76 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h77 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h78 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h79 :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h7a :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h7b :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h7c :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h7d :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h7e :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	7'h7f :
		rl_a87_t8 = RG_quantized_block_rl_41 ;
	default :
		rl_a87_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_173 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a88_t8 = RG_rl_173 ;
	7'h01 :
		rl_a88_t8 = RG_rl_173 ;
	7'h02 :
		rl_a88_t8 = RG_rl_173 ;
	7'h03 :
		rl_a88_t8 = RG_rl_173 ;
	7'h04 :
		rl_a88_t8 = RG_rl_173 ;
	7'h05 :
		rl_a88_t8 = RG_rl_173 ;
	7'h06 :
		rl_a88_t8 = RG_rl_173 ;
	7'h07 :
		rl_a88_t8 = RG_rl_173 ;
	7'h08 :
		rl_a88_t8 = RG_rl_173 ;
	7'h09 :
		rl_a88_t8 = RG_rl_173 ;
	7'h0a :
		rl_a88_t8 = RG_rl_173 ;
	7'h0b :
		rl_a88_t8 = RG_rl_173 ;
	7'h0c :
		rl_a88_t8 = RG_rl_173 ;
	7'h0d :
		rl_a88_t8 = RG_rl_173 ;
	7'h0e :
		rl_a88_t8 = RG_rl_173 ;
	7'h0f :
		rl_a88_t8 = RG_rl_173 ;
	7'h10 :
		rl_a88_t8 = RG_rl_173 ;
	7'h11 :
		rl_a88_t8 = RG_rl_173 ;
	7'h12 :
		rl_a88_t8 = RG_rl_173 ;
	7'h13 :
		rl_a88_t8 = RG_rl_173 ;
	7'h14 :
		rl_a88_t8 = RG_rl_173 ;
	7'h15 :
		rl_a88_t8 = RG_rl_173 ;
	7'h16 :
		rl_a88_t8 = RG_rl_173 ;
	7'h17 :
		rl_a88_t8 = RG_rl_173 ;
	7'h18 :
		rl_a88_t8 = RG_rl_173 ;
	7'h19 :
		rl_a88_t8 = RG_rl_173 ;
	7'h1a :
		rl_a88_t8 = RG_rl_173 ;
	7'h1b :
		rl_a88_t8 = RG_rl_173 ;
	7'h1c :
		rl_a88_t8 = RG_rl_173 ;
	7'h1d :
		rl_a88_t8 = RG_rl_173 ;
	7'h1e :
		rl_a88_t8 = RG_rl_173 ;
	7'h1f :
		rl_a88_t8 = RG_rl_173 ;
	7'h20 :
		rl_a88_t8 = RG_rl_173 ;
	7'h21 :
		rl_a88_t8 = RG_rl_173 ;
	7'h22 :
		rl_a88_t8 = RG_rl_173 ;
	7'h23 :
		rl_a88_t8 = RG_rl_173 ;
	7'h24 :
		rl_a88_t8 = RG_rl_173 ;
	7'h25 :
		rl_a88_t8 = RG_rl_173 ;
	7'h26 :
		rl_a88_t8 = RG_rl_173 ;
	7'h27 :
		rl_a88_t8 = RG_rl_173 ;
	7'h28 :
		rl_a88_t8 = RG_rl_173 ;
	7'h29 :
		rl_a88_t8 = RG_rl_173 ;
	7'h2a :
		rl_a88_t8 = RG_rl_173 ;
	7'h2b :
		rl_a88_t8 = RG_rl_173 ;
	7'h2c :
		rl_a88_t8 = RG_rl_173 ;
	7'h2d :
		rl_a88_t8 = RG_rl_173 ;
	7'h2e :
		rl_a88_t8 = RG_rl_173 ;
	7'h2f :
		rl_a88_t8 = RG_rl_173 ;
	7'h30 :
		rl_a88_t8 = RG_rl_173 ;
	7'h31 :
		rl_a88_t8 = RG_rl_173 ;
	7'h32 :
		rl_a88_t8 = RG_rl_173 ;
	7'h33 :
		rl_a88_t8 = RG_rl_173 ;
	7'h34 :
		rl_a88_t8 = RG_rl_173 ;
	7'h35 :
		rl_a88_t8 = RG_rl_173 ;
	7'h36 :
		rl_a88_t8 = RG_rl_173 ;
	7'h37 :
		rl_a88_t8 = RG_rl_173 ;
	7'h38 :
		rl_a88_t8 = RG_rl_173 ;
	7'h39 :
		rl_a88_t8 = RG_rl_173 ;
	7'h3a :
		rl_a88_t8 = RG_rl_173 ;
	7'h3b :
		rl_a88_t8 = RG_rl_173 ;
	7'h3c :
		rl_a88_t8 = RG_rl_173 ;
	7'h3d :
		rl_a88_t8 = RG_rl_173 ;
	7'h3e :
		rl_a88_t8 = RG_rl_173 ;
	7'h3f :
		rl_a88_t8 = RG_rl_173 ;
	7'h40 :
		rl_a88_t8 = RG_rl_173 ;
	7'h41 :
		rl_a88_t8 = RG_rl_173 ;
	7'h42 :
		rl_a88_t8 = RG_rl_173 ;
	7'h43 :
		rl_a88_t8 = RG_rl_173 ;
	7'h44 :
		rl_a88_t8 = RG_rl_173 ;
	7'h45 :
		rl_a88_t8 = RG_rl_173 ;
	7'h46 :
		rl_a88_t8 = RG_rl_173 ;
	7'h47 :
		rl_a88_t8 = RG_rl_173 ;
	7'h48 :
		rl_a88_t8 = RG_rl_173 ;
	7'h49 :
		rl_a88_t8 = RG_rl_173 ;
	7'h4a :
		rl_a88_t8 = RG_rl_173 ;
	7'h4b :
		rl_a88_t8 = RG_rl_173 ;
	7'h4c :
		rl_a88_t8 = RG_rl_173 ;
	7'h4d :
		rl_a88_t8 = RG_rl_173 ;
	7'h4e :
		rl_a88_t8 = RG_rl_173 ;
	7'h4f :
		rl_a88_t8 = RG_rl_173 ;
	7'h50 :
		rl_a88_t8 = RG_rl_173 ;
	7'h51 :
		rl_a88_t8 = RG_rl_173 ;
	7'h52 :
		rl_a88_t8 = RG_rl_173 ;
	7'h53 :
		rl_a88_t8 = RG_rl_173 ;
	7'h54 :
		rl_a88_t8 = RG_rl_173 ;
	7'h55 :
		rl_a88_t8 = RG_rl_173 ;
	7'h56 :
		rl_a88_t8 = RG_rl_173 ;
	7'h57 :
		rl_a88_t8 = RG_rl_173 ;
	7'h58 :
		rl_a88_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h59 :
		rl_a88_t8 = RG_rl_173 ;
	7'h5a :
		rl_a88_t8 = RG_rl_173 ;
	7'h5b :
		rl_a88_t8 = RG_rl_173 ;
	7'h5c :
		rl_a88_t8 = RG_rl_173 ;
	7'h5d :
		rl_a88_t8 = RG_rl_173 ;
	7'h5e :
		rl_a88_t8 = RG_rl_173 ;
	7'h5f :
		rl_a88_t8 = RG_rl_173 ;
	7'h60 :
		rl_a88_t8 = RG_rl_173 ;
	7'h61 :
		rl_a88_t8 = RG_rl_173 ;
	7'h62 :
		rl_a88_t8 = RG_rl_173 ;
	7'h63 :
		rl_a88_t8 = RG_rl_173 ;
	7'h64 :
		rl_a88_t8 = RG_rl_173 ;
	7'h65 :
		rl_a88_t8 = RG_rl_173 ;
	7'h66 :
		rl_a88_t8 = RG_rl_173 ;
	7'h67 :
		rl_a88_t8 = RG_rl_173 ;
	7'h68 :
		rl_a88_t8 = RG_rl_173 ;
	7'h69 :
		rl_a88_t8 = RG_rl_173 ;
	7'h6a :
		rl_a88_t8 = RG_rl_173 ;
	7'h6b :
		rl_a88_t8 = RG_rl_173 ;
	7'h6c :
		rl_a88_t8 = RG_rl_173 ;
	7'h6d :
		rl_a88_t8 = RG_rl_173 ;
	7'h6e :
		rl_a88_t8 = RG_rl_173 ;
	7'h6f :
		rl_a88_t8 = RG_rl_173 ;
	7'h70 :
		rl_a88_t8 = RG_rl_173 ;
	7'h71 :
		rl_a88_t8 = RG_rl_173 ;
	7'h72 :
		rl_a88_t8 = RG_rl_173 ;
	7'h73 :
		rl_a88_t8 = RG_rl_173 ;
	7'h74 :
		rl_a88_t8 = RG_rl_173 ;
	7'h75 :
		rl_a88_t8 = RG_rl_173 ;
	7'h76 :
		rl_a88_t8 = RG_rl_173 ;
	7'h77 :
		rl_a88_t8 = RG_rl_173 ;
	7'h78 :
		rl_a88_t8 = RG_rl_173 ;
	7'h79 :
		rl_a88_t8 = RG_rl_173 ;
	7'h7a :
		rl_a88_t8 = RG_rl_173 ;
	7'h7b :
		rl_a88_t8 = RG_rl_173 ;
	7'h7c :
		rl_a88_t8 = RG_rl_173 ;
	7'h7d :
		rl_a88_t8 = RG_rl_173 ;
	7'h7e :
		rl_a88_t8 = RG_rl_173 ;
	7'h7f :
		rl_a88_t8 = RG_rl_173 ;
	default :
		rl_a88_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_42 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h01 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h02 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h03 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h04 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h05 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h06 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h07 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h08 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h09 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h0a :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h0b :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h0c :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h0d :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h0e :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h0f :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h10 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h11 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h12 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h13 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h14 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h15 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h16 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h17 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h18 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h19 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h1a :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h1b :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h1c :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h1d :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h1e :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h1f :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h20 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h21 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h22 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h23 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h24 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h25 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h26 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h27 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h28 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h29 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h2a :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h2b :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h2c :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h2d :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h2e :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h2f :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h30 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h31 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h32 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h33 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h34 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h35 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h36 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h37 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h38 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h39 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h3a :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h3b :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h3c :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h3d :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h3e :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h3f :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h40 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h41 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h42 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h43 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h44 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h45 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h46 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h47 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h48 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h49 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h4a :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h4b :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h4c :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h4d :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h4e :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h4f :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h50 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h51 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h52 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h53 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h54 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h55 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h56 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h57 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h58 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h59 :
		rl_a89_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h5a :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h5b :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h5c :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h5d :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h5e :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h5f :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h60 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h61 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h62 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h63 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h64 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h65 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h66 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h67 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h68 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h69 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h6a :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h6b :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h6c :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h6d :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h6e :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h6f :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h70 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h71 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h72 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h73 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h74 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h75 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h76 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h77 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h78 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h79 :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h7a :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h7b :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h7c :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h7d :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h7e :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	7'h7f :
		rl_a89_t8 = RG_quantized_block_rl_42 ;
	default :
		rl_a89_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_174 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a90_t8 = RG_rl_174 ;
	7'h01 :
		rl_a90_t8 = RG_rl_174 ;
	7'h02 :
		rl_a90_t8 = RG_rl_174 ;
	7'h03 :
		rl_a90_t8 = RG_rl_174 ;
	7'h04 :
		rl_a90_t8 = RG_rl_174 ;
	7'h05 :
		rl_a90_t8 = RG_rl_174 ;
	7'h06 :
		rl_a90_t8 = RG_rl_174 ;
	7'h07 :
		rl_a90_t8 = RG_rl_174 ;
	7'h08 :
		rl_a90_t8 = RG_rl_174 ;
	7'h09 :
		rl_a90_t8 = RG_rl_174 ;
	7'h0a :
		rl_a90_t8 = RG_rl_174 ;
	7'h0b :
		rl_a90_t8 = RG_rl_174 ;
	7'h0c :
		rl_a90_t8 = RG_rl_174 ;
	7'h0d :
		rl_a90_t8 = RG_rl_174 ;
	7'h0e :
		rl_a90_t8 = RG_rl_174 ;
	7'h0f :
		rl_a90_t8 = RG_rl_174 ;
	7'h10 :
		rl_a90_t8 = RG_rl_174 ;
	7'h11 :
		rl_a90_t8 = RG_rl_174 ;
	7'h12 :
		rl_a90_t8 = RG_rl_174 ;
	7'h13 :
		rl_a90_t8 = RG_rl_174 ;
	7'h14 :
		rl_a90_t8 = RG_rl_174 ;
	7'h15 :
		rl_a90_t8 = RG_rl_174 ;
	7'h16 :
		rl_a90_t8 = RG_rl_174 ;
	7'h17 :
		rl_a90_t8 = RG_rl_174 ;
	7'h18 :
		rl_a90_t8 = RG_rl_174 ;
	7'h19 :
		rl_a90_t8 = RG_rl_174 ;
	7'h1a :
		rl_a90_t8 = RG_rl_174 ;
	7'h1b :
		rl_a90_t8 = RG_rl_174 ;
	7'h1c :
		rl_a90_t8 = RG_rl_174 ;
	7'h1d :
		rl_a90_t8 = RG_rl_174 ;
	7'h1e :
		rl_a90_t8 = RG_rl_174 ;
	7'h1f :
		rl_a90_t8 = RG_rl_174 ;
	7'h20 :
		rl_a90_t8 = RG_rl_174 ;
	7'h21 :
		rl_a90_t8 = RG_rl_174 ;
	7'h22 :
		rl_a90_t8 = RG_rl_174 ;
	7'h23 :
		rl_a90_t8 = RG_rl_174 ;
	7'h24 :
		rl_a90_t8 = RG_rl_174 ;
	7'h25 :
		rl_a90_t8 = RG_rl_174 ;
	7'h26 :
		rl_a90_t8 = RG_rl_174 ;
	7'h27 :
		rl_a90_t8 = RG_rl_174 ;
	7'h28 :
		rl_a90_t8 = RG_rl_174 ;
	7'h29 :
		rl_a90_t8 = RG_rl_174 ;
	7'h2a :
		rl_a90_t8 = RG_rl_174 ;
	7'h2b :
		rl_a90_t8 = RG_rl_174 ;
	7'h2c :
		rl_a90_t8 = RG_rl_174 ;
	7'h2d :
		rl_a90_t8 = RG_rl_174 ;
	7'h2e :
		rl_a90_t8 = RG_rl_174 ;
	7'h2f :
		rl_a90_t8 = RG_rl_174 ;
	7'h30 :
		rl_a90_t8 = RG_rl_174 ;
	7'h31 :
		rl_a90_t8 = RG_rl_174 ;
	7'h32 :
		rl_a90_t8 = RG_rl_174 ;
	7'h33 :
		rl_a90_t8 = RG_rl_174 ;
	7'h34 :
		rl_a90_t8 = RG_rl_174 ;
	7'h35 :
		rl_a90_t8 = RG_rl_174 ;
	7'h36 :
		rl_a90_t8 = RG_rl_174 ;
	7'h37 :
		rl_a90_t8 = RG_rl_174 ;
	7'h38 :
		rl_a90_t8 = RG_rl_174 ;
	7'h39 :
		rl_a90_t8 = RG_rl_174 ;
	7'h3a :
		rl_a90_t8 = RG_rl_174 ;
	7'h3b :
		rl_a90_t8 = RG_rl_174 ;
	7'h3c :
		rl_a90_t8 = RG_rl_174 ;
	7'h3d :
		rl_a90_t8 = RG_rl_174 ;
	7'h3e :
		rl_a90_t8 = RG_rl_174 ;
	7'h3f :
		rl_a90_t8 = RG_rl_174 ;
	7'h40 :
		rl_a90_t8 = RG_rl_174 ;
	7'h41 :
		rl_a90_t8 = RG_rl_174 ;
	7'h42 :
		rl_a90_t8 = RG_rl_174 ;
	7'h43 :
		rl_a90_t8 = RG_rl_174 ;
	7'h44 :
		rl_a90_t8 = RG_rl_174 ;
	7'h45 :
		rl_a90_t8 = RG_rl_174 ;
	7'h46 :
		rl_a90_t8 = RG_rl_174 ;
	7'h47 :
		rl_a90_t8 = RG_rl_174 ;
	7'h48 :
		rl_a90_t8 = RG_rl_174 ;
	7'h49 :
		rl_a90_t8 = RG_rl_174 ;
	7'h4a :
		rl_a90_t8 = RG_rl_174 ;
	7'h4b :
		rl_a90_t8 = RG_rl_174 ;
	7'h4c :
		rl_a90_t8 = RG_rl_174 ;
	7'h4d :
		rl_a90_t8 = RG_rl_174 ;
	7'h4e :
		rl_a90_t8 = RG_rl_174 ;
	7'h4f :
		rl_a90_t8 = RG_rl_174 ;
	7'h50 :
		rl_a90_t8 = RG_rl_174 ;
	7'h51 :
		rl_a90_t8 = RG_rl_174 ;
	7'h52 :
		rl_a90_t8 = RG_rl_174 ;
	7'h53 :
		rl_a90_t8 = RG_rl_174 ;
	7'h54 :
		rl_a90_t8 = RG_rl_174 ;
	7'h55 :
		rl_a90_t8 = RG_rl_174 ;
	7'h56 :
		rl_a90_t8 = RG_rl_174 ;
	7'h57 :
		rl_a90_t8 = RG_rl_174 ;
	7'h58 :
		rl_a90_t8 = RG_rl_174 ;
	7'h59 :
		rl_a90_t8 = RG_rl_174 ;
	7'h5a :
		rl_a90_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h5b :
		rl_a90_t8 = RG_rl_174 ;
	7'h5c :
		rl_a90_t8 = RG_rl_174 ;
	7'h5d :
		rl_a90_t8 = RG_rl_174 ;
	7'h5e :
		rl_a90_t8 = RG_rl_174 ;
	7'h5f :
		rl_a90_t8 = RG_rl_174 ;
	7'h60 :
		rl_a90_t8 = RG_rl_174 ;
	7'h61 :
		rl_a90_t8 = RG_rl_174 ;
	7'h62 :
		rl_a90_t8 = RG_rl_174 ;
	7'h63 :
		rl_a90_t8 = RG_rl_174 ;
	7'h64 :
		rl_a90_t8 = RG_rl_174 ;
	7'h65 :
		rl_a90_t8 = RG_rl_174 ;
	7'h66 :
		rl_a90_t8 = RG_rl_174 ;
	7'h67 :
		rl_a90_t8 = RG_rl_174 ;
	7'h68 :
		rl_a90_t8 = RG_rl_174 ;
	7'h69 :
		rl_a90_t8 = RG_rl_174 ;
	7'h6a :
		rl_a90_t8 = RG_rl_174 ;
	7'h6b :
		rl_a90_t8 = RG_rl_174 ;
	7'h6c :
		rl_a90_t8 = RG_rl_174 ;
	7'h6d :
		rl_a90_t8 = RG_rl_174 ;
	7'h6e :
		rl_a90_t8 = RG_rl_174 ;
	7'h6f :
		rl_a90_t8 = RG_rl_174 ;
	7'h70 :
		rl_a90_t8 = RG_rl_174 ;
	7'h71 :
		rl_a90_t8 = RG_rl_174 ;
	7'h72 :
		rl_a90_t8 = RG_rl_174 ;
	7'h73 :
		rl_a90_t8 = RG_rl_174 ;
	7'h74 :
		rl_a90_t8 = RG_rl_174 ;
	7'h75 :
		rl_a90_t8 = RG_rl_174 ;
	7'h76 :
		rl_a90_t8 = RG_rl_174 ;
	7'h77 :
		rl_a90_t8 = RG_rl_174 ;
	7'h78 :
		rl_a90_t8 = RG_rl_174 ;
	7'h79 :
		rl_a90_t8 = RG_rl_174 ;
	7'h7a :
		rl_a90_t8 = RG_rl_174 ;
	7'h7b :
		rl_a90_t8 = RG_rl_174 ;
	7'h7c :
		rl_a90_t8 = RG_rl_174 ;
	7'h7d :
		rl_a90_t8 = RG_rl_174 ;
	7'h7e :
		rl_a90_t8 = RG_rl_174 ;
	7'h7f :
		rl_a90_t8 = RG_rl_174 ;
	default :
		rl_a90_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_43 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h01 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h02 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h03 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h04 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h05 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h06 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h07 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h08 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h09 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h0a :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h0b :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h0c :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h0d :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h0e :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h0f :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h10 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h11 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h12 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h13 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h14 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h15 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h16 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h17 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h18 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h19 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h1a :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h1b :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h1c :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h1d :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h1e :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h1f :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h20 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h21 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h22 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h23 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h24 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h25 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h26 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h27 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h28 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h29 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h2a :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h2b :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h2c :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h2d :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h2e :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h2f :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h30 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h31 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h32 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h33 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h34 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h35 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h36 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h37 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h38 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h39 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h3a :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h3b :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h3c :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h3d :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h3e :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h3f :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h40 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h41 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h42 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h43 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h44 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h45 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h46 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h47 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h48 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h49 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h4a :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h4b :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h4c :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h4d :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h4e :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h4f :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h50 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h51 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h52 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h53 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h54 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h55 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h56 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h57 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h58 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h59 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h5a :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h5b :
		rl_a91_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h5c :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h5d :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h5e :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h5f :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h60 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h61 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h62 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h63 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h64 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h65 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h66 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h67 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h68 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h69 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h6a :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h6b :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h6c :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h6d :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h6e :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h6f :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h70 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h71 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h72 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h73 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h74 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h75 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h76 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h77 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h78 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h79 :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h7a :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h7b :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h7c :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h7d :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h7e :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	7'h7f :
		rl_a91_t8 = RG_quantized_block_rl_43 ;
	default :
		rl_a91_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_175 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a92_t8 = RG_rl_175 ;
	7'h01 :
		rl_a92_t8 = RG_rl_175 ;
	7'h02 :
		rl_a92_t8 = RG_rl_175 ;
	7'h03 :
		rl_a92_t8 = RG_rl_175 ;
	7'h04 :
		rl_a92_t8 = RG_rl_175 ;
	7'h05 :
		rl_a92_t8 = RG_rl_175 ;
	7'h06 :
		rl_a92_t8 = RG_rl_175 ;
	7'h07 :
		rl_a92_t8 = RG_rl_175 ;
	7'h08 :
		rl_a92_t8 = RG_rl_175 ;
	7'h09 :
		rl_a92_t8 = RG_rl_175 ;
	7'h0a :
		rl_a92_t8 = RG_rl_175 ;
	7'h0b :
		rl_a92_t8 = RG_rl_175 ;
	7'h0c :
		rl_a92_t8 = RG_rl_175 ;
	7'h0d :
		rl_a92_t8 = RG_rl_175 ;
	7'h0e :
		rl_a92_t8 = RG_rl_175 ;
	7'h0f :
		rl_a92_t8 = RG_rl_175 ;
	7'h10 :
		rl_a92_t8 = RG_rl_175 ;
	7'h11 :
		rl_a92_t8 = RG_rl_175 ;
	7'h12 :
		rl_a92_t8 = RG_rl_175 ;
	7'h13 :
		rl_a92_t8 = RG_rl_175 ;
	7'h14 :
		rl_a92_t8 = RG_rl_175 ;
	7'h15 :
		rl_a92_t8 = RG_rl_175 ;
	7'h16 :
		rl_a92_t8 = RG_rl_175 ;
	7'h17 :
		rl_a92_t8 = RG_rl_175 ;
	7'h18 :
		rl_a92_t8 = RG_rl_175 ;
	7'h19 :
		rl_a92_t8 = RG_rl_175 ;
	7'h1a :
		rl_a92_t8 = RG_rl_175 ;
	7'h1b :
		rl_a92_t8 = RG_rl_175 ;
	7'h1c :
		rl_a92_t8 = RG_rl_175 ;
	7'h1d :
		rl_a92_t8 = RG_rl_175 ;
	7'h1e :
		rl_a92_t8 = RG_rl_175 ;
	7'h1f :
		rl_a92_t8 = RG_rl_175 ;
	7'h20 :
		rl_a92_t8 = RG_rl_175 ;
	7'h21 :
		rl_a92_t8 = RG_rl_175 ;
	7'h22 :
		rl_a92_t8 = RG_rl_175 ;
	7'h23 :
		rl_a92_t8 = RG_rl_175 ;
	7'h24 :
		rl_a92_t8 = RG_rl_175 ;
	7'h25 :
		rl_a92_t8 = RG_rl_175 ;
	7'h26 :
		rl_a92_t8 = RG_rl_175 ;
	7'h27 :
		rl_a92_t8 = RG_rl_175 ;
	7'h28 :
		rl_a92_t8 = RG_rl_175 ;
	7'h29 :
		rl_a92_t8 = RG_rl_175 ;
	7'h2a :
		rl_a92_t8 = RG_rl_175 ;
	7'h2b :
		rl_a92_t8 = RG_rl_175 ;
	7'h2c :
		rl_a92_t8 = RG_rl_175 ;
	7'h2d :
		rl_a92_t8 = RG_rl_175 ;
	7'h2e :
		rl_a92_t8 = RG_rl_175 ;
	7'h2f :
		rl_a92_t8 = RG_rl_175 ;
	7'h30 :
		rl_a92_t8 = RG_rl_175 ;
	7'h31 :
		rl_a92_t8 = RG_rl_175 ;
	7'h32 :
		rl_a92_t8 = RG_rl_175 ;
	7'h33 :
		rl_a92_t8 = RG_rl_175 ;
	7'h34 :
		rl_a92_t8 = RG_rl_175 ;
	7'h35 :
		rl_a92_t8 = RG_rl_175 ;
	7'h36 :
		rl_a92_t8 = RG_rl_175 ;
	7'h37 :
		rl_a92_t8 = RG_rl_175 ;
	7'h38 :
		rl_a92_t8 = RG_rl_175 ;
	7'h39 :
		rl_a92_t8 = RG_rl_175 ;
	7'h3a :
		rl_a92_t8 = RG_rl_175 ;
	7'h3b :
		rl_a92_t8 = RG_rl_175 ;
	7'h3c :
		rl_a92_t8 = RG_rl_175 ;
	7'h3d :
		rl_a92_t8 = RG_rl_175 ;
	7'h3e :
		rl_a92_t8 = RG_rl_175 ;
	7'h3f :
		rl_a92_t8 = RG_rl_175 ;
	7'h40 :
		rl_a92_t8 = RG_rl_175 ;
	7'h41 :
		rl_a92_t8 = RG_rl_175 ;
	7'h42 :
		rl_a92_t8 = RG_rl_175 ;
	7'h43 :
		rl_a92_t8 = RG_rl_175 ;
	7'h44 :
		rl_a92_t8 = RG_rl_175 ;
	7'h45 :
		rl_a92_t8 = RG_rl_175 ;
	7'h46 :
		rl_a92_t8 = RG_rl_175 ;
	7'h47 :
		rl_a92_t8 = RG_rl_175 ;
	7'h48 :
		rl_a92_t8 = RG_rl_175 ;
	7'h49 :
		rl_a92_t8 = RG_rl_175 ;
	7'h4a :
		rl_a92_t8 = RG_rl_175 ;
	7'h4b :
		rl_a92_t8 = RG_rl_175 ;
	7'h4c :
		rl_a92_t8 = RG_rl_175 ;
	7'h4d :
		rl_a92_t8 = RG_rl_175 ;
	7'h4e :
		rl_a92_t8 = RG_rl_175 ;
	7'h4f :
		rl_a92_t8 = RG_rl_175 ;
	7'h50 :
		rl_a92_t8 = RG_rl_175 ;
	7'h51 :
		rl_a92_t8 = RG_rl_175 ;
	7'h52 :
		rl_a92_t8 = RG_rl_175 ;
	7'h53 :
		rl_a92_t8 = RG_rl_175 ;
	7'h54 :
		rl_a92_t8 = RG_rl_175 ;
	7'h55 :
		rl_a92_t8 = RG_rl_175 ;
	7'h56 :
		rl_a92_t8 = RG_rl_175 ;
	7'h57 :
		rl_a92_t8 = RG_rl_175 ;
	7'h58 :
		rl_a92_t8 = RG_rl_175 ;
	7'h59 :
		rl_a92_t8 = RG_rl_175 ;
	7'h5a :
		rl_a92_t8 = RG_rl_175 ;
	7'h5b :
		rl_a92_t8 = RG_rl_175 ;
	7'h5c :
		rl_a92_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h5d :
		rl_a92_t8 = RG_rl_175 ;
	7'h5e :
		rl_a92_t8 = RG_rl_175 ;
	7'h5f :
		rl_a92_t8 = RG_rl_175 ;
	7'h60 :
		rl_a92_t8 = RG_rl_175 ;
	7'h61 :
		rl_a92_t8 = RG_rl_175 ;
	7'h62 :
		rl_a92_t8 = RG_rl_175 ;
	7'h63 :
		rl_a92_t8 = RG_rl_175 ;
	7'h64 :
		rl_a92_t8 = RG_rl_175 ;
	7'h65 :
		rl_a92_t8 = RG_rl_175 ;
	7'h66 :
		rl_a92_t8 = RG_rl_175 ;
	7'h67 :
		rl_a92_t8 = RG_rl_175 ;
	7'h68 :
		rl_a92_t8 = RG_rl_175 ;
	7'h69 :
		rl_a92_t8 = RG_rl_175 ;
	7'h6a :
		rl_a92_t8 = RG_rl_175 ;
	7'h6b :
		rl_a92_t8 = RG_rl_175 ;
	7'h6c :
		rl_a92_t8 = RG_rl_175 ;
	7'h6d :
		rl_a92_t8 = RG_rl_175 ;
	7'h6e :
		rl_a92_t8 = RG_rl_175 ;
	7'h6f :
		rl_a92_t8 = RG_rl_175 ;
	7'h70 :
		rl_a92_t8 = RG_rl_175 ;
	7'h71 :
		rl_a92_t8 = RG_rl_175 ;
	7'h72 :
		rl_a92_t8 = RG_rl_175 ;
	7'h73 :
		rl_a92_t8 = RG_rl_175 ;
	7'h74 :
		rl_a92_t8 = RG_rl_175 ;
	7'h75 :
		rl_a92_t8 = RG_rl_175 ;
	7'h76 :
		rl_a92_t8 = RG_rl_175 ;
	7'h77 :
		rl_a92_t8 = RG_rl_175 ;
	7'h78 :
		rl_a92_t8 = RG_rl_175 ;
	7'h79 :
		rl_a92_t8 = RG_rl_175 ;
	7'h7a :
		rl_a92_t8 = RG_rl_175 ;
	7'h7b :
		rl_a92_t8 = RG_rl_175 ;
	7'h7c :
		rl_a92_t8 = RG_rl_175 ;
	7'h7d :
		rl_a92_t8 = RG_rl_175 ;
	7'h7e :
		rl_a92_t8 = RG_rl_175 ;
	7'h7f :
		rl_a92_t8 = RG_rl_175 ;
	default :
		rl_a92_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_44 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h01 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h02 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h03 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h04 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h05 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h06 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h07 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h08 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h09 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h0a :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h0b :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h0c :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h0d :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h0e :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h0f :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h10 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h11 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h12 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h13 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h14 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h15 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h16 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h17 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h18 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h19 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h1a :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h1b :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h1c :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h1d :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h1e :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h1f :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h20 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h21 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h22 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h23 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h24 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h25 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h26 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h27 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h28 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h29 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h2a :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h2b :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h2c :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h2d :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h2e :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h2f :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h30 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h31 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h32 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h33 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h34 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h35 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h36 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h37 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h38 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h39 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h3a :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h3b :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h3c :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h3d :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h3e :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h3f :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h40 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h41 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h42 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h43 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h44 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h45 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h46 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h47 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h48 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h49 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h4a :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h4b :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h4c :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h4d :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h4e :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h4f :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h50 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h51 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h52 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h53 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h54 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h55 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h56 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h57 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h58 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h59 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h5a :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h5b :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h5c :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h5d :
		rl_a93_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h5e :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h5f :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h60 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h61 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h62 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h63 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h64 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h65 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h66 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h67 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h68 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h69 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h6a :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h6b :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h6c :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h6d :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h6e :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h6f :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h70 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h71 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h72 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h73 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h74 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h75 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h76 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h77 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h78 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h79 :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h7a :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h7b :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h7c :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h7d :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h7e :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	7'h7f :
		rl_a93_t8 = RG_quantized_block_rl_44 ;
	default :
		rl_a93_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_176 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a94_t8 = RG_rl_176 ;
	7'h01 :
		rl_a94_t8 = RG_rl_176 ;
	7'h02 :
		rl_a94_t8 = RG_rl_176 ;
	7'h03 :
		rl_a94_t8 = RG_rl_176 ;
	7'h04 :
		rl_a94_t8 = RG_rl_176 ;
	7'h05 :
		rl_a94_t8 = RG_rl_176 ;
	7'h06 :
		rl_a94_t8 = RG_rl_176 ;
	7'h07 :
		rl_a94_t8 = RG_rl_176 ;
	7'h08 :
		rl_a94_t8 = RG_rl_176 ;
	7'h09 :
		rl_a94_t8 = RG_rl_176 ;
	7'h0a :
		rl_a94_t8 = RG_rl_176 ;
	7'h0b :
		rl_a94_t8 = RG_rl_176 ;
	7'h0c :
		rl_a94_t8 = RG_rl_176 ;
	7'h0d :
		rl_a94_t8 = RG_rl_176 ;
	7'h0e :
		rl_a94_t8 = RG_rl_176 ;
	7'h0f :
		rl_a94_t8 = RG_rl_176 ;
	7'h10 :
		rl_a94_t8 = RG_rl_176 ;
	7'h11 :
		rl_a94_t8 = RG_rl_176 ;
	7'h12 :
		rl_a94_t8 = RG_rl_176 ;
	7'h13 :
		rl_a94_t8 = RG_rl_176 ;
	7'h14 :
		rl_a94_t8 = RG_rl_176 ;
	7'h15 :
		rl_a94_t8 = RG_rl_176 ;
	7'h16 :
		rl_a94_t8 = RG_rl_176 ;
	7'h17 :
		rl_a94_t8 = RG_rl_176 ;
	7'h18 :
		rl_a94_t8 = RG_rl_176 ;
	7'h19 :
		rl_a94_t8 = RG_rl_176 ;
	7'h1a :
		rl_a94_t8 = RG_rl_176 ;
	7'h1b :
		rl_a94_t8 = RG_rl_176 ;
	7'h1c :
		rl_a94_t8 = RG_rl_176 ;
	7'h1d :
		rl_a94_t8 = RG_rl_176 ;
	7'h1e :
		rl_a94_t8 = RG_rl_176 ;
	7'h1f :
		rl_a94_t8 = RG_rl_176 ;
	7'h20 :
		rl_a94_t8 = RG_rl_176 ;
	7'h21 :
		rl_a94_t8 = RG_rl_176 ;
	7'h22 :
		rl_a94_t8 = RG_rl_176 ;
	7'h23 :
		rl_a94_t8 = RG_rl_176 ;
	7'h24 :
		rl_a94_t8 = RG_rl_176 ;
	7'h25 :
		rl_a94_t8 = RG_rl_176 ;
	7'h26 :
		rl_a94_t8 = RG_rl_176 ;
	7'h27 :
		rl_a94_t8 = RG_rl_176 ;
	7'h28 :
		rl_a94_t8 = RG_rl_176 ;
	7'h29 :
		rl_a94_t8 = RG_rl_176 ;
	7'h2a :
		rl_a94_t8 = RG_rl_176 ;
	7'h2b :
		rl_a94_t8 = RG_rl_176 ;
	7'h2c :
		rl_a94_t8 = RG_rl_176 ;
	7'h2d :
		rl_a94_t8 = RG_rl_176 ;
	7'h2e :
		rl_a94_t8 = RG_rl_176 ;
	7'h2f :
		rl_a94_t8 = RG_rl_176 ;
	7'h30 :
		rl_a94_t8 = RG_rl_176 ;
	7'h31 :
		rl_a94_t8 = RG_rl_176 ;
	7'h32 :
		rl_a94_t8 = RG_rl_176 ;
	7'h33 :
		rl_a94_t8 = RG_rl_176 ;
	7'h34 :
		rl_a94_t8 = RG_rl_176 ;
	7'h35 :
		rl_a94_t8 = RG_rl_176 ;
	7'h36 :
		rl_a94_t8 = RG_rl_176 ;
	7'h37 :
		rl_a94_t8 = RG_rl_176 ;
	7'h38 :
		rl_a94_t8 = RG_rl_176 ;
	7'h39 :
		rl_a94_t8 = RG_rl_176 ;
	7'h3a :
		rl_a94_t8 = RG_rl_176 ;
	7'h3b :
		rl_a94_t8 = RG_rl_176 ;
	7'h3c :
		rl_a94_t8 = RG_rl_176 ;
	7'h3d :
		rl_a94_t8 = RG_rl_176 ;
	7'h3e :
		rl_a94_t8 = RG_rl_176 ;
	7'h3f :
		rl_a94_t8 = RG_rl_176 ;
	7'h40 :
		rl_a94_t8 = RG_rl_176 ;
	7'h41 :
		rl_a94_t8 = RG_rl_176 ;
	7'h42 :
		rl_a94_t8 = RG_rl_176 ;
	7'h43 :
		rl_a94_t8 = RG_rl_176 ;
	7'h44 :
		rl_a94_t8 = RG_rl_176 ;
	7'h45 :
		rl_a94_t8 = RG_rl_176 ;
	7'h46 :
		rl_a94_t8 = RG_rl_176 ;
	7'h47 :
		rl_a94_t8 = RG_rl_176 ;
	7'h48 :
		rl_a94_t8 = RG_rl_176 ;
	7'h49 :
		rl_a94_t8 = RG_rl_176 ;
	7'h4a :
		rl_a94_t8 = RG_rl_176 ;
	7'h4b :
		rl_a94_t8 = RG_rl_176 ;
	7'h4c :
		rl_a94_t8 = RG_rl_176 ;
	7'h4d :
		rl_a94_t8 = RG_rl_176 ;
	7'h4e :
		rl_a94_t8 = RG_rl_176 ;
	7'h4f :
		rl_a94_t8 = RG_rl_176 ;
	7'h50 :
		rl_a94_t8 = RG_rl_176 ;
	7'h51 :
		rl_a94_t8 = RG_rl_176 ;
	7'h52 :
		rl_a94_t8 = RG_rl_176 ;
	7'h53 :
		rl_a94_t8 = RG_rl_176 ;
	7'h54 :
		rl_a94_t8 = RG_rl_176 ;
	7'h55 :
		rl_a94_t8 = RG_rl_176 ;
	7'h56 :
		rl_a94_t8 = RG_rl_176 ;
	7'h57 :
		rl_a94_t8 = RG_rl_176 ;
	7'h58 :
		rl_a94_t8 = RG_rl_176 ;
	7'h59 :
		rl_a94_t8 = RG_rl_176 ;
	7'h5a :
		rl_a94_t8 = RG_rl_176 ;
	7'h5b :
		rl_a94_t8 = RG_rl_176 ;
	7'h5c :
		rl_a94_t8 = RG_rl_176 ;
	7'h5d :
		rl_a94_t8 = RG_rl_176 ;
	7'h5e :
		rl_a94_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h5f :
		rl_a94_t8 = RG_rl_176 ;
	7'h60 :
		rl_a94_t8 = RG_rl_176 ;
	7'h61 :
		rl_a94_t8 = RG_rl_176 ;
	7'h62 :
		rl_a94_t8 = RG_rl_176 ;
	7'h63 :
		rl_a94_t8 = RG_rl_176 ;
	7'h64 :
		rl_a94_t8 = RG_rl_176 ;
	7'h65 :
		rl_a94_t8 = RG_rl_176 ;
	7'h66 :
		rl_a94_t8 = RG_rl_176 ;
	7'h67 :
		rl_a94_t8 = RG_rl_176 ;
	7'h68 :
		rl_a94_t8 = RG_rl_176 ;
	7'h69 :
		rl_a94_t8 = RG_rl_176 ;
	7'h6a :
		rl_a94_t8 = RG_rl_176 ;
	7'h6b :
		rl_a94_t8 = RG_rl_176 ;
	7'h6c :
		rl_a94_t8 = RG_rl_176 ;
	7'h6d :
		rl_a94_t8 = RG_rl_176 ;
	7'h6e :
		rl_a94_t8 = RG_rl_176 ;
	7'h6f :
		rl_a94_t8 = RG_rl_176 ;
	7'h70 :
		rl_a94_t8 = RG_rl_176 ;
	7'h71 :
		rl_a94_t8 = RG_rl_176 ;
	7'h72 :
		rl_a94_t8 = RG_rl_176 ;
	7'h73 :
		rl_a94_t8 = RG_rl_176 ;
	7'h74 :
		rl_a94_t8 = RG_rl_176 ;
	7'h75 :
		rl_a94_t8 = RG_rl_176 ;
	7'h76 :
		rl_a94_t8 = RG_rl_176 ;
	7'h77 :
		rl_a94_t8 = RG_rl_176 ;
	7'h78 :
		rl_a94_t8 = RG_rl_176 ;
	7'h79 :
		rl_a94_t8 = RG_rl_176 ;
	7'h7a :
		rl_a94_t8 = RG_rl_176 ;
	7'h7b :
		rl_a94_t8 = RG_rl_176 ;
	7'h7c :
		rl_a94_t8 = RG_rl_176 ;
	7'h7d :
		rl_a94_t8 = RG_rl_176 ;
	7'h7e :
		rl_a94_t8 = RG_rl_176 ;
	7'h7f :
		rl_a94_t8 = RG_rl_176 ;
	default :
		rl_a94_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_45 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h01 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h02 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h03 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h04 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h05 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h06 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h07 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h08 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h09 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h0a :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h0b :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h0c :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h0d :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h0e :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h0f :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h10 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h11 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h12 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h13 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h14 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h15 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h16 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h17 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h18 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h19 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h1a :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h1b :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h1c :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h1d :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h1e :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h1f :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h20 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h21 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h22 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h23 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h24 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h25 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h26 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h27 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h28 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h29 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h2a :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h2b :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h2c :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h2d :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h2e :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h2f :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h30 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h31 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h32 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h33 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h34 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h35 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h36 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h37 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h38 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h39 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h3a :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h3b :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h3c :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h3d :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h3e :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h3f :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h40 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h41 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h42 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h43 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h44 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h45 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h46 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h47 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h48 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h49 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h4a :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h4b :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h4c :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h4d :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h4e :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h4f :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h50 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h51 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h52 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h53 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h54 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h55 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h56 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h57 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h58 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h59 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h5a :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h5b :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h5c :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h5d :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h5e :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h5f :
		rl_a95_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h60 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h61 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h62 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h63 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h64 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h65 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h66 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h67 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h68 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h69 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h6a :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h6b :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h6c :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h6d :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h6e :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h6f :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h70 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h71 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h72 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h73 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h74 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h75 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h76 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h77 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h78 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h79 :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h7a :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h7b :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h7c :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h7d :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h7e :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	7'h7f :
		rl_a95_t8 = RG_quantized_block_rl_45 ;
	default :
		rl_a95_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_177 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a96_t8 = RG_rl_177 ;
	7'h01 :
		rl_a96_t8 = RG_rl_177 ;
	7'h02 :
		rl_a96_t8 = RG_rl_177 ;
	7'h03 :
		rl_a96_t8 = RG_rl_177 ;
	7'h04 :
		rl_a96_t8 = RG_rl_177 ;
	7'h05 :
		rl_a96_t8 = RG_rl_177 ;
	7'h06 :
		rl_a96_t8 = RG_rl_177 ;
	7'h07 :
		rl_a96_t8 = RG_rl_177 ;
	7'h08 :
		rl_a96_t8 = RG_rl_177 ;
	7'h09 :
		rl_a96_t8 = RG_rl_177 ;
	7'h0a :
		rl_a96_t8 = RG_rl_177 ;
	7'h0b :
		rl_a96_t8 = RG_rl_177 ;
	7'h0c :
		rl_a96_t8 = RG_rl_177 ;
	7'h0d :
		rl_a96_t8 = RG_rl_177 ;
	7'h0e :
		rl_a96_t8 = RG_rl_177 ;
	7'h0f :
		rl_a96_t8 = RG_rl_177 ;
	7'h10 :
		rl_a96_t8 = RG_rl_177 ;
	7'h11 :
		rl_a96_t8 = RG_rl_177 ;
	7'h12 :
		rl_a96_t8 = RG_rl_177 ;
	7'h13 :
		rl_a96_t8 = RG_rl_177 ;
	7'h14 :
		rl_a96_t8 = RG_rl_177 ;
	7'h15 :
		rl_a96_t8 = RG_rl_177 ;
	7'h16 :
		rl_a96_t8 = RG_rl_177 ;
	7'h17 :
		rl_a96_t8 = RG_rl_177 ;
	7'h18 :
		rl_a96_t8 = RG_rl_177 ;
	7'h19 :
		rl_a96_t8 = RG_rl_177 ;
	7'h1a :
		rl_a96_t8 = RG_rl_177 ;
	7'h1b :
		rl_a96_t8 = RG_rl_177 ;
	7'h1c :
		rl_a96_t8 = RG_rl_177 ;
	7'h1d :
		rl_a96_t8 = RG_rl_177 ;
	7'h1e :
		rl_a96_t8 = RG_rl_177 ;
	7'h1f :
		rl_a96_t8 = RG_rl_177 ;
	7'h20 :
		rl_a96_t8 = RG_rl_177 ;
	7'h21 :
		rl_a96_t8 = RG_rl_177 ;
	7'h22 :
		rl_a96_t8 = RG_rl_177 ;
	7'h23 :
		rl_a96_t8 = RG_rl_177 ;
	7'h24 :
		rl_a96_t8 = RG_rl_177 ;
	7'h25 :
		rl_a96_t8 = RG_rl_177 ;
	7'h26 :
		rl_a96_t8 = RG_rl_177 ;
	7'h27 :
		rl_a96_t8 = RG_rl_177 ;
	7'h28 :
		rl_a96_t8 = RG_rl_177 ;
	7'h29 :
		rl_a96_t8 = RG_rl_177 ;
	7'h2a :
		rl_a96_t8 = RG_rl_177 ;
	7'h2b :
		rl_a96_t8 = RG_rl_177 ;
	7'h2c :
		rl_a96_t8 = RG_rl_177 ;
	7'h2d :
		rl_a96_t8 = RG_rl_177 ;
	7'h2e :
		rl_a96_t8 = RG_rl_177 ;
	7'h2f :
		rl_a96_t8 = RG_rl_177 ;
	7'h30 :
		rl_a96_t8 = RG_rl_177 ;
	7'h31 :
		rl_a96_t8 = RG_rl_177 ;
	7'h32 :
		rl_a96_t8 = RG_rl_177 ;
	7'h33 :
		rl_a96_t8 = RG_rl_177 ;
	7'h34 :
		rl_a96_t8 = RG_rl_177 ;
	7'h35 :
		rl_a96_t8 = RG_rl_177 ;
	7'h36 :
		rl_a96_t8 = RG_rl_177 ;
	7'h37 :
		rl_a96_t8 = RG_rl_177 ;
	7'h38 :
		rl_a96_t8 = RG_rl_177 ;
	7'h39 :
		rl_a96_t8 = RG_rl_177 ;
	7'h3a :
		rl_a96_t8 = RG_rl_177 ;
	7'h3b :
		rl_a96_t8 = RG_rl_177 ;
	7'h3c :
		rl_a96_t8 = RG_rl_177 ;
	7'h3d :
		rl_a96_t8 = RG_rl_177 ;
	7'h3e :
		rl_a96_t8 = RG_rl_177 ;
	7'h3f :
		rl_a96_t8 = RG_rl_177 ;
	7'h40 :
		rl_a96_t8 = RG_rl_177 ;
	7'h41 :
		rl_a96_t8 = RG_rl_177 ;
	7'h42 :
		rl_a96_t8 = RG_rl_177 ;
	7'h43 :
		rl_a96_t8 = RG_rl_177 ;
	7'h44 :
		rl_a96_t8 = RG_rl_177 ;
	7'h45 :
		rl_a96_t8 = RG_rl_177 ;
	7'h46 :
		rl_a96_t8 = RG_rl_177 ;
	7'h47 :
		rl_a96_t8 = RG_rl_177 ;
	7'h48 :
		rl_a96_t8 = RG_rl_177 ;
	7'h49 :
		rl_a96_t8 = RG_rl_177 ;
	7'h4a :
		rl_a96_t8 = RG_rl_177 ;
	7'h4b :
		rl_a96_t8 = RG_rl_177 ;
	7'h4c :
		rl_a96_t8 = RG_rl_177 ;
	7'h4d :
		rl_a96_t8 = RG_rl_177 ;
	7'h4e :
		rl_a96_t8 = RG_rl_177 ;
	7'h4f :
		rl_a96_t8 = RG_rl_177 ;
	7'h50 :
		rl_a96_t8 = RG_rl_177 ;
	7'h51 :
		rl_a96_t8 = RG_rl_177 ;
	7'h52 :
		rl_a96_t8 = RG_rl_177 ;
	7'h53 :
		rl_a96_t8 = RG_rl_177 ;
	7'h54 :
		rl_a96_t8 = RG_rl_177 ;
	7'h55 :
		rl_a96_t8 = RG_rl_177 ;
	7'h56 :
		rl_a96_t8 = RG_rl_177 ;
	7'h57 :
		rl_a96_t8 = RG_rl_177 ;
	7'h58 :
		rl_a96_t8 = RG_rl_177 ;
	7'h59 :
		rl_a96_t8 = RG_rl_177 ;
	7'h5a :
		rl_a96_t8 = RG_rl_177 ;
	7'h5b :
		rl_a96_t8 = RG_rl_177 ;
	7'h5c :
		rl_a96_t8 = RG_rl_177 ;
	7'h5d :
		rl_a96_t8 = RG_rl_177 ;
	7'h5e :
		rl_a96_t8 = RG_rl_177 ;
	7'h5f :
		rl_a96_t8 = RG_rl_177 ;
	7'h60 :
		rl_a96_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h61 :
		rl_a96_t8 = RG_rl_177 ;
	7'h62 :
		rl_a96_t8 = RG_rl_177 ;
	7'h63 :
		rl_a96_t8 = RG_rl_177 ;
	7'h64 :
		rl_a96_t8 = RG_rl_177 ;
	7'h65 :
		rl_a96_t8 = RG_rl_177 ;
	7'h66 :
		rl_a96_t8 = RG_rl_177 ;
	7'h67 :
		rl_a96_t8 = RG_rl_177 ;
	7'h68 :
		rl_a96_t8 = RG_rl_177 ;
	7'h69 :
		rl_a96_t8 = RG_rl_177 ;
	7'h6a :
		rl_a96_t8 = RG_rl_177 ;
	7'h6b :
		rl_a96_t8 = RG_rl_177 ;
	7'h6c :
		rl_a96_t8 = RG_rl_177 ;
	7'h6d :
		rl_a96_t8 = RG_rl_177 ;
	7'h6e :
		rl_a96_t8 = RG_rl_177 ;
	7'h6f :
		rl_a96_t8 = RG_rl_177 ;
	7'h70 :
		rl_a96_t8 = RG_rl_177 ;
	7'h71 :
		rl_a96_t8 = RG_rl_177 ;
	7'h72 :
		rl_a96_t8 = RG_rl_177 ;
	7'h73 :
		rl_a96_t8 = RG_rl_177 ;
	7'h74 :
		rl_a96_t8 = RG_rl_177 ;
	7'h75 :
		rl_a96_t8 = RG_rl_177 ;
	7'h76 :
		rl_a96_t8 = RG_rl_177 ;
	7'h77 :
		rl_a96_t8 = RG_rl_177 ;
	7'h78 :
		rl_a96_t8 = RG_rl_177 ;
	7'h79 :
		rl_a96_t8 = RG_rl_177 ;
	7'h7a :
		rl_a96_t8 = RG_rl_177 ;
	7'h7b :
		rl_a96_t8 = RG_rl_177 ;
	7'h7c :
		rl_a96_t8 = RG_rl_177 ;
	7'h7d :
		rl_a96_t8 = RG_rl_177 ;
	7'h7e :
		rl_a96_t8 = RG_rl_177 ;
	7'h7f :
		rl_a96_t8 = RG_rl_177 ;
	default :
		rl_a96_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_46 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h01 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h02 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h03 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h04 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h05 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h06 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h07 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h08 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h09 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h0a :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h0b :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h0c :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h0d :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h0e :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h0f :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h10 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h11 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h12 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h13 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h14 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h15 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h16 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h17 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h18 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h19 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h1a :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h1b :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h1c :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h1d :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h1e :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h1f :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h20 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h21 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h22 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h23 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h24 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h25 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h26 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h27 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h28 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h29 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h2a :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h2b :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h2c :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h2d :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h2e :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h2f :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h30 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h31 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h32 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h33 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h34 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h35 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h36 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h37 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h38 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h39 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h3a :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h3b :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h3c :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h3d :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h3e :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h3f :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h40 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h41 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h42 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h43 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h44 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h45 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h46 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h47 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h48 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h49 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h4a :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h4b :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h4c :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h4d :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h4e :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h4f :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h50 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h51 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h52 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h53 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h54 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h55 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h56 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h57 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h58 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h59 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h5a :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h5b :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h5c :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h5d :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h5e :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h5f :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h60 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h61 :
		rl_a97_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h62 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h63 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h64 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h65 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h66 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h67 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h68 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h69 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h6a :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h6b :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h6c :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h6d :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h6e :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h6f :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h70 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h71 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h72 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h73 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h74 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h75 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h76 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h77 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h78 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h79 :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h7a :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h7b :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h7c :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h7d :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h7e :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	7'h7f :
		rl_a97_t8 = RG_quantized_block_rl_46 ;
	default :
		rl_a97_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_178 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a98_t8 = RG_rl_178 ;
	7'h01 :
		rl_a98_t8 = RG_rl_178 ;
	7'h02 :
		rl_a98_t8 = RG_rl_178 ;
	7'h03 :
		rl_a98_t8 = RG_rl_178 ;
	7'h04 :
		rl_a98_t8 = RG_rl_178 ;
	7'h05 :
		rl_a98_t8 = RG_rl_178 ;
	7'h06 :
		rl_a98_t8 = RG_rl_178 ;
	7'h07 :
		rl_a98_t8 = RG_rl_178 ;
	7'h08 :
		rl_a98_t8 = RG_rl_178 ;
	7'h09 :
		rl_a98_t8 = RG_rl_178 ;
	7'h0a :
		rl_a98_t8 = RG_rl_178 ;
	7'h0b :
		rl_a98_t8 = RG_rl_178 ;
	7'h0c :
		rl_a98_t8 = RG_rl_178 ;
	7'h0d :
		rl_a98_t8 = RG_rl_178 ;
	7'h0e :
		rl_a98_t8 = RG_rl_178 ;
	7'h0f :
		rl_a98_t8 = RG_rl_178 ;
	7'h10 :
		rl_a98_t8 = RG_rl_178 ;
	7'h11 :
		rl_a98_t8 = RG_rl_178 ;
	7'h12 :
		rl_a98_t8 = RG_rl_178 ;
	7'h13 :
		rl_a98_t8 = RG_rl_178 ;
	7'h14 :
		rl_a98_t8 = RG_rl_178 ;
	7'h15 :
		rl_a98_t8 = RG_rl_178 ;
	7'h16 :
		rl_a98_t8 = RG_rl_178 ;
	7'h17 :
		rl_a98_t8 = RG_rl_178 ;
	7'h18 :
		rl_a98_t8 = RG_rl_178 ;
	7'h19 :
		rl_a98_t8 = RG_rl_178 ;
	7'h1a :
		rl_a98_t8 = RG_rl_178 ;
	7'h1b :
		rl_a98_t8 = RG_rl_178 ;
	7'h1c :
		rl_a98_t8 = RG_rl_178 ;
	7'h1d :
		rl_a98_t8 = RG_rl_178 ;
	7'h1e :
		rl_a98_t8 = RG_rl_178 ;
	7'h1f :
		rl_a98_t8 = RG_rl_178 ;
	7'h20 :
		rl_a98_t8 = RG_rl_178 ;
	7'h21 :
		rl_a98_t8 = RG_rl_178 ;
	7'h22 :
		rl_a98_t8 = RG_rl_178 ;
	7'h23 :
		rl_a98_t8 = RG_rl_178 ;
	7'h24 :
		rl_a98_t8 = RG_rl_178 ;
	7'h25 :
		rl_a98_t8 = RG_rl_178 ;
	7'h26 :
		rl_a98_t8 = RG_rl_178 ;
	7'h27 :
		rl_a98_t8 = RG_rl_178 ;
	7'h28 :
		rl_a98_t8 = RG_rl_178 ;
	7'h29 :
		rl_a98_t8 = RG_rl_178 ;
	7'h2a :
		rl_a98_t8 = RG_rl_178 ;
	7'h2b :
		rl_a98_t8 = RG_rl_178 ;
	7'h2c :
		rl_a98_t8 = RG_rl_178 ;
	7'h2d :
		rl_a98_t8 = RG_rl_178 ;
	7'h2e :
		rl_a98_t8 = RG_rl_178 ;
	7'h2f :
		rl_a98_t8 = RG_rl_178 ;
	7'h30 :
		rl_a98_t8 = RG_rl_178 ;
	7'h31 :
		rl_a98_t8 = RG_rl_178 ;
	7'h32 :
		rl_a98_t8 = RG_rl_178 ;
	7'h33 :
		rl_a98_t8 = RG_rl_178 ;
	7'h34 :
		rl_a98_t8 = RG_rl_178 ;
	7'h35 :
		rl_a98_t8 = RG_rl_178 ;
	7'h36 :
		rl_a98_t8 = RG_rl_178 ;
	7'h37 :
		rl_a98_t8 = RG_rl_178 ;
	7'h38 :
		rl_a98_t8 = RG_rl_178 ;
	7'h39 :
		rl_a98_t8 = RG_rl_178 ;
	7'h3a :
		rl_a98_t8 = RG_rl_178 ;
	7'h3b :
		rl_a98_t8 = RG_rl_178 ;
	7'h3c :
		rl_a98_t8 = RG_rl_178 ;
	7'h3d :
		rl_a98_t8 = RG_rl_178 ;
	7'h3e :
		rl_a98_t8 = RG_rl_178 ;
	7'h3f :
		rl_a98_t8 = RG_rl_178 ;
	7'h40 :
		rl_a98_t8 = RG_rl_178 ;
	7'h41 :
		rl_a98_t8 = RG_rl_178 ;
	7'h42 :
		rl_a98_t8 = RG_rl_178 ;
	7'h43 :
		rl_a98_t8 = RG_rl_178 ;
	7'h44 :
		rl_a98_t8 = RG_rl_178 ;
	7'h45 :
		rl_a98_t8 = RG_rl_178 ;
	7'h46 :
		rl_a98_t8 = RG_rl_178 ;
	7'h47 :
		rl_a98_t8 = RG_rl_178 ;
	7'h48 :
		rl_a98_t8 = RG_rl_178 ;
	7'h49 :
		rl_a98_t8 = RG_rl_178 ;
	7'h4a :
		rl_a98_t8 = RG_rl_178 ;
	7'h4b :
		rl_a98_t8 = RG_rl_178 ;
	7'h4c :
		rl_a98_t8 = RG_rl_178 ;
	7'h4d :
		rl_a98_t8 = RG_rl_178 ;
	7'h4e :
		rl_a98_t8 = RG_rl_178 ;
	7'h4f :
		rl_a98_t8 = RG_rl_178 ;
	7'h50 :
		rl_a98_t8 = RG_rl_178 ;
	7'h51 :
		rl_a98_t8 = RG_rl_178 ;
	7'h52 :
		rl_a98_t8 = RG_rl_178 ;
	7'h53 :
		rl_a98_t8 = RG_rl_178 ;
	7'h54 :
		rl_a98_t8 = RG_rl_178 ;
	7'h55 :
		rl_a98_t8 = RG_rl_178 ;
	7'h56 :
		rl_a98_t8 = RG_rl_178 ;
	7'h57 :
		rl_a98_t8 = RG_rl_178 ;
	7'h58 :
		rl_a98_t8 = RG_rl_178 ;
	7'h59 :
		rl_a98_t8 = RG_rl_178 ;
	7'h5a :
		rl_a98_t8 = RG_rl_178 ;
	7'h5b :
		rl_a98_t8 = RG_rl_178 ;
	7'h5c :
		rl_a98_t8 = RG_rl_178 ;
	7'h5d :
		rl_a98_t8 = RG_rl_178 ;
	7'h5e :
		rl_a98_t8 = RG_rl_178 ;
	7'h5f :
		rl_a98_t8 = RG_rl_178 ;
	7'h60 :
		rl_a98_t8 = RG_rl_178 ;
	7'h61 :
		rl_a98_t8 = RG_rl_178 ;
	7'h62 :
		rl_a98_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h63 :
		rl_a98_t8 = RG_rl_178 ;
	7'h64 :
		rl_a98_t8 = RG_rl_178 ;
	7'h65 :
		rl_a98_t8 = RG_rl_178 ;
	7'h66 :
		rl_a98_t8 = RG_rl_178 ;
	7'h67 :
		rl_a98_t8 = RG_rl_178 ;
	7'h68 :
		rl_a98_t8 = RG_rl_178 ;
	7'h69 :
		rl_a98_t8 = RG_rl_178 ;
	7'h6a :
		rl_a98_t8 = RG_rl_178 ;
	7'h6b :
		rl_a98_t8 = RG_rl_178 ;
	7'h6c :
		rl_a98_t8 = RG_rl_178 ;
	7'h6d :
		rl_a98_t8 = RG_rl_178 ;
	7'h6e :
		rl_a98_t8 = RG_rl_178 ;
	7'h6f :
		rl_a98_t8 = RG_rl_178 ;
	7'h70 :
		rl_a98_t8 = RG_rl_178 ;
	7'h71 :
		rl_a98_t8 = RG_rl_178 ;
	7'h72 :
		rl_a98_t8 = RG_rl_178 ;
	7'h73 :
		rl_a98_t8 = RG_rl_178 ;
	7'h74 :
		rl_a98_t8 = RG_rl_178 ;
	7'h75 :
		rl_a98_t8 = RG_rl_178 ;
	7'h76 :
		rl_a98_t8 = RG_rl_178 ;
	7'h77 :
		rl_a98_t8 = RG_rl_178 ;
	7'h78 :
		rl_a98_t8 = RG_rl_178 ;
	7'h79 :
		rl_a98_t8 = RG_rl_178 ;
	7'h7a :
		rl_a98_t8 = RG_rl_178 ;
	7'h7b :
		rl_a98_t8 = RG_rl_178 ;
	7'h7c :
		rl_a98_t8 = RG_rl_178 ;
	7'h7d :
		rl_a98_t8 = RG_rl_178 ;
	7'h7e :
		rl_a98_t8 = RG_rl_178 ;
	7'h7f :
		rl_a98_t8 = RG_rl_178 ;
	default :
		rl_a98_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_47 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h01 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h02 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h03 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h04 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h05 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h06 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h07 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h08 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h09 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h0a :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h0b :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h0c :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h0d :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h0e :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h0f :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h10 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h11 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h12 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h13 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h14 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h15 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h16 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h17 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h18 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h19 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h1a :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h1b :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h1c :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h1d :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h1e :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h1f :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h20 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h21 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h22 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h23 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h24 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h25 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h26 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h27 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h28 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h29 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h2a :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h2b :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h2c :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h2d :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h2e :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h2f :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h30 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h31 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h32 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h33 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h34 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h35 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h36 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h37 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h38 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h39 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h3a :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h3b :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h3c :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h3d :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h3e :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h3f :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h40 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h41 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h42 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h43 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h44 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h45 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h46 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h47 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h48 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h49 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h4a :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h4b :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h4c :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h4d :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h4e :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h4f :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h50 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h51 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h52 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h53 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h54 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h55 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h56 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h57 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h58 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h59 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h5a :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h5b :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h5c :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h5d :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h5e :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h5f :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h60 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h61 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h62 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h63 :
		rl_a99_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h64 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h65 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h66 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h67 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h68 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h69 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h6a :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h6b :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h6c :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h6d :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h6e :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h6f :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h70 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h71 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h72 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h73 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h74 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h75 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h76 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h77 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h78 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h79 :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h7a :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h7b :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h7c :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h7d :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h7e :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	7'h7f :
		rl_a99_t8 = RG_quantized_block_rl_47 ;
	default :
		rl_a99_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_179 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a100_t8 = RG_rl_179 ;
	7'h01 :
		rl_a100_t8 = RG_rl_179 ;
	7'h02 :
		rl_a100_t8 = RG_rl_179 ;
	7'h03 :
		rl_a100_t8 = RG_rl_179 ;
	7'h04 :
		rl_a100_t8 = RG_rl_179 ;
	7'h05 :
		rl_a100_t8 = RG_rl_179 ;
	7'h06 :
		rl_a100_t8 = RG_rl_179 ;
	7'h07 :
		rl_a100_t8 = RG_rl_179 ;
	7'h08 :
		rl_a100_t8 = RG_rl_179 ;
	7'h09 :
		rl_a100_t8 = RG_rl_179 ;
	7'h0a :
		rl_a100_t8 = RG_rl_179 ;
	7'h0b :
		rl_a100_t8 = RG_rl_179 ;
	7'h0c :
		rl_a100_t8 = RG_rl_179 ;
	7'h0d :
		rl_a100_t8 = RG_rl_179 ;
	7'h0e :
		rl_a100_t8 = RG_rl_179 ;
	7'h0f :
		rl_a100_t8 = RG_rl_179 ;
	7'h10 :
		rl_a100_t8 = RG_rl_179 ;
	7'h11 :
		rl_a100_t8 = RG_rl_179 ;
	7'h12 :
		rl_a100_t8 = RG_rl_179 ;
	7'h13 :
		rl_a100_t8 = RG_rl_179 ;
	7'h14 :
		rl_a100_t8 = RG_rl_179 ;
	7'h15 :
		rl_a100_t8 = RG_rl_179 ;
	7'h16 :
		rl_a100_t8 = RG_rl_179 ;
	7'h17 :
		rl_a100_t8 = RG_rl_179 ;
	7'h18 :
		rl_a100_t8 = RG_rl_179 ;
	7'h19 :
		rl_a100_t8 = RG_rl_179 ;
	7'h1a :
		rl_a100_t8 = RG_rl_179 ;
	7'h1b :
		rl_a100_t8 = RG_rl_179 ;
	7'h1c :
		rl_a100_t8 = RG_rl_179 ;
	7'h1d :
		rl_a100_t8 = RG_rl_179 ;
	7'h1e :
		rl_a100_t8 = RG_rl_179 ;
	7'h1f :
		rl_a100_t8 = RG_rl_179 ;
	7'h20 :
		rl_a100_t8 = RG_rl_179 ;
	7'h21 :
		rl_a100_t8 = RG_rl_179 ;
	7'h22 :
		rl_a100_t8 = RG_rl_179 ;
	7'h23 :
		rl_a100_t8 = RG_rl_179 ;
	7'h24 :
		rl_a100_t8 = RG_rl_179 ;
	7'h25 :
		rl_a100_t8 = RG_rl_179 ;
	7'h26 :
		rl_a100_t8 = RG_rl_179 ;
	7'h27 :
		rl_a100_t8 = RG_rl_179 ;
	7'h28 :
		rl_a100_t8 = RG_rl_179 ;
	7'h29 :
		rl_a100_t8 = RG_rl_179 ;
	7'h2a :
		rl_a100_t8 = RG_rl_179 ;
	7'h2b :
		rl_a100_t8 = RG_rl_179 ;
	7'h2c :
		rl_a100_t8 = RG_rl_179 ;
	7'h2d :
		rl_a100_t8 = RG_rl_179 ;
	7'h2e :
		rl_a100_t8 = RG_rl_179 ;
	7'h2f :
		rl_a100_t8 = RG_rl_179 ;
	7'h30 :
		rl_a100_t8 = RG_rl_179 ;
	7'h31 :
		rl_a100_t8 = RG_rl_179 ;
	7'h32 :
		rl_a100_t8 = RG_rl_179 ;
	7'h33 :
		rl_a100_t8 = RG_rl_179 ;
	7'h34 :
		rl_a100_t8 = RG_rl_179 ;
	7'h35 :
		rl_a100_t8 = RG_rl_179 ;
	7'h36 :
		rl_a100_t8 = RG_rl_179 ;
	7'h37 :
		rl_a100_t8 = RG_rl_179 ;
	7'h38 :
		rl_a100_t8 = RG_rl_179 ;
	7'h39 :
		rl_a100_t8 = RG_rl_179 ;
	7'h3a :
		rl_a100_t8 = RG_rl_179 ;
	7'h3b :
		rl_a100_t8 = RG_rl_179 ;
	7'h3c :
		rl_a100_t8 = RG_rl_179 ;
	7'h3d :
		rl_a100_t8 = RG_rl_179 ;
	7'h3e :
		rl_a100_t8 = RG_rl_179 ;
	7'h3f :
		rl_a100_t8 = RG_rl_179 ;
	7'h40 :
		rl_a100_t8 = RG_rl_179 ;
	7'h41 :
		rl_a100_t8 = RG_rl_179 ;
	7'h42 :
		rl_a100_t8 = RG_rl_179 ;
	7'h43 :
		rl_a100_t8 = RG_rl_179 ;
	7'h44 :
		rl_a100_t8 = RG_rl_179 ;
	7'h45 :
		rl_a100_t8 = RG_rl_179 ;
	7'h46 :
		rl_a100_t8 = RG_rl_179 ;
	7'h47 :
		rl_a100_t8 = RG_rl_179 ;
	7'h48 :
		rl_a100_t8 = RG_rl_179 ;
	7'h49 :
		rl_a100_t8 = RG_rl_179 ;
	7'h4a :
		rl_a100_t8 = RG_rl_179 ;
	7'h4b :
		rl_a100_t8 = RG_rl_179 ;
	7'h4c :
		rl_a100_t8 = RG_rl_179 ;
	7'h4d :
		rl_a100_t8 = RG_rl_179 ;
	7'h4e :
		rl_a100_t8 = RG_rl_179 ;
	7'h4f :
		rl_a100_t8 = RG_rl_179 ;
	7'h50 :
		rl_a100_t8 = RG_rl_179 ;
	7'h51 :
		rl_a100_t8 = RG_rl_179 ;
	7'h52 :
		rl_a100_t8 = RG_rl_179 ;
	7'h53 :
		rl_a100_t8 = RG_rl_179 ;
	7'h54 :
		rl_a100_t8 = RG_rl_179 ;
	7'h55 :
		rl_a100_t8 = RG_rl_179 ;
	7'h56 :
		rl_a100_t8 = RG_rl_179 ;
	7'h57 :
		rl_a100_t8 = RG_rl_179 ;
	7'h58 :
		rl_a100_t8 = RG_rl_179 ;
	7'h59 :
		rl_a100_t8 = RG_rl_179 ;
	7'h5a :
		rl_a100_t8 = RG_rl_179 ;
	7'h5b :
		rl_a100_t8 = RG_rl_179 ;
	7'h5c :
		rl_a100_t8 = RG_rl_179 ;
	7'h5d :
		rl_a100_t8 = RG_rl_179 ;
	7'h5e :
		rl_a100_t8 = RG_rl_179 ;
	7'h5f :
		rl_a100_t8 = RG_rl_179 ;
	7'h60 :
		rl_a100_t8 = RG_rl_179 ;
	7'h61 :
		rl_a100_t8 = RG_rl_179 ;
	7'h62 :
		rl_a100_t8 = RG_rl_179 ;
	7'h63 :
		rl_a100_t8 = RG_rl_179 ;
	7'h64 :
		rl_a100_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h65 :
		rl_a100_t8 = RG_rl_179 ;
	7'h66 :
		rl_a100_t8 = RG_rl_179 ;
	7'h67 :
		rl_a100_t8 = RG_rl_179 ;
	7'h68 :
		rl_a100_t8 = RG_rl_179 ;
	7'h69 :
		rl_a100_t8 = RG_rl_179 ;
	7'h6a :
		rl_a100_t8 = RG_rl_179 ;
	7'h6b :
		rl_a100_t8 = RG_rl_179 ;
	7'h6c :
		rl_a100_t8 = RG_rl_179 ;
	7'h6d :
		rl_a100_t8 = RG_rl_179 ;
	7'h6e :
		rl_a100_t8 = RG_rl_179 ;
	7'h6f :
		rl_a100_t8 = RG_rl_179 ;
	7'h70 :
		rl_a100_t8 = RG_rl_179 ;
	7'h71 :
		rl_a100_t8 = RG_rl_179 ;
	7'h72 :
		rl_a100_t8 = RG_rl_179 ;
	7'h73 :
		rl_a100_t8 = RG_rl_179 ;
	7'h74 :
		rl_a100_t8 = RG_rl_179 ;
	7'h75 :
		rl_a100_t8 = RG_rl_179 ;
	7'h76 :
		rl_a100_t8 = RG_rl_179 ;
	7'h77 :
		rl_a100_t8 = RG_rl_179 ;
	7'h78 :
		rl_a100_t8 = RG_rl_179 ;
	7'h79 :
		rl_a100_t8 = RG_rl_179 ;
	7'h7a :
		rl_a100_t8 = RG_rl_179 ;
	7'h7b :
		rl_a100_t8 = RG_rl_179 ;
	7'h7c :
		rl_a100_t8 = RG_rl_179 ;
	7'h7d :
		rl_a100_t8 = RG_rl_179 ;
	7'h7e :
		rl_a100_t8 = RG_rl_179 ;
	7'h7f :
		rl_a100_t8 = RG_rl_179 ;
	default :
		rl_a100_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_48 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h01 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h02 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h03 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h04 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h05 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h06 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h07 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h08 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h09 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h0a :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h0b :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h0c :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h0d :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h0e :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h0f :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h10 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h11 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h12 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h13 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h14 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h15 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h16 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h17 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h18 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h19 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h1a :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h1b :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h1c :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h1d :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h1e :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h1f :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h20 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h21 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h22 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h23 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h24 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h25 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h26 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h27 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h28 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h29 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h2a :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h2b :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h2c :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h2d :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h2e :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h2f :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h30 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h31 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h32 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h33 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h34 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h35 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h36 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h37 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h38 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h39 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h3a :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h3b :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h3c :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h3d :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h3e :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h3f :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h40 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h41 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h42 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h43 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h44 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h45 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h46 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h47 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h48 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h49 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h4a :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h4b :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h4c :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h4d :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h4e :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h4f :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h50 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h51 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h52 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h53 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h54 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h55 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h56 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h57 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h58 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h59 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h5a :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h5b :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h5c :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h5d :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h5e :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h5f :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h60 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h61 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h62 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h63 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h64 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h65 :
		rl_a101_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h66 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h67 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h68 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h69 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h6a :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h6b :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h6c :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h6d :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h6e :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h6f :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h70 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h71 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h72 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h73 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h74 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h75 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h76 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h77 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h78 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h79 :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h7a :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h7b :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h7c :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h7d :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h7e :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	7'h7f :
		rl_a101_t8 = RG_quantized_block_rl_48 ;
	default :
		rl_a101_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_180 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a102_t8 = RG_rl_180 ;
	7'h01 :
		rl_a102_t8 = RG_rl_180 ;
	7'h02 :
		rl_a102_t8 = RG_rl_180 ;
	7'h03 :
		rl_a102_t8 = RG_rl_180 ;
	7'h04 :
		rl_a102_t8 = RG_rl_180 ;
	7'h05 :
		rl_a102_t8 = RG_rl_180 ;
	7'h06 :
		rl_a102_t8 = RG_rl_180 ;
	7'h07 :
		rl_a102_t8 = RG_rl_180 ;
	7'h08 :
		rl_a102_t8 = RG_rl_180 ;
	7'h09 :
		rl_a102_t8 = RG_rl_180 ;
	7'h0a :
		rl_a102_t8 = RG_rl_180 ;
	7'h0b :
		rl_a102_t8 = RG_rl_180 ;
	7'h0c :
		rl_a102_t8 = RG_rl_180 ;
	7'h0d :
		rl_a102_t8 = RG_rl_180 ;
	7'h0e :
		rl_a102_t8 = RG_rl_180 ;
	7'h0f :
		rl_a102_t8 = RG_rl_180 ;
	7'h10 :
		rl_a102_t8 = RG_rl_180 ;
	7'h11 :
		rl_a102_t8 = RG_rl_180 ;
	7'h12 :
		rl_a102_t8 = RG_rl_180 ;
	7'h13 :
		rl_a102_t8 = RG_rl_180 ;
	7'h14 :
		rl_a102_t8 = RG_rl_180 ;
	7'h15 :
		rl_a102_t8 = RG_rl_180 ;
	7'h16 :
		rl_a102_t8 = RG_rl_180 ;
	7'h17 :
		rl_a102_t8 = RG_rl_180 ;
	7'h18 :
		rl_a102_t8 = RG_rl_180 ;
	7'h19 :
		rl_a102_t8 = RG_rl_180 ;
	7'h1a :
		rl_a102_t8 = RG_rl_180 ;
	7'h1b :
		rl_a102_t8 = RG_rl_180 ;
	7'h1c :
		rl_a102_t8 = RG_rl_180 ;
	7'h1d :
		rl_a102_t8 = RG_rl_180 ;
	7'h1e :
		rl_a102_t8 = RG_rl_180 ;
	7'h1f :
		rl_a102_t8 = RG_rl_180 ;
	7'h20 :
		rl_a102_t8 = RG_rl_180 ;
	7'h21 :
		rl_a102_t8 = RG_rl_180 ;
	7'h22 :
		rl_a102_t8 = RG_rl_180 ;
	7'h23 :
		rl_a102_t8 = RG_rl_180 ;
	7'h24 :
		rl_a102_t8 = RG_rl_180 ;
	7'h25 :
		rl_a102_t8 = RG_rl_180 ;
	7'h26 :
		rl_a102_t8 = RG_rl_180 ;
	7'h27 :
		rl_a102_t8 = RG_rl_180 ;
	7'h28 :
		rl_a102_t8 = RG_rl_180 ;
	7'h29 :
		rl_a102_t8 = RG_rl_180 ;
	7'h2a :
		rl_a102_t8 = RG_rl_180 ;
	7'h2b :
		rl_a102_t8 = RG_rl_180 ;
	7'h2c :
		rl_a102_t8 = RG_rl_180 ;
	7'h2d :
		rl_a102_t8 = RG_rl_180 ;
	7'h2e :
		rl_a102_t8 = RG_rl_180 ;
	7'h2f :
		rl_a102_t8 = RG_rl_180 ;
	7'h30 :
		rl_a102_t8 = RG_rl_180 ;
	7'h31 :
		rl_a102_t8 = RG_rl_180 ;
	7'h32 :
		rl_a102_t8 = RG_rl_180 ;
	7'h33 :
		rl_a102_t8 = RG_rl_180 ;
	7'h34 :
		rl_a102_t8 = RG_rl_180 ;
	7'h35 :
		rl_a102_t8 = RG_rl_180 ;
	7'h36 :
		rl_a102_t8 = RG_rl_180 ;
	7'h37 :
		rl_a102_t8 = RG_rl_180 ;
	7'h38 :
		rl_a102_t8 = RG_rl_180 ;
	7'h39 :
		rl_a102_t8 = RG_rl_180 ;
	7'h3a :
		rl_a102_t8 = RG_rl_180 ;
	7'h3b :
		rl_a102_t8 = RG_rl_180 ;
	7'h3c :
		rl_a102_t8 = RG_rl_180 ;
	7'h3d :
		rl_a102_t8 = RG_rl_180 ;
	7'h3e :
		rl_a102_t8 = RG_rl_180 ;
	7'h3f :
		rl_a102_t8 = RG_rl_180 ;
	7'h40 :
		rl_a102_t8 = RG_rl_180 ;
	7'h41 :
		rl_a102_t8 = RG_rl_180 ;
	7'h42 :
		rl_a102_t8 = RG_rl_180 ;
	7'h43 :
		rl_a102_t8 = RG_rl_180 ;
	7'h44 :
		rl_a102_t8 = RG_rl_180 ;
	7'h45 :
		rl_a102_t8 = RG_rl_180 ;
	7'h46 :
		rl_a102_t8 = RG_rl_180 ;
	7'h47 :
		rl_a102_t8 = RG_rl_180 ;
	7'h48 :
		rl_a102_t8 = RG_rl_180 ;
	7'h49 :
		rl_a102_t8 = RG_rl_180 ;
	7'h4a :
		rl_a102_t8 = RG_rl_180 ;
	7'h4b :
		rl_a102_t8 = RG_rl_180 ;
	7'h4c :
		rl_a102_t8 = RG_rl_180 ;
	7'h4d :
		rl_a102_t8 = RG_rl_180 ;
	7'h4e :
		rl_a102_t8 = RG_rl_180 ;
	7'h4f :
		rl_a102_t8 = RG_rl_180 ;
	7'h50 :
		rl_a102_t8 = RG_rl_180 ;
	7'h51 :
		rl_a102_t8 = RG_rl_180 ;
	7'h52 :
		rl_a102_t8 = RG_rl_180 ;
	7'h53 :
		rl_a102_t8 = RG_rl_180 ;
	7'h54 :
		rl_a102_t8 = RG_rl_180 ;
	7'h55 :
		rl_a102_t8 = RG_rl_180 ;
	7'h56 :
		rl_a102_t8 = RG_rl_180 ;
	7'h57 :
		rl_a102_t8 = RG_rl_180 ;
	7'h58 :
		rl_a102_t8 = RG_rl_180 ;
	7'h59 :
		rl_a102_t8 = RG_rl_180 ;
	7'h5a :
		rl_a102_t8 = RG_rl_180 ;
	7'h5b :
		rl_a102_t8 = RG_rl_180 ;
	7'h5c :
		rl_a102_t8 = RG_rl_180 ;
	7'h5d :
		rl_a102_t8 = RG_rl_180 ;
	7'h5e :
		rl_a102_t8 = RG_rl_180 ;
	7'h5f :
		rl_a102_t8 = RG_rl_180 ;
	7'h60 :
		rl_a102_t8 = RG_rl_180 ;
	7'h61 :
		rl_a102_t8 = RG_rl_180 ;
	7'h62 :
		rl_a102_t8 = RG_rl_180 ;
	7'h63 :
		rl_a102_t8 = RG_rl_180 ;
	7'h64 :
		rl_a102_t8 = RG_rl_180 ;
	7'h65 :
		rl_a102_t8 = RG_rl_180 ;
	7'h66 :
		rl_a102_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h67 :
		rl_a102_t8 = RG_rl_180 ;
	7'h68 :
		rl_a102_t8 = RG_rl_180 ;
	7'h69 :
		rl_a102_t8 = RG_rl_180 ;
	7'h6a :
		rl_a102_t8 = RG_rl_180 ;
	7'h6b :
		rl_a102_t8 = RG_rl_180 ;
	7'h6c :
		rl_a102_t8 = RG_rl_180 ;
	7'h6d :
		rl_a102_t8 = RG_rl_180 ;
	7'h6e :
		rl_a102_t8 = RG_rl_180 ;
	7'h6f :
		rl_a102_t8 = RG_rl_180 ;
	7'h70 :
		rl_a102_t8 = RG_rl_180 ;
	7'h71 :
		rl_a102_t8 = RG_rl_180 ;
	7'h72 :
		rl_a102_t8 = RG_rl_180 ;
	7'h73 :
		rl_a102_t8 = RG_rl_180 ;
	7'h74 :
		rl_a102_t8 = RG_rl_180 ;
	7'h75 :
		rl_a102_t8 = RG_rl_180 ;
	7'h76 :
		rl_a102_t8 = RG_rl_180 ;
	7'h77 :
		rl_a102_t8 = RG_rl_180 ;
	7'h78 :
		rl_a102_t8 = RG_rl_180 ;
	7'h79 :
		rl_a102_t8 = RG_rl_180 ;
	7'h7a :
		rl_a102_t8 = RG_rl_180 ;
	7'h7b :
		rl_a102_t8 = RG_rl_180 ;
	7'h7c :
		rl_a102_t8 = RG_rl_180 ;
	7'h7d :
		rl_a102_t8 = RG_rl_180 ;
	7'h7e :
		rl_a102_t8 = RG_rl_180 ;
	7'h7f :
		rl_a102_t8 = RG_rl_180 ;
	default :
		rl_a102_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_49 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h01 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h02 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h03 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h04 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h05 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h06 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h07 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h08 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h09 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h0a :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h0b :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h0c :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h0d :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h0e :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h0f :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h10 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h11 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h12 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h13 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h14 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h15 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h16 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h17 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h18 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h19 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h1a :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h1b :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h1c :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h1d :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h1e :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h1f :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h20 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h21 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h22 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h23 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h24 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h25 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h26 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h27 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h28 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h29 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h2a :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h2b :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h2c :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h2d :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h2e :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h2f :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h30 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h31 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h32 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h33 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h34 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h35 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h36 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h37 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h38 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h39 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h3a :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h3b :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h3c :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h3d :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h3e :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h3f :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h40 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h41 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h42 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h43 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h44 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h45 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h46 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h47 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h48 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h49 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h4a :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h4b :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h4c :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h4d :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h4e :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h4f :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h50 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h51 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h52 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h53 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h54 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h55 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h56 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h57 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h58 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h59 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h5a :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h5b :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h5c :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h5d :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h5e :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h5f :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h60 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h61 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h62 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h63 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h64 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h65 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h66 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h67 :
		rl_a103_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h68 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h69 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h6a :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h6b :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h6c :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h6d :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h6e :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h6f :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h70 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h71 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h72 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h73 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h74 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h75 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h76 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h77 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h78 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h79 :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h7a :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h7b :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h7c :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h7d :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h7e :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	7'h7f :
		rl_a103_t8 = RG_quantized_block_rl_49 ;
	default :
		rl_a103_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_181 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a104_t8 = RG_rl_181 ;
	7'h01 :
		rl_a104_t8 = RG_rl_181 ;
	7'h02 :
		rl_a104_t8 = RG_rl_181 ;
	7'h03 :
		rl_a104_t8 = RG_rl_181 ;
	7'h04 :
		rl_a104_t8 = RG_rl_181 ;
	7'h05 :
		rl_a104_t8 = RG_rl_181 ;
	7'h06 :
		rl_a104_t8 = RG_rl_181 ;
	7'h07 :
		rl_a104_t8 = RG_rl_181 ;
	7'h08 :
		rl_a104_t8 = RG_rl_181 ;
	7'h09 :
		rl_a104_t8 = RG_rl_181 ;
	7'h0a :
		rl_a104_t8 = RG_rl_181 ;
	7'h0b :
		rl_a104_t8 = RG_rl_181 ;
	7'h0c :
		rl_a104_t8 = RG_rl_181 ;
	7'h0d :
		rl_a104_t8 = RG_rl_181 ;
	7'h0e :
		rl_a104_t8 = RG_rl_181 ;
	7'h0f :
		rl_a104_t8 = RG_rl_181 ;
	7'h10 :
		rl_a104_t8 = RG_rl_181 ;
	7'h11 :
		rl_a104_t8 = RG_rl_181 ;
	7'h12 :
		rl_a104_t8 = RG_rl_181 ;
	7'h13 :
		rl_a104_t8 = RG_rl_181 ;
	7'h14 :
		rl_a104_t8 = RG_rl_181 ;
	7'h15 :
		rl_a104_t8 = RG_rl_181 ;
	7'h16 :
		rl_a104_t8 = RG_rl_181 ;
	7'h17 :
		rl_a104_t8 = RG_rl_181 ;
	7'h18 :
		rl_a104_t8 = RG_rl_181 ;
	7'h19 :
		rl_a104_t8 = RG_rl_181 ;
	7'h1a :
		rl_a104_t8 = RG_rl_181 ;
	7'h1b :
		rl_a104_t8 = RG_rl_181 ;
	7'h1c :
		rl_a104_t8 = RG_rl_181 ;
	7'h1d :
		rl_a104_t8 = RG_rl_181 ;
	7'h1e :
		rl_a104_t8 = RG_rl_181 ;
	7'h1f :
		rl_a104_t8 = RG_rl_181 ;
	7'h20 :
		rl_a104_t8 = RG_rl_181 ;
	7'h21 :
		rl_a104_t8 = RG_rl_181 ;
	7'h22 :
		rl_a104_t8 = RG_rl_181 ;
	7'h23 :
		rl_a104_t8 = RG_rl_181 ;
	7'h24 :
		rl_a104_t8 = RG_rl_181 ;
	7'h25 :
		rl_a104_t8 = RG_rl_181 ;
	7'h26 :
		rl_a104_t8 = RG_rl_181 ;
	7'h27 :
		rl_a104_t8 = RG_rl_181 ;
	7'h28 :
		rl_a104_t8 = RG_rl_181 ;
	7'h29 :
		rl_a104_t8 = RG_rl_181 ;
	7'h2a :
		rl_a104_t8 = RG_rl_181 ;
	7'h2b :
		rl_a104_t8 = RG_rl_181 ;
	7'h2c :
		rl_a104_t8 = RG_rl_181 ;
	7'h2d :
		rl_a104_t8 = RG_rl_181 ;
	7'h2e :
		rl_a104_t8 = RG_rl_181 ;
	7'h2f :
		rl_a104_t8 = RG_rl_181 ;
	7'h30 :
		rl_a104_t8 = RG_rl_181 ;
	7'h31 :
		rl_a104_t8 = RG_rl_181 ;
	7'h32 :
		rl_a104_t8 = RG_rl_181 ;
	7'h33 :
		rl_a104_t8 = RG_rl_181 ;
	7'h34 :
		rl_a104_t8 = RG_rl_181 ;
	7'h35 :
		rl_a104_t8 = RG_rl_181 ;
	7'h36 :
		rl_a104_t8 = RG_rl_181 ;
	7'h37 :
		rl_a104_t8 = RG_rl_181 ;
	7'h38 :
		rl_a104_t8 = RG_rl_181 ;
	7'h39 :
		rl_a104_t8 = RG_rl_181 ;
	7'h3a :
		rl_a104_t8 = RG_rl_181 ;
	7'h3b :
		rl_a104_t8 = RG_rl_181 ;
	7'h3c :
		rl_a104_t8 = RG_rl_181 ;
	7'h3d :
		rl_a104_t8 = RG_rl_181 ;
	7'h3e :
		rl_a104_t8 = RG_rl_181 ;
	7'h3f :
		rl_a104_t8 = RG_rl_181 ;
	7'h40 :
		rl_a104_t8 = RG_rl_181 ;
	7'h41 :
		rl_a104_t8 = RG_rl_181 ;
	7'h42 :
		rl_a104_t8 = RG_rl_181 ;
	7'h43 :
		rl_a104_t8 = RG_rl_181 ;
	7'h44 :
		rl_a104_t8 = RG_rl_181 ;
	7'h45 :
		rl_a104_t8 = RG_rl_181 ;
	7'h46 :
		rl_a104_t8 = RG_rl_181 ;
	7'h47 :
		rl_a104_t8 = RG_rl_181 ;
	7'h48 :
		rl_a104_t8 = RG_rl_181 ;
	7'h49 :
		rl_a104_t8 = RG_rl_181 ;
	7'h4a :
		rl_a104_t8 = RG_rl_181 ;
	7'h4b :
		rl_a104_t8 = RG_rl_181 ;
	7'h4c :
		rl_a104_t8 = RG_rl_181 ;
	7'h4d :
		rl_a104_t8 = RG_rl_181 ;
	7'h4e :
		rl_a104_t8 = RG_rl_181 ;
	7'h4f :
		rl_a104_t8 = RG_rl_181 ;
	7'h50 :
		rl_a104_t8 = RG_rl_181 ;
	7'h51 :
		rl_a104_t8 = RG_rl_181 ;
	7'h52 :
		rl_a104_t8 = RG_rl_181 ;
	7'h53 :
		rl_a104_t8 = RG_rl_181 ;
	7'h54 :
		rl_a104_t8 = RG_rl_181 ;
	7'h55 :
		rl_a104_t8 = RG_rl_181 ;
	7'h56 :
		rl_a104_t8 = RG_rl_181 ;
	7'h57 :
		rl_a104_t8 = RG_rl_181 ;
	7'h58 :
		rl_a104_t8 = RG_rl_181 ;
	7'h59 :
		rl_a104_t8 = RG_rl_181 ;
	7'h5a :
		rl_a104_t8 = RG_rl_181 ;
	7'h5b :
		rl_a104_t8 = RG_rl_181 ;
	7'h5c :
		rl_a104_t8 = RG_rl_181 ;
	7'h5d :
		rl_a104_t8 = RG_rl_181 ;
	7'h5e :
		rl_a104_t8 = RG_rl_181 ;
	7'h5f :
		rl_a104_t8 = RG_rl_181 ;
	7'h60 :
		rl_a104_t8 = RG_rl_181 ;
	7'h61 :
		rl_a104_t8 = RG_rl_181 ;
	7'h62 :
		rl_a104_t8 = RG_rl_181 ;
	7'h63 :
		rl_a104_t8 = RG_rl_181 ;
	7'h64 :
		rl_a104_t8 = RG_rl_181 ;
	7'h65 :
		rl_a104_t8 = RG_rl_181 ;
	7'h66 :
		rl_a104_t8 = RG_rl_181 ;
	7'h67 :
		rl_a104_t8 = RG_rl_181 ;
	7'h68 :
		rl_a104_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h69 :
		rl_a104_t8 = RG_rl_181 ;
	7'h6a :
		rl_a104_t8 = RG_rl_181 ;
	7'h6b :
		rl_a104_t8 = RG_rl_181 ;
	7'h6c :
		rl_a104_t8 = RG_rl_181 ;
	7'h6d :
		rl_a104_t8 = RG_rl_181 ;
	7'h6e :
		rl_a104_t8 = RG_rl_181 ;
	7'h6f :
		rl_a104_t8 = RG_rl_181 ;
	7'h70 :
		rl_a104_t8 = RG_rl_181 ;
	7'h71 :
		rl_a104_t8 = RG_rl_181 ;
	7'h72 :
		rl_a104_t8 = RG_rl_181 ;
	7'h73 :
		rl_a104_t8 = RG_rl_181 ;
	7'h74 :
		rl_a104_t8 = RG_rl_181 ;
	7'h75 :
		rl_a104_t8 = RG_rl_181 ;
	7'h76 :
		rl_a104_t8 = RG_rl_181 ;
	7'h77 :
		rl_a104_t8 = RG_rl_181 ;
	7'h78 :
		rl_a104_t8 = RG_rl_181 ;
	7'h79 :
		rl_a104_t8 = RG_rl_181 ;
	7'h7a :
		rl_a104_t8 = RG_rl_181 ;
	7'h7b :
		rl_a104_t8 = RG_rl_181 ;
	7'h7c :
		rl_a104_t8 = RG_rl_181 ;
	7'h7d :
		rl_a104_t8 = RG_rl_181 ;
	7'h7e :
		rl_a104_t8 = RG_rl_181 ;
	7'h7f :
		rl_a104_t8 = RG_rl_181 ;
	default :
		rl_a104_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_50 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h01 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h02 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h03 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h04 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h05 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h06 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h07 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h08 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h09 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h0a :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h0b :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h0c :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h0d :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h0e :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h0f :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h10 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h11 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h12 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h13 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h14 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h15 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h16 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h17 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h18 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h19 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h1a :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h1b :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h1c :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h1d :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h1e :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h1f :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h20 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h21 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h22 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h23 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h24 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h25 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h26 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h27 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h28 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h29 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h2a :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h2b :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h2c :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h2d :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h2e :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h2f :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h30 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h31 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h32 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h33 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h34 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h35 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h36 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h37 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h38 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h39 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h3a :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h3b :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h3c :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h3d :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h3e :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h3f :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h40 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h41 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h42 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h43 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h44 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h45 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h46 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h47 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h48 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h49 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h4a :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h4b :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h4c :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h4d :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h4e :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h4f :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h50 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h51 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h52 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h53 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h54 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h55 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h56 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h57 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h58 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h59 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h5a :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h5b :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h5c :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h5d :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h5e :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h5f :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h60 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h61 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h62 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h63 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h64 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h65 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h66 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h67 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h68 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h69 :
		rl_a105_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h6a :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h6b :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h6c :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h6d :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h6e :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h6f :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h70 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h71 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h72 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h73 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h74 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h75 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h76 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h77 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h78 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h79 :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h7a :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h7b :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h7c :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h7d :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h7e :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	7'h7f :
		rl_a105_t8 = RG_quantized_block_rl_50 ;
	default :
		rl_a105_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_182 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a106_t8 = RG_rl_182 ;
	7'h01 :
		rl_a106_t8 = RG_rl_182 ;
	7'h02 :
		rl_a106_t8 = RG_rl_182 ;
	7'h03 :
		rl_a106_t8 = RG_rl_182 ;
	7'h04 :
		rl_a106_t8 = RG_rl_182 ;
	7'h05 :
		rl_a106_t8 = RG_rl_182 ;
	7'h06 :
		rl_a106_t8 = RG_rl_182 ;
	7'h07 :
		rl_a106_t8 = RG_rl_182 ;
	7'h08 :
		rl_a106_t8 = RG_rl_182 ;
	7'h09 :
		rl_a106_t8 = RG_rl_182 ;
	7'h0a :
		rl_a106_t8 = RG_rl_182 ;
	7'h0b :
		rl_a106_t8 = RG_rl_182 ;
	7'h0c :
		rl_a106_t8 = RG_rl_182 ;
	7'h0d :
		rl_a106_t8 = RG_rl_182 ;
	7'h0e :
		rl_a106_t8 = RG_rl_182 ;
	7'h0f :
		rl_a106_t8 = RG_rl_182 ;
	7'h10 :
		rl_a106_t8 = RG_rl_182 ;
	7'h11 :
		rl_a106_t8 = RG_rl_182 ;
	7'h12 :
		rl_a106_t8 = RG_rl_182 ;
	7'h13 :
		rl_a106_t8 = RG_rl_182 ;
	7'h14 :
		rl_a106_t8 = RG_rl_182 ;
	7'h15 :
		rl_a106_t8 = RG_rl_182 ;
	7'h16 :
		rl_a106_t8 = RG_rl_182 ;
	7'h17 :
		rl_a106_t8 = RG_rl_182 ;
	7'h18 :
		rl_a106_t8 = RG_rl_182 ;
	7'h19 :
		rl_a106_t8 = RG_rl_182 ;
	7'h1a :
		rl_a106_t8 = RG_rl_182 ;
	7'h1b :
		rl_a106_t8 = RG_rl_182 ;
	7'h1c :
		rl_a106_t8 = RG_rl_182 ;
	7'h1d :
		rl_a106_t8 = RG_rl_182 ;
	7'h1e :
		rl_a106_t8 = RG_rl_182 ;
	7'h1f :
		rl_a106_t8 = RG_rl_182 ;
	7'h20 :
		rl_a106_t8 = RG_rl_182 ;
	7'h21 :
		rl_a106_t8 = RG_rl_182 ;
	7'h22 :
		rl_a106_t8 = RG_rl_182 ;
	7'h23 :
		rl_a106_t8 = RG_rl_182 ;
	7'h24 :
		rl_a106_t8 = RG_rl_182 ;
	7'h25 :
		rl_a106_t8 = RG_rl_182 ;
	7'h26 :
		rl_a106_t8 = RG_rl_182 ;
	7'h27 :
		rl_a106_t8 = RG_rl_182 ;
	7'h28 :
		rl_a106_t8 = RG_rl_182 ;
	7'h29 :
		rl_a106_t8 = RG_rl_182 ;
	7'h2a :
		rl_a106_t8 = RG_rl_182 ;
	7'h2b :
		rl_a106_t8 = RG_rl_182 ;
	7'h2c :
		rl_a106_t8 = RG_rl_182 ;
	7'h2d :
		rl_a106_t8 = RG_rl_182 ;
	7'h2e :
		rl_a106_t8 = RG_rl_182 ;
	7'h2f :
		rl_a106_t8 = RG_rl_182 ;
	7'h30 :
		rl_a106_t8 = RG_rl_182 ;
	7'h31 :
		rl_a106_t8 = RG_rl_182 ;
	7'h32 :
		rl_a106_t8 = RG_rl_182 ;
	7'h33 :
		rl_a106_t8 = RG_rl_182 ;
	7'h34 :
		rl_a106_t8 = RG_rl_182 ;
	7'h35 :
		rl_a106_t8 = RG_rl_182 ;
	7'h36 :
		rl_a106_t8 = RG_rl_182 ;
	7'h37 :
		rl_a106_t8 = RG_rl_182 ;
	7'h38 :
		rl_a106_t8 = RG_rl_182 ;
	7'h39 :
		rl_a106_t8 = RG_rl_182 ;
	7'h3a :
		rl_a106_t8 = RG_rl_182 ;
	7'h3b :
		rl_a106_t8 = RG_rl_182 ;
	7'h3c :
		rl_a106_t8 = RG_rl_182 ;
	7'h3d :
		rl_a106_t8 = RG_rl_182 ;
	7'h3e :
		rl_a106_t8 = RG_rl_182 ;
	7'h3f :
		rl_a106_t8 = RG_rl_182 ;
	7'h40 :
		rl_a106_t8 = RG_rl_182 ;
	7'h41 :
		rl_a106_t8 = RG_rl_182 ;
	7'h42 :
		rl_a106_t8 = RG_rl_182 ;
	7'h43 :
		rl_a106_t8 = RG_rl_182 ;
	7'h44 :
		rl_a106_t8 = RG_rl_182 ;
	7'h45 :
		rl_a106_t8 = RG_rl_182 ;
	7'h46 :
		rl_a106_t8 = RG_rl_182 ;
	7'h47 :
		rl_a106_t8 = RG_rl_182 ;
	7'h48 :
		rl_a106_t8 = RG_rl_182 ;
	7'h49 :
		rl_a106_t8 = RG_rl_182 ;
	7'h4a :
		rl_a106_t8 = RG_rl_182 ;
	7'h4b :
		rl_a106_t8 = RG_rl_182 ;
	7'h4c :
		rl_a106_t8 = RG_rl_182 ;
	7'h4d :
		rl_a106_t8 = RG_rl_182 ;
	7'h4e :
		rl_a106_t8 = RG_rl_182 ;
	7'h4f :
		rl_a106_t8 = RG_rl_182 ;
	7'h50 :
		rl_a106_t8 = RG_rl_182 ;
	7'h51 :
		rl_a106_t8 = RG_rl_182 ;
	7'h52 :
		rl_a106_t8 = RG_rl_182 ;
	7'h53 :
		rl_a106_t8 = RG_rl_182 ;
	7'h54 :
		rl_a106_t8 = RG_rl_182 ;
	7'h55 :
		rl_a106_t8 = RG_rl_182 ;
	7'h56 :
		rl_a106_t8 = RG_rl_182 ;
	7'h57 :
		rl_a106_t8 = RG_rl_182 ;
	7'h58 :
		rl_a106_t8 = RG_rl_182 ;
	7'h59 :
		rl_a106_t8 = RG_rl_182 ;
	7'h5a :
		rl_a106_t8 = RG_rl_182 ;
	7'h5b :
		rl_a106_t8 = RG_rl_182 ;
	7'h5c :
		rl_a106_t8 = RG_rl_182 ;
	7'h5d :
		rl_a106_t8 = RG_rl_182 ;
	7'h5e :
		rl_a106_t8 = RG_rl_182 ;
	7'h5f :
		rl_a106_t8 = RG_rl_182 ;
	7'h60 :
		rl_a106_t8 = RG_rl_182 ;
	7'h61 :
		rl_a106_t8 = RG_rl_182 ;
	7'h62 :
		rl_a106_t8 = RG_rl_182 ;
	7'h63 :
		rl_a106_t8 = RG_rl_182 ;
	7'h64 :
		rl_a106_t8 = RG_rl_182 ;
	7'h65 :
		rl_a106_t8 = RG_rl_182 ;
	7'h66 :
		rl_a106_t8 = RG_rl_182 ;
	7'h67 :
		rl_a106_t8 = RG_rl_182 ;
	7'h68 :
		rl_a106_t8 = RG_rl_182 ;
	7'h69 :
		rl_a106_t8 = RG_rl_182 ;
	7'h6a :
		rl_a106_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h6b :
		rl_a106_t8 = RG_rl_182 ;
	7'h6c :
		rl_a106_t8 = RG_rl_182 ;
	7'h6d :
		rl_a106_t8 = RG_rl_182 ;
	7'h6e :
		rl_a106_t8 = RG_rl_182 ;
	7'h6f :
		rl_a106_t8 = RG_rl_182 ;
	7'h70 :
		rl_a106_t8 = RG_rl_182 ;
	7'h71 :
		rl_a106_t8 = RG_rl_182 ;
	7'h72 :
		rl_a106_t8 = RG_rl_182 ;
	7'h73 :
		rl_a106_t8 = RG_rl_182 ;
	7'h74 :
		rl_a106_t8 = RG_rl_182 ;
	7'h75 :
		rl_a106_t8 = RG_rl_182 ;
	7'h76 :
		rl_a106_t8 = RG_rl_182 ;
	7'h77 :
		rl_a106_t8 = RG_rl_182 ;
	7'h78 :
		rl_a106_t8 = RG_rl_182 ;
	7'h79 :
		rl_a106_t8 = RG_rl_182 ;
	7'h7a :
		rl_a106_t8 = RG_rl_182 ;
	7'h7b :
		rl_a106_t8 = RG_rl_182 ;
	7'h7c :
		rl_a106_t8 = RG_rl_182 ;
	7'h7d :
		rl_a106_t8 = RG_rl_182 ;
	7'h7e :
		rl_a106_t8 = RG_rl_182 ;
	7'h7f :
		rl_a106_t8 = RG_rl_182 ;
	default :
		rl_a106_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_51 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h01 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h02 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h03 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h04 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h05 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h06 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h07 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h08 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h09 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h0a :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h0b :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h0c :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h0d :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h0e :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h0f :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h10 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h11 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h12 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h13 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h14 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h15 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h16 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h17 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h18 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h19 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h1a :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h1b :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h1c :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h1d :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h1e :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h1f :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h20 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h21 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h22 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h23 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h24 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h25 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h26 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h27 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h28 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h29 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h2a :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h2b :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h2c :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h2d :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h2e :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h2f :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h30 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h31 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h32 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h33 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h34 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h35 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h36 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h37 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h38 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h39 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h3a :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h3b :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h3c :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h3d :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h3e :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h3f :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h40 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h41 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h42 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h43 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h44 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h45 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h46 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h47 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h48 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h49 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h4a :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h4b :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h4c :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h4d :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h4e :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h4f :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h50 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h51 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h52 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h53 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h54 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h55 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h56 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h57 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h58 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h59 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h5a :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h5b :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h5c :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h5d :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h5e :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h5f :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h60 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h61 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h62 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h63 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h64 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h65 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h66 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h67 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h68 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h69 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h6a :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h6b :
		rl_a107_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h6c :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h6d :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h6e :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h6f :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h70 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h71 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h72 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h73 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h74 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h75 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h76 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h77 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h78 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h79 :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h7a :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h7b :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h7c :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h7d :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h7e :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	7'h7f :
		rl_a107_t8 = RG_quantized_block_rl_51 ;
	default :
		rl_a107_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_183 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a108_t8 = RG_rl_183 ;
	7'h01 :
		rl_a108_t8 = RG_rl_183 ;
	7'h02 :
		rl_a108_t8 = RG_rl_183 ;
	7'h03 :
		rl_a108_t8 = RG_rl_183 ;
	7'h04 :
		rl_a108_t8 = RG_rl_183 ;
	7'h05 :
		rl_a108_t8 = RG_rl_183 ;
	7'h06 :
		rl_a108_t8 = RG_rl_183 ;
	7'h07 :
		rl_a108_t8 = RG_rl_183 ;
	7'h08 :
		rl_a108_t8 = RG_rl_183 ;
	7'h09 :
		rl_a108_t8 = RG_rl_183 ;
	7'h0a :
		rl_a108_t8 = RG_rl_183 ;
	7'h0b :
		rl_a108_t8 = RG_rl_183 ;
	7'h0c :
		rl_a108_t8 = RG_rl_183 ;
	7'h0d :
		rl_a108_t8 = RG_rl_183 ;
	7'h0e :
		rl_a108_t8 = RG_rl_183 ;
	7'h0f :
		rl_a108_t8 = RG_rl_183 ;
	7'h10 :
		rl_a108_t8 = RG_rl_183 ;
	7'h11 :
		rl_a108_t8 = RG_rl_183 ;
	7'h12 :
		rl_a108_t8 = RG_rl_183 ;
	7'h13 :
		rl_a108_t8 = RG_rl_183 ;
	7'h14 :
		rl_a108_t8 = RG_rl_183 ;
	7'h15 :
		rl_a108_t8 = RG_rl_183 ;
	7'h16 :
		rl_a108_t8 = RG_rl_183 ;
	7'h17 :
		rl_a108_t8 = RG_rl_183 ;
	7'h18 :
		rl_a108_t8 = RG_rl_183 ;
	7'h19 :
		rl_a108_t8 = RG_rl_183 ;
	7'h1a :
		rl_a108_t8 = RG_rl_183 ;
	7'h1b :
		rl_a108_t8 = RG_rl_183 ;
	7'h1c :
		rl_a108_t8 = RG_rl_183 ;
	7'h1d :
		rl_a108_t8 = RG_rl_183 ;
	7'h1e :
		rl_a108_t8 = RG_rl_183 ;
	7'h1f :
		rl_a108_t8 = RG_rl_183 ;
	7'h20 :
		rl_a108_t8 = RG_rl_183 ;
	7'h21 :
		rl_a108_t8 = RG_rl_183 ;
	7'h22 :
		rl_a108_t8 = RG_rl_183 ;
	7'h23 :
		rl_a108_t8 = RG_rl_183 ;
	7'h24 :
		rl_a108_t8 = RG_rl_183 ;
	7'h25 :
		rl_a108_t8 = RG_rl_183 ;
	7'h26 :
		rl_a108_t8 = RG_rl_183 ;
	7'h27 :
		rl_a108_t8 = RG_rl_183 ;
	7'h28 :
		rl_a108_t8 = RG_rl_183 ;
	7'h29 :
		rl_a108_t8 = RG_rl_183 ;
	7'h2a :
		rl_a108_t8 = RG_rl_183 ;
	7'h2b :
		rl_a108_t8 = RG_rl_183 ;
	7'h2c :
		rl_a108_t8 = RG_rl_183 ;
	7'h2d :
		rl_a108_t8 = RG_rl_183 ;
	7'h2e :
		rl_a108_t8 = RG_rl_183 ;
	7'h2f :
		rl_a108_t8 = RG_rl_183 ;
	7'h30 :
		rl_a108_t8 = RG_rl_183 ;
	7'h31 :
		rl_a108_t8 = RG_rl_183 ;
	7'h32 :
		rl_a108_t8 = RG_rl_183 ;
	7'h33 :
		rl_a108_t8 = RG_rl_183 ;
	7'h34 :
		rl_a108_t8 = RG_rl_183 ;
	7'h35 :
		rl_a108_t8 = RG_rl_183 ;
	7'h36 :
		rl_a108_t8 = RG_rl_183 ;
	7'h37 :
		rl_a108_t8 = RG_rl_183 ;
	7'h38 :
		rl_a108_t8 = RG_rl_183 ;
	7'h39 :
		rl_a108_t8 = RG_rl_183 ;
	7'h3a :
		rl_a108_t8 = RG_rl_183 ;
	7'h3b :
		rl_a108_t8 = RG_rl_183 ;
	7'h3c :
		rl_a108_t8 = RG_rl_183 ;
	7'h3d :
		rl_a108_t8 = RG_rl_183 ;
	7'h3e :
		rl_a108_t8 = RG_rl_183 ;
	7'h3f :
		rl_a108_t8 = RG_rl_183 ;
	7'h40 :
		rl_a108_t8 = RG_rl_183 ;
	7'h41 :
		rl_a108_t8 = RG_rl_183 ;
	7'h42 :
		rl_a108_t8 = RG_rl_183 ;
	7'h43 :
		rl_a108_t8 = RG_rl_183 ;
	7'h44 :
		rl_a108_t8 = RG_rl_183 ;
	7'h45 :
		rl_a108_t8 = RG_rl_183 ;
	7'h46 :
		rl_a108_t8 = RG_rl_183 ;
	7'h47 :
		rl_a108_t8 = RG_rl_183 ;
	7'h48 :
		rl_a108_t8 = RG_rl_183 ;
	7'h49 :
		rl_a108_t8 = RG_rl_183 ;
	7'h4a :
		rl_a108_t8 = RG_rl_183 ;
	7'h4b :
		rl_a108_t8 = RG_rl_183 ;
	7'h4c :
		rl_a108_t8 = RG_rl_183 ;
	7'h4d :
		rl_a108_t8 = RG_rl_183 ;
	7'h4e :
		rl_a108_t8 = RG_rl_183 ;
	7'h4f :
		rl_a108_t8 = RG_rl_183 ;
	7'h50 :
		rl_a108_t8 = RG_rl_183 ;
	7'h51 :
		rl_a108_t8 = RG_rl_183 ;
	7'h52 :
		rl_a108_t8 = RG_rl_183 ;
	7'h53 :
		rl_a108_t8 = RG_rl_183 ;
	7'h54 :
		rl_a108_t8 = RG_rl_183 ;
	7'h55 :
		rl_a108_t8 = RG_rl_183 ;
	7'h56 :
		rl_a108_t8 = RG_rl_183 ;
	7'h57 :
		rl_a108_t8 = RG_rl_183 ;
	7'h58 :
		rl_a108_t8 = RG_rl_183 ;
	7'h59 :
		rl_a108_t8 = RG_rl_183 ;
	7'h5a :
		rl_a108_t8 = RG_rl_183 ;
	7'h5b :
		rl_a108_t8 = RG_rl_183 ;
	7'h5c :
		rl_a108_t8 = RG_rl_183 ;
	7'h5d :
		rl_a108_t8 = RG_rl_183 ;
	7'h5e :
		rl_a108_t8 = RG_rl_183 ;
	7'h5f :
		rl_a108_t8 = RG_rl_183 ;
	7'h60 :
		rl_a108_t8 = RG_rl_183 ;
	7'h61 :
		rl_a108_t8 = RG_rl_183 ;
	7'h62 :
		rl_a108_t8 = RG_rl_183 ;
	7'h63 :
		rl_a108_t8 = RG_rl_183 ;
	7'h64 :
		rl_a108_t8 = RG_rl_183 ;
	7'h65 :
		rl_a108_t8 = RG_rl_183 ;
	7'h66 :
		rl_a108_t8 = RG_rl_183 ;
	7'h67 :
		rl_a108_t8 = RG_rl_183 ;
	7'h68 :
		rl_a108_t8 = RG_rl_183 ;
	7'h69 :
		rl_a108_t8 = RG_rl_183 ;
	7'h6a :
		rl_a108_t8 = RG_rl_183 ;
	7'h6b :
		rl_a108_t8 = RG_rl_183 ;
	7'h6c :
		rl_a108_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h6d :
		rl_a108_t8 = RG_rl_183 ;
	7'h6e :
		rl_a108_t8 = RG_rl_183 ;
	7'h6f :
		rl_a108_t8 = RG_rl_183 ;
	7'h70 :
		rl_a108_t8 = RG_rl_183 ;
	7'h71 :
		rl_a108_t8 = RG_rl_183 ;
	7'h72 :
		rl_a108_t8 = RG_rl_183 ;
	7'h73 :
		rl_a108_t8 = RG_rl_183 ;
	7'h74 :
		rl_a108_t8 = RG_rl_183 ;
	7'h75 :
		rl_a108_t8 = RG_rl_183 ;
	7'h76 :
		rl_a108_t8 = RG_rl_183 ;
	7'h77 :
		rl_a108_t8 = RG_rl_183 ;
	7'h78 :
		rl_a108_t8 = RG_rl_183 ;
	7'h79 :
		rl_a108_t8 = RG_rl_183 ;
	7'h7a :
		rl_a108_t8 = RG_rl_183 ;
	7'h7b :
		rl_a108_t8 = RG_rl_183 ;
	7'h7c :
		rl_a108_t8 = RG_rl_183 ;
	7'h7d :
		rl_a108_t8 = RG_rl_183 ;
	7'h7e :
		rl_a108_t8 = RG_rl_183 ;
	7'h7f :
		rl_a108_t8 = RG_rl_183 ;
	default :
		rl_a108_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_52 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h01 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h02 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h03 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h04 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h05 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h06 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h07 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h08 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h09 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h0a :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h0b :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h0c :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h0d :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h0e :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h0f :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h10 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h11 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h12 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h13 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h14 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h15 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h16 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h17 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h18 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h19 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h1a :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h1b :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h1c :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h1d :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h1e :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h1f :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h20 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h21 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h22 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h23 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h24 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h25 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h26 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h27 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h28 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h29 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h2a :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h2b :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h2c :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h2d :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h2e :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h2f :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h30 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h31 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h32 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h33 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h34 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h35 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h36 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h37 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h38 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h39 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h3a :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h3b :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h3c :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h3d :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h3e :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h3f :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h40 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h41 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h42 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h43 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h44 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h45 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h46 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h47 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h48 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h49 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h4a :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h4b :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h4c :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h4d :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h4e :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h4f :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h50 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h51 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h52 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h53 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h54 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h55 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h56 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h57 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h58 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h59 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h5a :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h5b :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h5c :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h5d :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h5e :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h5f :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h60 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h61 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h62 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h63 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h64 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h65 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h66 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h67 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h68 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h69 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h6a :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h6b :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h6c :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h6d :
		rl_a109_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h6e :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h6f :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h70 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h71 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h72 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h73 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h74 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h75 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h76 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h77 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h78 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h79 :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h7a :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h7b :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h7c :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h7d :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h7e :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	7'h7f :
		rl_a109_t8 = RG_quantized_block_rl_52 ;
	default :
		rl_a109_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_184 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a110_t8 = RG_rl_184 ;
	7'h01 :
		rl_a110_t8 = RG_rl_184 ;
	7'h02 :
		rl_a110_t8 = RG_rl_184 ;
	7'h03 :
		rl_a110_t8 = RG_rl_184 ;
	7'h04 :
		rl_a110_t8 = RG_rl_184 ;
	7'h05 :
		rl_a110_t8 = RG_rl_184 ;
	7'h06 :
		rl_a110_t8 = RG_rl_184 ;
	7'h07 :
		rl_a110_t8 = RG_rl_184 ;
	7'h08 :
		rl_a110_t8 = RG_rl_184 ;
	7'h09 :
		rl_a110_t8 = RG_rl_184 ;
	7'h0a :
		rl_a110_t8 = RG_rl_184 ;
	7'h0b :
		rl_a110_t8 = RG_rl_184 ;
	7'h0c :
		rl_a110_t8 = RG_rl_184 ;
	7'h0d :
		rl_a110_t8 = RG_rl_184 ;
	7'h0e :
		rl_a110_t8 = RG_rl_184 ;
	7'h0f :
		rl_a110_t8 = RG_rl_184 ;
	7'h10 :
		rl_a110_t8 = RG_rl_184 ;
	7'h11 :
		rl_a110_t8 = RG_rl_184 ;
	7'h12 :
		rl_a110_t8 = RG_rl_184 ;
	7'h13 :
		rl_a110_t8 = RG_rl_184 ;
	7'h14 :
		rl_a110_t8 = RG_rl_184 ;
	7'h15 :
		rl_a110_t8 = RG_rl_184 ;
	7'h16 :
		rl_a110_t8 = RG_rl_184 ;
	7'h17 :
		rl_a110_t8 = RG_rl_184 ;
	7'h18 :
		rl_a110_t8 = RG_rl_184 ;
	7'h19 :
		rl_a110_t8 = RG_rl_184 ;
	7'h1a :
		rl_a110_t8 = RG_rl_184 ;
	7'h1b :
		rl_a110_t8 = RG_rl_184 ;
	7'h1c :
		rl_a110_t8 = RG_rl_184 ;
	7'h1d :
		rl_a110_t8 = RG_rl_184 ;
	7'h1e :
		rl_a110_t8 = RG_rl_184 ;
	7'h1f :
		rl_a110_t8 = RG_rl_184 ;
	7'h20 :
		rl_a110_t8 = RG_rl_184 ;
	7'h21 :
		rl_a110_t8 = RG_rl_184 ;
	7'h22 :
		rl_a110_t8 = RG_rl_184 ;
	7'h23 :
		rl_a110_t8 = RG_rl_184 ;
	7'h24 :
		rl_a110_t8 = RG_rl_184 ;
	7'h25 :
		rl_a110_t8 = RG_rl_184 ;
	7'h26 :
		rl_a110_t8 = RG_rl_184 ;
	7'h27 :
		rl_a110_t8 = RG_rl_184 ;
	7'h28 :
		rl_a110_t8 = RG_rl_184 ;
	7'h29 :
		rl_a110_t8 = RG_rl_184 ;
	7'h2a :
		rl_a110_t8 = RG_rl_184 ;
	7'h2b :
		rl_a110_t8 = RG_rl_184 ;
	7'h2c :
		rl_a110_t8 = RG_rl_184 ;
	7'h2d :
		rl_a110_t8 = RG_rl_184 ;
	7'h2e :
		rl_a110_t8 = RG_rl_184 ;
	7'h2f :
		rl_a110_t8 = RG_rl_184 ;
	7'h30 :
		rl_a110_t8 = RG_rl_184 ;
	7'h31 :
		rl_a110_t8 = RG_rl_184 ;
	7'h32 :
		rl_a110_t8 = RG_rl_184 ;
	7'h33 :
		rl_a110_t8 = RG_rl_184 ;
	7'h34 :
		rl_a110_t8 = RG_rl_184 ;
	7'h35 :
		rl_a110_t8 = RG_rl_184 ;
	7'h36 :
		rl_a110_t8 = RG_rl_184 ;
	7'h37 :
		rl_a110_t8 = RG_rl_184 ;
	7'h38 :
		rl_a110_t8 = RG_rl_184 ;
	7'h39 :
		rl_a110_t8 = RG_rl_184 ;
	7'h3a :
		rl_a110_t8 = RG_rl_184 ;
	7'h3b :
		rl_a110_t8 = RG_rl_184 ;
	7'h3c :
		rl_a110_t8 = RG_rl_184 ;
	7'h3d :
		rl_a110_t8 = RG_rl_184 ;
	7'h3e :
		rl_a110_t8 = RG_rl_184 ;
	7'h3f :
		rl_a110_t8 = RG_rl_184 ;
	7'h40 :
		rl_a110_t8 = RG_rl_184 ;
	7'h41 :
		rl_a110_t8 = RG_rl_184 ;
	7'h42 :
		rl_a110_t8 = RG_rl_184 ;
	7'h43 :
		rl_a110_t8 = RG_rl_184 ;
	7'h44 :
		rl_a110_t8 = RG_rl_184 ;
	7'h45 :
		rl_a110_t8 = RG_rl_184 ;
	7'h46 :
		rl_a110_t8 = RG_rl_184 ;
	7'h47 :
		rl_a110_t8 = RG_rl_184 ;
	7'h48 :
		rl_a110_t8 = RG_rl_184 ;
	7'h49 :
		rl_a110_t8 = RG_rl_184 ;
	7'h4a :
		rl_a110_t8 = RG_rl_184 ;
	7'h4b :
		rl_a110_t8 = RG_rl_184 ;
	7'h4c :
		rl_a110_t8 = RG_rl_184 ;
	7'h4d :
		rl_a110_t8 = RG_rl_184 ;
	7'h4e :
		rl_a110_t8 = RG_rl_184 ;
	7'h4f :
		rl_a110_t8 = RG_rl_184 ;
	7'h50 :
		rl_a110_t8 = RG_rl_184 ;
	7'h51 :
		rl_a110_t8 = RG_rl_184 ;
	7'h52 :
		rl_a110_t8 = RG_rl_184 ;
	7'h53 :
		rl_a110_t8 = RG_rl_184 ;
	7'h54 :
		rl_a110_t8 = RG_rl_184 ;
	7'h55 :
		rl_a110_t8 = RG_rl_184 ;
	7'h56 :
		rl_a110_t8 = RG_rl_184 ;
	7'h57 :
		rl_a110_t8 = RG_rl_184 ;
	7'h58 :
		rl_a110_t8 = RG_rl_184 ;
	7'h59 :
		rl_a110_t8 = RG_rl_184 ;
	7'h5a :
		rl_a110_t8 = RG_rl_184 ;
	7'h5b :
		rl_a110_t8 = RG_rl_184 ;
	7'h5c :
		rl_a110_t8 = RG_rl_184 ;
	7'h5d :
		rl_a110_t8 = RG_rl_184 ;
	7'h5e :
		rl_a110_t8 = RG_rl_184 ;
	7'h5f :
		rl_a110_t8 = RG_rl_184 ;
	7'h60 :
		rl_a110_t8 = RG_rl_184 ;
	7'h61 :
		rl_a110_t8 = RG_rl_184 ;
	7'h62 :
		rl_a110_t8 = RG_rl_184 ;
	7'h63 :
		rl_a110_t8 = RG_rl_184 ;
	7'h64 :
		rl_a110_t8 = RG_rl_184 ;
	7'h65 :
		rl_a110_t8 = RG_rl_184 ;
	7'h66 :
		rl_a110_t8 = RG_rl_184 ;
	7'h67 :
		rl_a110_t8 = RG_rl_184 ;
	7'h68 :
		rl_a110_t8 = RG_rl_184 ;
	7'h69 :
		rl_a110_t8 = RG_rl_184 ;
	7'h6a :
		rl_a110_t8 = RG_rl_184 ;
	7'h6b :
		rl_a110_t8 = RG_rl_184 ;
	7'h6c :
		rl_a110_t8 = RG_rl_184 ;
	7'h6d :
		rl_a110_t8 = RG_rl_184 ;
	7'h6e :
		rl_a110_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h6f :
		rl_a110_t8 = RG_rl_184 ;
	7'h70 :
		rl_a110_t8 = RG_rl_184 ;
	7'h71 :
		rl_a110_t8 = RG_rl_184 ;
	7'h72 :
		rl_a110_t8 = RG_rl_184 ;
	7'h73 :
		rl_a110_t8 = RG_rl_184 ;
	7'h74 :
		rl_a110_t8 = RG_rl_184 ;
	7'h75 :
		rl_a110_t8 = RG_rl_184 ;
	7'h76 :
		rl_a110_t8 = RG_rl_184 ;
	7'h77 :
		rl_a110_t8 = RG_rl_184 ;
	7'h78 :
		rl_a110_t8 = RG_rl_184 ;
	7'h79 :
		rl_a110_t8 = RG_rl_184 ;
	7'h7a :
		rl_a110_t8 = RG_rl_184 ;
	7'h7b :
		rl_a110_t8 = RG_rl_184 ;
	7'h7c :
		rl_a110_t8 = RG_rl_184 ;
	7'h7d :
		rl_a110_t8 = RG_rl_184 ;
	7'h7e :
		rl_a110_t8 = RG_rl_184 ;
	7'h7f :
		rl_a110_t8 = RG_rl_184 ;
	default :
		rl_a110_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_53 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h01 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h02 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h03 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h04 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h05 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h06 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h07 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h08 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h09 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h0a :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h0b :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h0c :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h0d :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h0e :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h0f :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h10 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h11 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h12 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h13 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h14 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h15 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h16 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h17 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h18 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h19 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h1a :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h1b :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h1c :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h1d :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h1e :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h1f :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h20 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h21 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h22 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h23 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h24 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h25 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h26 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h27 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h28 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h29 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h2a :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h2b :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h2c :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h2d :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h2e :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h2f :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h30 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h31 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h32 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h33 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h34 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h35 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h36 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h37 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h38 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h39 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h3a :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h3b :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h3c :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h3d :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h3e :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h3f :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h40 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h41 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h42 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h43 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h44 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h45 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h46 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h47 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h48 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h49 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h4a :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h4b :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h4c :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h4d :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h4e :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h4f :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h50 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h51 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h52 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h53 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h54 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h55 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h56 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h57 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h58 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h59 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h5a :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h5b :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h5c :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h5d :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h5e :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h5f :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h60 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h61 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h62 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h63 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h64 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h65 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h66 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h67 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h68 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h69 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h6a :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h6b :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h6c :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h6d :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h6e :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h6f :
		rl_a111_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h70 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h71 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h72 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h73 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h74 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h75 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h76 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h77 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h78 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h79 :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h7a :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h7b :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h7c :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h7d :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h7e :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	7'h7f :
		rl_a111_t8 = RG_quantized_block_rl_53 ;
	default :
		rl_a111_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_185 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a112_t8 = RG_rl_185 ;
	7'h01 :
		rl_a112_t8 = RG_rl_185 ;
	7'h02 :
		rl_a112_t8 = RG_rl_185 ;
	7'h03 :
		rl_a112_t8 = RG_rl_185 ;
	7'h04 :
		rl_a112_t8 = RG_rl_185 ;
	7'h05 :
		rl_a112_t8 = RG_rl_185 ;
	7'h06 :
		rl_a112_t8 = RG_rl_185 ;
	7'h07 :
		rl_a112_t8 = RG_rl_185 ;
	7'h08 :
		rl_a112_t8 = RG_rl_185 ;
	7'h09 :
		rl_a112_t8 = RG_rl_185 ;
	7'h0a :
		rl_a112_t8 = RG_rl_185 ;
	7'h0b :
		rl_a112_t8 = RG_rl_185 ;
	7'h0c :
		rl_a112_t8 = RG_rl_185 ;
	7'h0d :
		rl_a112_t8 = RG_rl_185 ;
	7'h0e :
		rl_a112_t8 = RG_rl_185 ;
	7'h0f :
		rl_a112_t8 = RG_rl_185 ;
	7'h10 :
		rl_a112_t8 = RG_rl_185 ;
	7'h11 :
		rl_a112_t8 = RG_rl_185 ;
	7'h12 :
		rl_a112_t8 = RG_rl_185 ;
	7'h13 :
		rl_a112_t8 = RG_rl_185 ;
	7'h14 :
		rl_a112_t8 = RG_rl_185 ;
	7'h15 :
		rl_a112_t8 = RG_rl_185 ;
	7'h16 :
		rl_a112_t8 = RG_rl_185 ;
	7'h17 :
		rl_a112_t8 = RG_rl_185 ;
	7'h18 :
		rl_a112_t8 = RG_rl_185 ;
	7'h19 :
		rl_a112_t8 = RG_rl_185 ;
	7'h1a :
		rl_a112_t8 = RG_rl_185 ;
	7'h1b :
		rl_a112_t8 = RG_rl_185 ;
	7'h1c :
		rl_a112_t8 = RG_rl_185 ;
	7'h1d :
		rl_a112_t8 = RG_rl_185 ;
	7'h1e :
		rl_a112_t8 = RG_rl_185 ;
	7'h1f :
		rl_a112_t8 = RG_rl_185 ;
	7'h20 :
		rl_a112_t8 = RG_rl_185 ;
	7'h21 :
		rl_a112_t8 = RG_rl_185 ;
	7'h22 :
		rl_a112_t8 = RG_rl_185 ;
	7'h23 :
		rl_a112_t8 = RG_rl_185 ;
	7'h24 :
		rl_a112_t8 = RG_rl_185 ;
	7'h25 :
		rl_a112_t8 = RG_rl_185 ;
	7'h26 :
		rl_a112_t8 = RG_rl_185 ;
	7'h27 :
		rl_a112_t8 = RG_rl_185 ;
	7'h28 :
		rl_a112_t8 = RG_rl_185 ;
	7'h29 :
		rl_a112_t8 = RG_rl_185 ;
	7'h2a :
		rl_a112_t8 = RG_rl_185 ;
	7'h2b :
		rl_a112_t8 = RG_rl_185 ;
	7'h2c :
		rl_a112_t8 = RG_rl_185 ;
	7'h2d :
		rl_a112_t8 = RG_rl_185 ;
	7'h2e :
		rl_a112_t8 = RG_rl_185 ;
	7'h2f :
		rl_a112_t8 = RG_rl_185 ;
	7'h30 :
		rl_a112_t8 = RG_rl_185 ;
	7'h31 :
		rl_a112_t8 = RG_rl_185 ;
	7'h32 :
		rl_a112_t8 = RG_rl_185 ;
	7'h33 :
		rl_a112_t8 = RG_rl_185 ;
	7'h34 :
		rl_a112_t8 = RG_rl_185 ;
	7'h35 :
		rl_a112_t8 = RG_rl_185 ;
	7'h36 :
		rl_a112_t8 = RG_rl_185 ;
	7'h37 :
		rl_a112_t8 = RG_rl_185 ;
	7'h38 :
		rl_a112_t8 = RG_rl_185 ;
	7'h39 :
		rl_a112_t8 = RG_rl_185 ;
	7'h3a :
		rl_a112_t8 = RG_rl_185 ;
	7'h3b :
		rl_a112_t8 = RG_rl_185 ;
	7'h3c :
		rl_a112_t8 = RG_rl_185 ;
	7'h3d :
		rl_a112_t8 = RG_rl_185 ;
	7'h3e :
		rl_a112_t8 = RG_rl_185 ;
	7'h3f :
		rl_a112_t8 = RG_rl_185 ;
	7'h40 :
		rl_a112_t8 = RG_rl_185 ;
	7'h41 :
		rl_a112_t8 = RG_rl_185 ;
	7'h42 :
		rl_a112_t8 = RG_rl_185 ;
	7'h43 :
		rl_a112_t8 = RG_rl_185 ;
	7'h44 :
		rl_a112_t8 = RG_rl_185 ;
	7'h45 :
		rl_a112_t8 = RG_rl_185 ;
	7'h46 :
		rl_a112_t8 = RG_rl_185 ;
	7'h47 :
		rl_a112_t8 = RG_rl_185 ;
	7'h48 :
		rl_a112_t8 = RG_rl_185 ;
	7'h49 :
		rl_a112_t8 = RG_rl_185 ;
	7'h4a :
		rl_a112_t8 = RG_rl_185 ;
	7'h4b :
		rl_a112_t8 = RG_rl_185 ;
	7'h4c :
		rl_a112_t8 = RG_rl_185 ;
	7'h4d :
		rl_a112_t8 = RG_rl_185 ;
	7'h4e :
		rl_a112_t8 = RG_rl_185 ;
	7'h4f :
		rl_a112_t8 = RG_rl_185 ;
	7'h50 :
		rl_a112_t8 = RG_rl_185 ;
	7'h51 :
		rl_a112_t8 = RG_rl_185 ;
	7'h52 :
		rl_a112_t8 = RG_rl_185 ;
	7'h53 :
		rl_a112_t8 = RG_rl_185 ;
	7'h54 :
		rl_a112_t8 = RG_rl_185 ;
	7'h55 :
		rl_a112_t8 = RG_rl_185 ;
	7'h56 :
		rl_a112_t8 = RG_rl_185 ;
	7'h57 :
		rl_a112_t8 = RG_rl_185 ;
	7'h58 :
		rl_a112_t8 = RG_rl_185 ;
	7'h59 :
		rl_a112_t8 = RG_rl_185 ;
	7'h5a :
		rl_a112_t8 = RG_rl_185 ;
	7'h5b :
		rl_a112_t8 = RG_rl_185 ;
	7'h5c :
		rl_a112_t8 = RG_rl_185 ;
	7'h5d :
		rl_a112_t8 = RG_rl_185 ;
	7'h5e :
		rl_a112_t8 = RG_rl_185 ;
	7'h5f :
		rl_a112_t8 = RG_rl_185 ;
	7'h60 :
		rl_a112_t8 = RG_rl_185 ;
	7'h61 :
		rl_a112_t8 = RG_rl_185 ;
	7'h62 :
		rl_a112_t8 = RG_rl_185 ;
	7'h63 :
		rl_a112_t8 = RG_rl_185 ;
	7'h64 :
		rl_a112_t8 = RG_rl_185 ;
	7'h65 :
		rl_a112_t8 = RG_rl_185 ;
	7'h66 :
		rl_a112_t8 = RG_rl_185 ;
	7'h67 :
		rl_a112_t8 = RG_rl_185 ;
	7'h68 :
		rl_a112_t8 = RG_rl_185 ;
	7'h69 :
		rl_a112_t8 = RG_rl_185 ;
	7'h6a :
		rl_a112_t8 = RG_rl_185 ;
	7'h6b :
		rl_a112_t8 = RG_rl_185 ;
	7'h6c :
		rl_a112_t8 = RG_rl_185 ;
	7'h6d :
		rl_a112_t8 = RG_rl_185 ;
	7'h6e :
		rl_a112_t8 = RG_rl_185 ;
	7'h6f :
		rl_a112_t8 = RG_rl_185 ;
	7'h70 :
		rl_a112_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h71 :
		rl_a112_t8 = RG_rl_185 ;
	7'h72 :
		rl_a112_t8 = RG_rl_185 ;
	7'h73 :
		rl_a112_t8 = RG_rl_185 ;
	7'h74 :
		rl_a112_t8 = RG_rl_185 ;
	7'h75 :
		rl_a112_t8 = RG_rl_185 ;
	7'h76 :
		rl_a112_t8 = RG_rl_185 ;
	7'h77 :
		rl_a112_t8 = RG_rl_185 ;
	7'h78 :
		rl_a112_t8 = RG_rl_185 ;
	7'h79 :
		rl_a112_t8 = RG_rl_185 ;
	7'h7a :
		rl_a112_t8 = RG_rl_185 ;
	7'h7b :
		rl_a112_t8 = RG_rl_185 ;
	7'h7c :
		rl_a112_t8 = RG_rl_185 ;
	7'h7d :
		rl_a112_t8 = RG_rl_185 ;
	7'h7e :
		rl_a112_t8 = RG_rl_185 ;
	7'h7f :
		rl_a112_t8 = RG_rl_185 ;
	default :
		rl_a112_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_54 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h01 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h02 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h03 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h04 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h05 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h06 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h07 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h08 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h09 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h0a :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h0b :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h0c :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h0d :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h0e :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h0f :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h10 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h11 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h12 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h13 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h14 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h15 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h16 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h17 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h18 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h19 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h1a :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h1b :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h1c :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h1d :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h1e :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h1f :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h20 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h21 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h22 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h23 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h24 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h25 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h26 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h27 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h28 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h29 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h2a :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h2b :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h2c :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h2d :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h2e :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h2f :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h30 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h31 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h32 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h33 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h34 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h35 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h36 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h37 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h38 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h39 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h3a :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h3b :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h3c :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h3d :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h3e :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h3f :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h40 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h41 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h42 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h43 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h44 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h45 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h46 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h47 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h48 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h49 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h4a :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h4b :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h4c :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h4d :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h4e :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h4f :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h50 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h51 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h52 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h53 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h54 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h55 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h56 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h57 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h58 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h59 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h5a :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h5b :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h5c :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h5d :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h5e :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h5f :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h60 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h61 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h62 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h63 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h64 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h65 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h66 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h67 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h68 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h69 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h6a :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h6b :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h6c :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h6d :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h6e :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h6f :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h70 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h71 :
		rl_a113_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h72 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h73 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h74 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h75 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h76 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h77 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h78 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h79 :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h7a :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h7b :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h7c :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h7d :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h7e :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	7'h7f :
		rl_a113_t8 = RG_quantized_block_rl_54 ;
	default :
		rl_a113_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_186 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a114_t8 = RG_rl_186 ;
	7'h01 :
		rl_a114_t8 = RG_rl_186 ;
	7'h02 :
		rl_a114_t8 = RG_rl_186 ;
	7'h03 :
		rl_a114_t8 = RG_rl_186 ;
	7'h04 :
		rl_a114_t8 = RG_rl_186 ;
	7'h05 :
		rl_a114_t8 = RG_rl_186 ;
	7'h06 :
		rl_a114_t8 = RG_rl_186 ;
	7'h07 :
		rl_a114_t8 = RG_rl_186 ;
	7'h08 :
		rl_a114_t8 = RG_rl_186 ;
	7'h09 :
		rl_a114_t8 = RG_rl_186 ;
	7'h0a :
		rl_a114_t8 = RG_rl_186 ;
	7'h0b :
		rl_a114_t8 = RG_rl_186 ;
	7'h0c :
		rl_a114_t8 = RG_rl_186 ;
	7'h0d :
		rl_a114_t8 = RG_rl_186 ;
	7'h0e :
		rl_a114_t8 = RG_rl_186 ;
	7'h0f :
		rl_a114_t8 = RG_rl_186 ;
	7'h10 :
		rl_a114_t8 = RG_rl_186 ;
	7'h11 :
		rl_a114_t8 = RG_rl_186 ;
	7'h12 :
		rl_a114_t8 = RG_rl_186 ;
	7'h13 :
		rl_a114_t8 = RG_rl_186 ;
	7'h14 :
		rl_a114_t8 = RG_rl_186 ;
	7'h15 :
		rl_a114_t8 = RG_rl_186 ;
	7'h16 :
		rl_a114_t8 = RG_rl_186 ;
	7'h17 :
		rl_a114_t8 = RG_rl_186 ;
	7'h18 :
		rl_a114_t8 = RG_rl_186 ;
	7'h19 :
		rl_a114_t8 = RG_rl_186 ;
	7'h1a :
		rl_a114_t8 = RG_rl_186 ;
	7'h1b :
		rl_a114_t8 = RG_rl_186 ;
	7'h1c :
		rl_a114_t8 = RG_rl_186 ;
	7'h1d :
		rl_a114_t8 = RG_rl_186 ;
	7'h1e :
		rl_a114_t8 = RG_rl_186 ;
	7'h1f :
		rl_a114_t8 = RG_rl_186 ;
	7'h20 :
		rl_a114_t8 = RG_rl_186 ;
	7'h21 :
		rl_a114_t8 = RG_rl_186 ;
	7'h22 :
		rl_a114_t8 = RG_rl_186 ;
	7'h23 :
		rl_a114_t8 = RG_rl_186 ;
	7'h24 :
		rl_a114_t8 = RG_rl_186 ;
	7'h25 :
		rl_a114_t8 = RG_rl_186 ;
	7'h26 :
		rl_a114_t8 = RG_rl_186 ;
	7'h27 :
		rl_a114_t8 = RG_rl_186 ;
	7'h28 :
		rl_a114_t8 = RG_rl_186 ;
	7'h29 :
		rl_a114_t8 = RG_rl_186 ;
	7'h2a :
		rl_a114_t8 = RG_rl_186 ;
	7'h2b :
		rl_a114_t8 = RG_rl_186 ;
	7'h2c :
		rl_a114_t8 = RG_rl_186 ;
	7'h2d :
		rl_a114_t8 = RG_rl_186 ;
	7'h2e :
		rl_a114_t8 = RG_rl_186 ;
	7'h2f :
		rl_a114_t8 = RG_rl_186 ;
	7'h30 :
		rl_a114_t8 = RG_rl_186 ;
	7'h31 :
		rl_a114_t8 = RG_rl_186 ;
	7'h32 :
		rl_a114_t8 = RG_rl_186 ;
	7'h33 :
		rl_a114_t8 = RG_rl_186 ;
	7'h34 :
		rl_a114_t8 = RG_rl_186 ;
	7'h35 :
		rl_a114_t8 = RG_rl_186 ;
	7'h36 :
		rl_a114_t8 = RG_rl_186 ;
	7'h37 :
		rl_a114_t8 = RG_rl_186 ;
	7'h38 :
		rl_a114_t8 = RG_rl_186 ;
	7'h39 :
		rl_a114_t8 = RG_rl_186 ;
	7'h3a :
		rl_a114_t8 = RG_rl_186 ;
	7'h3b :
		rl_a114_t8 = RG_rl_186 ;
	7'h3c :
		rl_a114_t8 = RG_rl_186 ;
	7'h3d :
		rl_a114_t8 = RG_rl_186 ;
	7'h3e :
		rl_a114_t8 = RG_rl_186 ;
	7'h3f :
		rl_a114_t8 = RG_rl_186 ;
	7'h40 :
		rl_a114_t8 = RG_rl_186 ;
	7'h41 :
		rl_a114_t8 = RG_rl_186 ;
	7'h42 :
		rl_a114_t8 = RG_rl_186 ;
	7'h43 :
		rl_a114_t8 = RG_rl_186 ;
	7'h44 :
		rl_a114_t8 = RG_rl_186 ;
	7'h45 :
		rl_a114_t8 = RG_rl_186 ;
	7'h46 :
		rl_a114_t8 = RG_rl_186 ;
	7'h47 :
		rl_a114_t8 = RG_rl_186 ;
	7'h48 :
		rl_a114_t8 = RG_rl_186 ;
	7'h49 :
		rl_a114_t8 = RG_rl_186 ;
	7'h4a :
		rl_a114_t8 = RG_rl_186 ;
	7'h4b :
		rl_a114_t8 = RG_rl_186 ;
	7'h4c :
		rl_a114_t8 = RG_rl_186 ;
	7'h4d :
		rl_a114_t8 = RG_rl_186 ;
	7'h4e :
		rl_a114_t8 = RG_rl_186 ;
	7'h4f :
		rl_a114_t8 = RG_rl_186 ;
	7'h50 :
		rl_a114_t8 = RG_rl_186 ;
	7'h51 :
		rl_a114_t8 = RG_rl_186 ;
	7'h52 :
		rl_a114_t8 = RG_rl_186 ;
	7'h53 :
		rl_a114_t8 = RG_rl_186 ;
	7'h54 :
		rl_a114_t8 = RG_rl_186 ;
	7'h55 :
		rl_a114_t8 = RG_rl_186 ;
	7'h56 :
		rl_a114_t8 = RG_rl_186 ;
	7'h57 :
		rl_a114_t8 = RG_rl_186 ;
	7'h58 :
		rl_a114_t8 = RG_rl_186 ;
	7'h59 :
		rl_a114_t8 = RG_rl_186 ;
	7'h5a :
		rl_a114_t8 = RG_rl_186 ;
	7'h5b :
		rl_a114_t8 = RG_rl_186 ;
	7'h5c :
		rl_a114_t8 = RG_rl_186 ;
	7'h5d :
		rl_a114_t8 = RG_rl_186 ;
	7'h5e :
		rl_a114_t8 = RG_rl_186 ;
	7'h5f :
		rl_a114_t8 = RG_rl_186 ;
	7'h60 :
		rl_a114_t8 = RG_rl_186 ;
	7'h61 :
		rl_a114_t8 = RG_rl_186 ;
	7'h62 :
		rl_a114_t8 = RG_rl_186 ;
	7'h63 :
		rl_a114_t8 = RG_rl_186 ;
	7'h64 :
		rl_a114_t8 = RG_rl_186 ;
	7'h65 :
		rl_a114_t8 = RG_rl_186 ;
	7'h66 :
		rl_a114_t8 = RG_rl_186 ;
	7'h67 :
		rl_a114_t8 = RG_rl_186 ;
	7'h68 :
		rl_a114_t8 = RG_rl_186 ;
	7'h69 :
		rl_a114_t8 = RG_rl_186 ;
	7'h6a :
		rl_a114_t8 = RG_rl_186 ;
	7'h6b :
		rl_a114_t8 = RG_rl_186 ;
	7'h6c :
		rl_a114_t8 = RG_rl_186 ;
	7'h6d :
		rl_a114_t8 = RG_rl_186 ;
	7'h6e :
		rl_a114_t8 = RG_rl_186 ;
	7'h6f :
		rl_a114_t8 = RG_rl_186 ;
	7'h70 :
		rl_a114_t8 = RG_rl_186 ;
	7'h71 :
		rl_a114_t8 = RG_rl_186 ;
	7'h72 :
		rl_a114_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h73 :
		rl_a114_t8 = RG_rl_186 ;
	7'h74 :
		rl_a114_t8 = RG_rl_186 ;
	7'h75 :
		rl_a114_t8 = RG_rl_186 ;
	7'h76 :
		rl_a114_t8 = RG_rl_186 ;
	7'h77 :
		rl_a114_t8 = RG_rl_186 ;
	7'h78 :
		rl_a114_t8 = RG_rl_186 ;
	7'h79 :
		rl_a114_t8 = RG_rl_186 ;
	7'h7a :
		rl_a114_t8 = RG_rl_186 ;
	7'h7b :
		rl_a114_t8 = RG_rl_186 ;
	7'h7c :
		rl_a114_t8 = RG_rl_186 ;
	7'h7d :
		rl_a114_t8 = RG_rl_186 ;
	7'h7e :
		rl_a114_t8 = RG_rl_186 ;
	7'h7f :
		rl_a114_t8 = RG_rl_186 ;
	default :
		rl_a114_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_55 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h01 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h02 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h03 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h04 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h05 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h06 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h07 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h08 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h09 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h0a :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h0b :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h0c :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h0d :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h0e :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h0f :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h10 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h11 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h12 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h13 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h14 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h15 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h16 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h17 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h18 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h19 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h1a :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h1b :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h1c :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h1d :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h1e :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h1f :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h20 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h21 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h22 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h23 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h24 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h25 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h26 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h27 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h28 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h29 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h2a :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h2b :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h2c :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h2d :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h2e :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h2f :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h30 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h31 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h32 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h33 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h34 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h35 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h36 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h37 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h38 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h39 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h3a :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h3b :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h3c :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h3d :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h3e :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h3f :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h40 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h41 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h42 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h43 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h44 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h45 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h46 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h47 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h48 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h49 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h4a :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h4b :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h4c :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h4d :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h4e :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h4f :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h50 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h51 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h52 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h53 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h54 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h55 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h56 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h57 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h58 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h59 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h5a :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h5b :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h5c :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h5d :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h5e :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h5f :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h60 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h61 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h62 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h63 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h64 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h65 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h66 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h67 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h68 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h69 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h6a :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h6b :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h6c :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h6d :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h6e :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h6f :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h70 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h71 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h72 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h73 :
		rl_a115_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h74 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h75 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h76 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h77 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h78 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h79 :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h7a :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h7b :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h7c :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h7d :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h7e :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	7'h7f :
		rl_a115_t8 = RG_quantized_block_rl_55 ;
	default :
		rl_a115_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_187 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a116_t8 = RG_rl_187 ;
	7'h01 :
		rl_a116_t8 = RG_rl_187 ;
	7'h02 :
		rl_a116_t8 = RG_rl_187 ;
	7'h03 :
		rl_a116_t8 = RG_rl_187 ;
	7'h04 :
		rl_a116_t8 = RG_rl_187 ;
	7'h05 :
		rl_a116_t8 = RG_rl_187 ;
	7'h06 :
		rl_a116_t8 = RG_rl_187 ;
	7'h07 :
		rl_a116_t8 = RG_rl_187 ;
	7'h08 :
		rl_a116_t8 = RG_rl_187 ;
	7'h09 :
		rl_a116_t8 = RG_rl_187 ;
	7'h0a :
		rl_a116_t8 = RG_rl_187 ;
	7'h0b :
		rl_a116_t8 = RG_rl_187 ;
	7'h0c :
		rl_a116_t8 = RG_rl_187 ;
	7'h0d :
		rl_a116_t8 = RG_rl_187 ;
	7'h0e :
		rl_a116_t8 = RG_rl_187 ;
	7'h0f :
		rl_a116_t8 = RG_rl_187 ;
	7'h10 :
		rl_a116_t8 = RG_rl_187 ;
	7'h11 :
		rl_a116_t8 = RG_rl_187 ;
	7'h12 :
		rl_a116_t8 = RG_rl_187 ;
	7'h13 :
		rl_a116_t8 = RG_rl_187 ;
	7'h14 :
		rl_a116_t8 = RG_rl_187 ;
	7'h15 :
		rl_a116_t8 = RG_rl_187 ;
	7'h16 :
		rl_a116_t8 = RG_rl_187 ;
	7'h17 :
		rl_a116_t8 = RG_rl_187 ;
	7'h18 :
		rl_a116_t8 = RG_rl_187 ;
	7'h19 :
		rl_a116_t8 = RG_rl_187 ;
	7'h1a :
		rl_a116_t8 = RG_rl_187 ;
	7'h1b :
		rl_a116_t8 = RG_rl_187 ;
	7'h1c :
		rl_a116_t8 = RG_rl_187 ;
	7'h1d :
		rl_a116_t8 = RG_rl_187 ;
	7'h1e :
		rl_a116_t8 = RG_rl_187 ;
	7'h1f :
		rl_a116_t8 = RG_rl_187 ;
	7'h20 :
		rl_a116_t8 = RG_rl_187 ;
	7'h21 :
		rl_a116_t8 = RG_rl_187 ;
	7'h22 :
		rl_a116_t8 = RG_rl_187 ;
	7'h23 :
		rl_a116_t8 = RG_rl_187 ;
	7'h24 :
		rl_a116_t8 = RG_rl_187 ;
	7'h25 :
		rl_a116_t8 = RG_rl_187 ;
	7'h26 :
		rl_a116_t8 = RG_rl_187 ;
	7'h27 :
		rl_a116_t8 = RG_rl_187 ;
	7'h28 :
		rl_a116_t8 = RG_rl_187 ;
	7'h29 :
		rl_a116_t8 = RG_rl_187 ;
	7'h2a :
		rl_a116_t8 = RG_rl_187 ;
	7'h2b :
		rl_a116_t8 = RG_rl_187 ;
	7'h2c :
		rl_a116_t8 = RG_rl_187 ;
	7'h2d :
		rl_a116_t8 = RG_rl_187 ;
	7'h2e :
		rl_a116_t8 = RG_rl_187 ;
	7'h2f :
		rl_a116_t8 = RG_rl_187 ;
	7'h30 :
		rl_a116_t8 = RG_rl_187 ;
	7'h31 :
		rl_a116_t8 = RG_rl_187 ;
	7'h32 :
		rl_a116_t8 = RG_rl_187 ;
	7'h33 :
		rl_a116_t8 = RG_rl_187 ;
	7'h34 :
		rl_a116_t8 = RG_rl_187 ;
	7'h35 :
		rl_a116_t8 = RG_rl_187 ;
	7'h36 :
		rl_a116_t8 = RG_rl_187 ;
	7'h37 :
		rl_a116_t8 = RG_rl_187 ;
	7'h38 :
		rl_a116_t8 = RG_rl_187 ;
	7'h39 :
		rl_a116_t8 = RG_rl_187 ;
	7'h3a :
		rl_a116_t8 = RG_rl_187 ;
	7'h3b :
		rl_a116_t8 = RG_rl_187 ;
	7'h3c :
		rl_a116_t8 = RG_rl_187 ;
	7'h3d :
		rl_a116_t8 = RG_rl_187 ;
	7'h3e :
		rl_a116_t8 = RG_rl_187 ;
	7'h3f :
		rl_a116_t8 = RG_rl_187 ;
	7'h40 :
		rl_a116_t8 = RG_rl_187 ;
	7'h41 :
		rl_a116_t8 = RG_rl_187 ;
	7'h42 :
		rl_a116_t8 = RG_rl_187 ;
	7'h43 :
		rl_a116_t8 = RG_rl_187 ;
	7'h44 :
		rl_a116_t8 = RG_rl_187 ;
	7'h45 :
		rl_a116_t8 = RG_rl_187 ;
	7'h46 :
		rl_a116_t8 = RG_rl_187 ;
	7'h47 :
		rl_a116_t8 = RG_rl_187 ;
	7'h48 :
		rl_a116_t8 = RG_rl_187 ;
	7'h49 :
		rl_a116_t8 = RG_rl_187 ;
	7'h4a :
		rl_a116_t8 = RG_rl_187 ;
	7'h4b :
		rl_a116_t8 = RG_rl_187 ;
	7'h4c :
		rl_a116_t8 = RG_rl_187 ;
	7'h4d :
		rl_a116_t8 = RG_rl_187 ;
	7'h4e :
		rl_a116_t8 = RG_rl_187 ;
	7'h4f :
		rl_a116_t8 = RG_rl_187 ;
	7'h50 :
		rl_a116_t8 = RG_rl_187 ;
	7'h51 :
		rl_a116_t8 = RG_rl_187 ;
	7'h52 :
		rl_a116_t8 = RG_rl_187 ;
	7'h53 :
		rl_a116_t8 = RG_rl_187 ;
	7'h54 :
		rl_a116_t8 = RG_rl_187 ;
	7'h55 :
		rl_a116_t8 = RG_rl_187 ;
	7'h56 :
		rl_a116_t8 = RG_rl_187 ;
	7'h57 :
		rl_a116_t8 = RG_rl_187 ;
	7'h58 :
		rl_a116_t8 = RG_rl_187 ;
	7'h59 :
		rl_a116_t8 = RG_rl_187 ;
	7'h5a :
		rl_a116_t8 = RG_rl_187 ;
	7'h5b :
		rl_a116_t8 = RG_rl_187 ;
	7'h5c :
		rl_a116_t8 = RG_rl_187 ;
	7'h5d :
		rl_a116_t8 = RG_rl_187 ;
	7'h5e :
		rl_a116_t8 = RG_rl_187 ;
	7'h5f :
		rl_a116_t8 = RG_rl_187 ;
	7'h60 :
		rl_a116_t8 = RG_rl_187 ;
	7'h61 :
		rl_a116_t8 = RG_rl_187 ;
	7'h62 :
		rl_a116_t8 = RG_rl_187 ;
	7'h63 :
		rl_a116_t8 = RG_rl_187 ;
	7'h64 :
		rl_a116_t8 = RG_rl_187 ;
	7'h65 :
		rl_a116_t8 = RG_rl_187 ;
	7'h66 :
		rl_a116_t8 = RG_rl_187 ;
	7'h67 :
		rl_a116_t8 = RG_rl_187 ;
	7'h68 :
		rl_a116_t8 = RG_rl_187 ;
	7'h69 :
		rl_a116_t8 = RG_rl_187 ;
	7'h6a :
		rl_a116_t8 = RG_rl_187 ;
	7'h6b :
		rl_a116_t8 = RG_rl_187 ;
	7'h6c :
		rl_a116_t8 = RG_rl_187 ;
	7'h6d :
		rl_a116_t8 = RG_rl_187 ;
	7'h6e :
		rl_a116_t8 = RG_rl_187 ;
	7'h6f :
		rl_a116_t8 = RG_rl_187 ;
	7'h70 :
		rl_a116_t8 = RG_rl_187 ;
	7'h71 :
		rl_a116_t8 = RG_rl_187 ;
	7'h72 :
		rl_a116_t8 = RG_rl_187 ;
	7'h73 :
		rl_a116_t8 = RG_rl_187 ;
	7'h74 :
		rl_a116_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h75 :
		rl_a116_t8 = RG_rl_187 ;
	7'h76 :
		rl_a116_t8 = RG_rl_187 ;
	7'h77 :
		rl_a116_t8 = RG_rl_187 ;
	7'h78 :
		rl_a116_t8 = RG_rl_187 ;
	7'h79 :
		rl_a116_t8 = RG_rl_187 ;
	7'h7a :
		rl_a116_t8 = RG_rl_187 ;
	7'h7b :
		rl_a116_t8 = RG_rl_187 ;
	7'h7c :
		rl_a116_t8 = RG_rl_187 ;
	7'h7d :
		rl_a116_t8 = RG_rl_187 ;
	7'h7e :
		rl_a116_t8 = RG_rl_187 ;
	7'h7f :
		rl_a116_t8 = RG_rl_187 ;
	default :
		rl_a116_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_56 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h01 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h02 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h03 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h04 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h05 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h06 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h07 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h08 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h09 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h0a :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h0b :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h0c :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h0d :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h0e :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h0f :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h10 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h11 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h12 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h13 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h14 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h15 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h16 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h17 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h18 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h19 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h1a :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h1b :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h1c :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h1d :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h1e :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h1f :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h20 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h21 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h22 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h23 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h24 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h25 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h26 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h27 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h28 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h29 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h2a :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h2b :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h2c :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h2d :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h2e :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h2f :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h30 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h31 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h32 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h33 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h34 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h35 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h36 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h37 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h38 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h39 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h3a :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h3b :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h3c :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h3d :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h3e :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h3f :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h40 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h41 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h42 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h43 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h44 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h45 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h46 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h47 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h48 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h49 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h4a :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h4b :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h4c :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h4d :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h4e :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h4f :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h50 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h51 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h52 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h53 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h54 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h55 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h56 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h57 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h58 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h59 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h5a :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h5b :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h5c :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h5d :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h5e :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h5f :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h60 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h61 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h62 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h63 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h64 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h65 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h66 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h67 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h68 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h69 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h6a :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h6b :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h6c :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h6d :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h6e :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h6f :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h70 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h71 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h72 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h73 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h74 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h75 :
		rl_a117_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h76 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h77 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h78 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h79 :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h7a :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h7b :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h7c :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h7d :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h7e :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	7'h7f :
		rl_a117_t8 = RG_quantized_block_rl_56 ;
	default :
		rl_a117_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_188 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a118_t8 = RG_rl_188 ;
	7'h01 :
		rl_a118_t8 = RG_rl_188 ;
	7'h02 :
		rl_a118_t8 = RG_rl_188 ;
	7'h03 :
		rl_a118_t8 = RG_rl_188 ;
	7'h04 :
		rl_a118_t8 = RG_rl_188 ;
	7'h05 :
		rl_a118_t8 = RG_rl_188 ;
	7'h06 :
		rl_a118_t8 = RG_rl_188 ;
	7'h07 :
		rl_a118_t8 = RG_rl_188 ;
	7'h08 :
		rl_a118_t8 = RG_rl_188 ;
	7'h09 :
		rl_a118_t8 = RG_rl_188 ;
	7'h0a :
		rl_a118_t8 = RG_rl_188 ;
	7'h0b :
		rl_a118_t8 = RG_rl_188 ;
	7'h0c :
		rl_a118_t8 = RG_rl_188 ;
	7'h0d :
		rl_a118_t8 = RG_rl_188 ;
	7'h0e :
		rl_a118_t8 = RG_rl_188 ;
	7'h0f :
		rl_a118_t8 = RG_rl_188 ;
	7'h10 :
		rl_a118_t8 = RG_rl_188 ;
	7'h11 :
		rl_a118_t8 = RG_rl_188 ;
	7'h12 :
		rl_a118_t8 = RG_rl_188 ;
	7'h13 :
		rl_a118_t8 = RG_rl_188 ;
	7'h14 :
		rl_a118_t8 = RG_rl_188 ;
	7'h15 :
		rl_a118_t8 = RG_rl_188 ;
	7'h16 :
		rl_a118_t8 = RG_rl_188 ;
	7'h17 :
		rl_a118_t8 = RG_rl_188 ;
	7'h18 :
		rl_a118_t8 = RG_rl_188 ;
	7'h19 :
		rl_a118_t8 = RG_rl_188 ;
	7'h1a :
		rl_a118_t8 = RG_rl_188 ;
	7'h1b :
		rl_a118_t8 = RG_rl_188 ;
	7'h1c :
		rl_a118_t8 = RG_rl_188 ;
	7'h1d :
		rl_a118_t8 = RG_rl_188 ;
	7'h1e :
		rl_a118_t8 = RG_rl_188 ;
	7'h1f :
		rl_a118_t8 = RG_rl_188 ;
	7'h20 :
		rl_a118_t8 = RG_rl_188 ;
	7'h21 :
		rl_a118_t8 = RG_rl_188 ;
	7'h22 :
		rl_a118_t8 = RG_rl_188 ;
	7'h23 :
		rl_a118_t8 = RG_rl_188 ;
	7'h24 :
		rl_a118_t8 = RG_rl_188 ;
	7'h25 :
		rl_a118_t8 = RG_rl_188 ;
	7'h26 :
		rl_a118_t8 = RG_rl_188 ;
	7'h27 :
		rl_a118_t8 = RG_rl_188 ;
	7'h28 :
		rl_a118_t8 = RG_rl_188 ;
	7'h29 :
		rl_a118_t8 = RG_rl_188 ;
	7'h2a :
		rl_a118_t8 = RG_rl_188 ;
	7'h2b :
		rl_a118_t8 = RG_rl_188 ;
	7'h2c :
		rl_a118_t8 = RG_rl_188 ;
	7'h2d :
		rl_a118_t8 = RG_rl_188 ;
	7'h2e :
		rl_a118_t8 = RG_rl_188 ;
	7'h2f :
		rl_a118_t8 = RG_rl_188 ;
	7'h30 :
		rl_a118_t8 = RG_rl_188 ;
	7'h31 :
		rl_a118_t8 = RG_rl_188 ;
	7'h32 :
		rl_a118_t8 = RG_rl_188 ;
	7'h33 :
		rl_a118_t8 = RG_rl_188 ;
	7'h34 :
		rl_a118_t8 = RG_rl_188 ;
	7'h35 :
		rl_a118_t8 = RG_rl_188 ;
	7'h36 :
		rl_a118_t8 = RG_rl_188 ;
	7'h37 :
		rl_a118_t8 = RG_rl_188 ;
	7'h38 :
		rl_a118_t8 = RG_rl_188 ;
	7'h39 :
		rl_a118_t8 = RG_rl_188 ;
	7'h3a :
		rl_a118_t8 = RG_rl_188 ;
	7'h3b :
		rl_a118_t8 = RG_rl_188 ;
	7'h3c :
		rl_a118_t8 = RG_rl_188 ;
	7'h3d :
		rl_a118_t8 = RG_rl_188 ;
	7'h3e :
		rl_a118_t8 = RG_rl_188 ;
	7'h3f :
		rl_a118_t8 = RG_rl_188 ;
	7'h40 :
		rl_a118_t8 = RG_rl_188 ;
	7'h41 :
		rl_a118_t8 = RG_rl_188 ;
	7'h42 :
		rl_a118_t8 = RG_rl_188 ;
	7'h43 :
		rl_a118_t8 = RG_rl_188 ;
	7'h44 :
		rl_a118_t8 = RG_rl_188 ;
	7'h45 :
		rl_a118_t8 = RG_rl_188 ;
	7'h46 :
		rl_a118_t8 = RG_rl_188 ;
	7'h47 :
		rl_a118_t8 = RG_rl_188 ;
	7'h48 :
		rl_a118_t8 = RG_rl_188 ;
	7'h49 :
		rl_a118_t8 = RG_rl_188 ;
	7'h4a :
		rl_a118_t8 = RG_rl_188 ;
	7'h4b :
		rl_a118_t8 = RG_rl_188 ;
	7'h4c :
		rl_a118_t8 = RG_rl_188 ;
	7'h4d :
		rl_a118_t8 = RG_rl_188 ;
	7'h4e :
		rl_a118_t8 = RG_rl_188 ;
	7'h4f :
		rl_a118_t8 = RG_rl_188 ;
	7'h50 :
		rl_a118_t8 = RG_rl_188 ;
	7'h51 :
		rl_a118_t8 = RG_rl_188 ;
	7'h52 :
		rl_a118_t8 = RG_rl_188 ;
	7'h53 :
		rl_a118_t8 = RG_rl_188 ;
	7'h54 :
		rl_a118_t8 = RG_rl_188 ;
	7'h55 :
		rl_a118_t8 = RG_rl_188 ;
	7'h56 :
		rl_a118_t8 = RG_rl_188 ;
	7'h57 :
		rl_a118_t8 = RG_rl_188 ;
	7'h58 :
		rl_a118_t8 = RG_rl_188 ;
	7'h59 :
		rl_a118_t8 = RG_rl_188 ;
	7'h5a :
		rl_a118_t8 = RG_rl_188 ;
	7'h5b :
		rl_a118_t8 = RG_rl_188 ;
	7'h5c :
		rl_a118_t8 = RG_rl_188 ;
	7'h5d :
		rl_a118_t8 = RG_rl_188 ;
	7'h5e :
		rl_a118_t8 = RG_rl_188 ;
	7'h5f :
		rl_a118_t8 = RG_rl_188 ;
	7'h60 :
		rl_a118_t8 = RG_rl_188 ;
	7'h61 :
		rl_a118_t8 = RG_rl_188 ;
	7'h62 :
		rl_a118_t8 = RG_rl_188 ;
	7'h63 :
		rl_a118_t8 = RG_rl_188 ;
	7'h64 :
		rl_a118_t8 = RG_rl_188 ;
	7'h65 :
		rl_a118_t8 = RG_rl_188 ;
	7'h66 :
		rl_a118_t8 = RG_rl_188 ;
	7'h67 :
		rl_a118_t8 = RG_rl_188 ;
	7'h68 :
		rl_a118_t8 = RG_rl_188 ;
	7'h69 :
		rl_a118_t8 = RG_rl_188 ;
	7'h6a :
		rl_a118_t8 = RG_rl_188 ;
	7'h6b :
		rl_a118_t8 = RG_rl_188 ;
	7'h6c :
		rl_a118_t8 = RG_rl_188 ;
	7'h6d :
		rl_a118_t8 = RG_rl_188 ;
	7'h6e :
		rl_a118_t8 = RG_rl_188 ;
	7'h6f :
		rl_a118_t8 = RG_rl_188 ;
	7'h70 :
		rl_a118_t8 = RG_rl_188 ;
	7'h71 :
		rl_a118_t8 = RG_rl_188 ;
	7'h72 :
		rl_a118_t8 = RG_rl_188 ;
	7'h73 :
		rl_a118_t8 = RG_rl_188 ;
	7'h74 :
		rl_a118_t8 = RG_rl_188 ;
	7'h75 :
		rl_a118_t8 = RG_rl_188 ;
	7'h76 :
		rl_a118_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h77 :
		rl_a118_t8 = RG_rl_188 ;
	7'h78 :
		rl_a118_t8 = RG_rl_188 ;
	7'h79 :
		rl_a118_t8 = RG_rl_188 ;
	7'h7a :
		rl_a118_t8 = RG_rl_188 ;
	7'h7b :
		rl_a118_t8 = RG_rl_188 ;
	7'h7c :
		rl_a118_t8 = RG_rl_188 ;
	7'h7d :
		rl_a118_t8 = RG_rl_188 ;
	7'h7e :
		rl_a118_t8 = RG_rl_188 ;
	7'h7f :
		rl_a118_t8 = RG_rl_188 ;
	default :
		rl_a118_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_57 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h01 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h02 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h03 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h04 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h05 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h06 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h07 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h08 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h09 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h0a :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h0b :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h0c :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h0d :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h0e :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h0f :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h10 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h11 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h12 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h13 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h14 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h15 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h16 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h17 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h18 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h19 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h1a :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h1b :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h1c :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h1d :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h1e :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h1f :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h20 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h21 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h22 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h23 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h24 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h25 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h26 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h27 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h28 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h29 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h2a :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h2b :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h2c :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h2d :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h2e :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h2f :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h30 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h31 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h32 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h33 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h34 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h35 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h36 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h37 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h38 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h39 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h3a :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h3b :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h3c :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h3d :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h3e :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h3f :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h40 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h41 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h42 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h43 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h44 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h45 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h46 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h47 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h48 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h49 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h4a :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h4b :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h4c :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h4d :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h4e :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h4f :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h50 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h51 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h52 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h53 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h54 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h55 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h56 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h57 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h58 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h59 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h5a :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h5b :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h5c :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h5d :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h5e :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h5f :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h60 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h61 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h62 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h63 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h64 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h65 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h66 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h67 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h68 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h69 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h6a :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h6b :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h6c :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h6d :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h6e :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h6f :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h70 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h71 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h72 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h73 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h74 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h75 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h76 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h77 :
		rl_a119_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h78 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h79 :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h7a :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h7b :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h7c :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h7d :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h7e :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	7'h7f :
		rl_a119_t8 = RG_quantized_block_rl_57 ;
	default :
		rl_a119_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_189 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a120_t8 = RG_rl_189 ;
	7'h01 :
		rl_a120_t8 = RG_rl_189 ;
	7'h02 :
		rl_a120_t8 = RG_rl_189 ;
	7'h03 :
		rl_a120_t8 = RG_rl_189 ;
	7'h04 :
		rl_a120_t8 = RG_rl_189 ;
	7'h05 :
		rl_a120_t8 = RG_rl_189 ;
	7'h06 :
		rl_a120_t8 = RG_rl_189 ;
	7'h07 :
		rl_a120_t8 = RG_rl_189 ;
	7'h08 :
		rl_a120_t8 = RG_rl_189 ;
	7'h09 :
		rl_a120_t8 = RG_rl_189 ;
	7'h0a :
		rl_a120_t8 = RG_rl_189 ;
	7'h0b :
		rl_a120_t8 = RG_rl_189 ;
	7'h0c :
		rl_a120_t8 = RG_rl_189 ;
	7'h0d :
		rl_a120_t8 = RG_rl_189 ;
	7'h0e :
		rl_a120_t8 = RG_rl_189 ;
	7'h0f :
		rl_a120_t8 = RG_rl_189 ;
	7'h10 :
		rl_a120_t8 = RG_rl_189 ;
	7'h11 :
		rl_a120_t8 = RG_rl_189 ;
	7'h12 :
		rl_a120_t8 = RG_rl_189 ;
	7'h13 :
		rl_a120_t8 = RG_rl_189 ;
	7'h14 :
		rl_a120_t8 = RG_rl_189 ;
	7'h15 :
		rl_a120_t8 = RG_rl_189 ;
	7'h16 :
		rl_a120_t8 = RG_rl_189 ;
	7'h17 :
		rl_a120_t8 = RG_rl_189 ;
	7'h18 :
		rl_a120_t8 = RG_rl_189 ;
	7'h19 :
		rl_a120_t8 = RG_rl_189 ;
	7'h1a :
		rl_a120_t8 = RG_rl_189 ;
	7'h1b :
		rl_a120_t8 = RG_rl_189 ;
	7'h1c :
		rl_a120_t8 = RG_rl_189 ;
	7'h1d :
		rl_a120_t8 = RG_rl_189 ;
	7'h1e :
		rl_a120_t8 = RG_rl_189 ;
	7'h1f :
		rl_a120_t8 = RG_rl_189 ;
	7'h20 :
		rl_a120_t8 = RG_rl_189 ;
	7'h21 :
		rl_a120_t8 = RG_rl_189 ;
	7'h22 :
		rl_a120_t8 = RG_rl_189 ;
	7'h23 :
		rl_a120_t8 = RG_rl_189 ;
	7'h24 :
		rl_a120_t8 = RG_rl_189 ;
	7'h25 :
		rl_a120_t8 = RG_rl_189 ;
	7'h26 :
		rl_a120_t8 = RG_rl_189 ;
	7'h27 :
		rl_a120_t8 = RG_rl_189 ;
	7'h28 :
		rl_a120_t8 = RG_rl_189 ;
	7'h29 :
		rl_a120_t8 = RG_rl_189 ;
	7'h2a :
		rl_a120_t8 = RG_rl_189 ;
	7'h2b :
		rl_a120_t8 = RG_rl_189 ;
	7'h2c :
		rl_a120_t8 = RG_rl_189 ;
	7'h2d :
		rl_a120_t8 = RG_rl_189 ;
	7'h2e :
		rl_a120_t8 = RG_rl_189 ;
	7'h2f :
		rl_a120_t8 = RG_rl_189 ;
	7'h30 :
		rl_a120_t8 = RG_rl_189 ;
	7'h31 :
		rl_a120_t8 = RG_rl_189 ;
	7'h32 :
		rl_a120_t8 = RG_rl_189 ;
	7'h33 :
		rl_a120_t8 = RG_rl_189 ;
	7'h34 :
		rl_a120_t8 = RG_rl_189 ;
	7'h35 :
		rl_a120_t8 = RG_rl_189 ;
	7'h36 :
		rl_a120_t8 = RG_rl_189 ;
	7'h37 :
		rl_a120_t8 = RG_rl_189 ;
	7'h38 :
		rl_a120_t8 = RG_rl_189 ;
	7'h39 :
		rl_a120_t8 = RG_rl_189 ;
	7'h3a :
		rl_a120_t8 = RG_rl_189 ;
	7'h3b :
		rl_a120_t8 = RG_rl_189 ;
	7'h3c :
		rl_a120_t8 = RG_rl_189 ;
	7'h3d :
		rl_a120_t8 = RG_rl_189 ;
	7'h3e :
		rl_a120_t8 = RG_rl_189 ;
	7'h3f :
		rl_a120_t8 = RG_rl_189 ;
	7'h40 :
		rl_a120_t8 = RG_rl_189 ;
	7'h41 :
		rl_a120_t8 = RG_rl_189 ;
	7'h42 :
		rl_a120_t8 = RG_rl_189 ;
	7'h43 :
		rl_a120_t8 = RG_rl_189 ;
	7'h44 :
		rl_a120_t8 = RG_rl_189 ;
	7'h45 :
		rl_a120_t8 = RG_rl_189 ;
	7'h46 :
		rl_a120_t8 = RG_rl_189 ;
	7'h47 :
		rl_a120_t8 = RG_rl_189 ;
	7'h48 :
		rl_a120_t8 = RG_rl_189 ;
	7'h49 :
		rl_a120_t8 = RG_rl_189 ;
	7'h4a :
		rl_a120_t8 = RG_rl_189 ;
	7'h4b :
		rl_a120_t8 = RG_rl_189 ;
	7'h4c :
		rl_a120_t8 = RG_rl_189 ;
	7'h4d :
		rl_a120_t8 = RG_rl_189 ;
	7'h4e :
		rl_a120_t8 = RG_rl_189 ;
	7'h4f :
		rl_a120_t8 = RG_rl_189 ;
	7'h50 :
		rl_a120_t8 = RG_rl_189 ;
	7'h51 :
		rl_a120_t8 = RG_rl_189 ;
	7'h52 :
		rl_a120_t8 = RG_rl_189 ;
	7'h53 :
		rl_a120_t8 = RG_rl_189 ;
	7'h54 :
		rl_a120_t8 = RG_rl_189 ;
	7'h55 :
		rl_a120_t8 = RG_rl_189 ;
	7'h56 :
		rl_a120_t8 = RG_rl_189 ;
	7'h57 :
		rl_a120_t8 = RG_rl_189 ;
	7'h58 :
		rl_a120_t8 = RG_rl_189 ;
	7'h59 :
		rl_a120_t8 = RG_rl_189 ;
	7'h5a :
		rl_a120_t8 = RG_rl_189 ;
	7'h5b :
		rl_a120_t8 = RG_rl_189 ;
	7'h5c :
		rl_a120_t8 = RG_rl_189 ;
	7'h5d :
		rl_a120_t8 = RG_rl_189 ;
	7'h5e :
		rl_a120_t8 = RG_rl_189 ;
	7'h5f :
		rl_a120_t8 = RG_rl_189 ;
	7'h60 :
		rl_a120_t8 = RG_rl_189 ;
	7'h61 :
		rl_a120_t8 = RG_rl_189 ;
	7'h62 :
		rl_a120_t8 = RG_rl_189 ;
	7'h63 :
		rl_a120_t8 = RG_rl_189 ;
	7'h64 :
		rl_a120_t8 = RG_rl_189 ;
	7'h65 :
		rl_a120_t8 = RG_rl_189 ;
	7'h66 :
		rl_a120_t8 = RG_rl_189 ;
	7'h67 :
		rl_a120_t8 = RG_rl_189 ;
	7'h68 :
		rl_a120_t8 = RG_rl_189 ;
	7'h69 :
		rl_a120_t8 = RG_rl_189 ;
	7'h6a :
		rl_a120_t8 = RG_rl_189 ;
	7'h6b :
		rl_a120_t8 = RG_rl_189 ;
	7'h6c :
		rl_a120_t8 = RG_rl_189 ;
	7'h6d :
		rl_a120_t8 = RG_rl_189 ;
	7'h6e :
		rl_a120_t8 = RG_rl_189 ;
	7'h6f :
		rl_a120_t8 = RG_rl_189 ;
	7'h70 :
		rl_a120_t8 = RG_rl_189 ;
	7'h71 :
		rl_a120_t8 = RG_rl_189 ;
	7'h72 :
		rl_a120_t8 = RG_rl_189 ;
	7'h73 :
		rl_a120_t8 = RG_rl_189 ;
	7'h74 :
		rl_a120_t8 = RG_rl_189 ;
	7'h75 :
		rl_a120_t8 = RG_rl_189 ;
	7'h76 :
		rl_a120_t8 = RG_rl_189 ;
	7'h77 :
		rl_a120_t8 = RG_rl_189 ;
	7'h78 :
		rl_a120_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h79 :
		rl_a120_t8 = RG_rl_189 ;
	7'h7a :
		rl_a120_t8 = RG_rl_189 ;
	7'h7b :
		rl_a120_t8 = RG_rl_189 ;
	7'h7c :
		rl_a120_t8 = RG_rl_189 ;
	7'h7d :
		rl_a120_t8 = RG_rl_189 ;
	7'h7e :
		rl_a120_t8 = RG_rl_189 ;
	7'h7f :
		rl_a120_t8 = RG_rl_189 ;
	default :
		rl_a120_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_58 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h01 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h02 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h03 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h04 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h05 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h06 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h07 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h08 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h09 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h0a :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h0b :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h0c :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h0d :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h0e :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h0f :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h10 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h11 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h12 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h13 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h14 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h15 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h16 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h17 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h18 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h19 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h1a :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h1b :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h1c :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h1d :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h1e :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h1f :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h20 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h21 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h22 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h23 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h24 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h25 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h26 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h27 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h28 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h29 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h2a :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h2b :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h2c :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h2d :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h2e :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h2f :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h30 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h31 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h32 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h33 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h34 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h35 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h36 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h37 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h38 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h39 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h3a :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h3b :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h3c :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h3d :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h3e :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h3f :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h40 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h41 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h42 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h43 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h44 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h45 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h46 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h47 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h48 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h49 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h4a :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h4b :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h4c :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h4d :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h4e :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h4f :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h50 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h51 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h52 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h53 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h54 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h55 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h56 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h57 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h58 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h59 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h5a :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h5b :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h5c :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h5d :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h5e :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h5f :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h60 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h61 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h62 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h63 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h64 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h65 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h66 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h67 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h68 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h69 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h6a :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h6b :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h6c :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h6d :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h6e :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h6f :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h70 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h71 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h72 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h73 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h74 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h75 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h76 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h77 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h78 :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h79 :
		rl_a121_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h7a :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h7b :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h7c :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h7d :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h7e :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	7'h7f :
		rl_a121_t8 = RG_quantized_block_rl_58 ;
	default :
		rl_a121_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_190 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a122_t8 = RG_rl_190 ;
	7'h01 :
		rl_a122_t8 = RG_rl_190 ;
	7'h02 :
		rl_a122_t8 = RG_rl_190 ;
	7'h03 :
		rl_a122_t8 = RG_rl_190 ;
	7'h04 :
		rl_a122_t8 = RG_rl_190 ;
	7'h05 :
		rl_a122_t8 = RG_rl_190 ;
	7'h06 :
		rl_a122_t8 = RG_rl_190 ;
	7'h07 :
		rl_a122_t8 = RG_rl_190 ;
	7'h08 :
		rl_a122_t8 = RG_rl_190 ;
	7'h09 :
		rl_a122_t8 = RG_rl_190 ;
	7'h0a :
		rl_a122_t8 = RG_rl_190 ;
	7'h0b :
		rl_a122_t8 = RG_rl_190 ;
	7'h0c :
		rl_a122_t8 = RG_rl_190 ;
	7'h0d :
		rl_a122_t8 = RG_rl_190 ;
	7'h0e :
		rl_a122_t8 = RG_rl_190 ;
	7'h0f :
		rl_a122_t8 = RG_rl_190 ;
	7'h10 :
		rl_a122_t8 = RG_rl_190 ;
	7'h11 :
		rl_a122_t8 = RG_rl_190 ;
	7'h12 :
		rl_a122_t8 = RG_rl_190 ;
	7'h13 :
		rl_a122_t8 = RG_rl_190 ;
	7'h14 :
		rl_a122_t8 = RG_rl_190 ;
	7'h15 :
		rl_a122_t8 = RG_rl_190 ;
	7'h16 :
		rl_a122_t8 = RG_rl_190 ;
	7'h17 :
		rl_a122_t8 = RG_rl_190 ;
	7'h18 :
		rl_a122_t8 = RG_rl_190 ;
	7'h19 :
		rl_a122_t8 = RG_rl_190 ;
	7'h1a :
		rl_a122_t8 = RG_rl_190 ;
	7'h1b :
		rl_a122_t8 = RG_rl_190 ;
	7'h1c :
		rl_a122_t8 = RG_rl_190 ;
	7'h1d :
		rl_a122_t8 = RG_rl_190 ;
	7'h1e :
		rl_a122_t8 = RG_rl_190 ;
	7'h1f :
		rl_a122_t8 = RG_rl_190 ;
	7'h20 :
		rl_a122_t8 = RG_rl_190 ;
	7'h21 :
		rl_a122_t8 = RG_rl_190 ;
	7'h22 :
		rl_a122_t8 = RG_rl_190 ;
	7'h23 :
		rl_a122_t8 = RG_rl_190 ;
	7'h24 :
		rl_a122_t8 = RG_rl_190 ;
	7'h25 :
		rl_a122_t8 = RG_rl_190 ;
	7'h26 :
		rl_a122_t8 = RG_rl_190 ;
	7'h27 :
		rl_a122_t8 = RG_rl_190 ;
	7'h28 :
		rl_a122_t8 = RG_rl_190 ;
	7'h29 :
		rl_a122_t8 = RG_rl_190 ;
	7'h2a :
		rl_a122_t8 = RG_rl_190 ;
	7'h2b :
		rl_a122_t8 = RG_rl_190 ;
	7'h2c :
		rl_a122_t8 = RG_rl_190 ;
	7'h2d :
		rl_a122_t8 = RG_rl_190 ;
	7'h2e :
		rl_a122_t8 = RG_rl_190 ;
	7'h2f :
		rl_a122_t8 = RG_rl_190 ;
	7'h30 :
		rl_a122_t8 = RG_rl_190 ;
	7'h31 :
		rl_a122_t8 = RG_rl_190 ;
	7'h32 :
		rl_a122_t8 = RG_rl_190 ;
	7'h33 :
		rl_a122_t8 = RG_rl_190 ;
	7'h34 :
		rl_a122_t8 = RG_rl_190 ;
	7'h35 :
		rl_a122_t8 = RG_rl_190 ;
	7'h36 :
		rl_a122_t8 = RG_rl_190 ;
	7'h37 :
		rl_a122_t8 = RG_rl_190 ;
	7'h38 :
		rl_a122_t8 = RG_rl_190 ;
	7'h39 :
		rl_a122_t8 = RG_rl_190 ;
	7'h3a :
		rl_a122_t8 = RG_rl_190 ;
	7'h3b :
		rl_a122_t8 = RG_rl_190 ;
	7'h3c :
		rl_a122_t8 = RG_rl_190 ;
	7'h3d :
		rl_a122_t8 = RG_rl_190 ;
	7'h3e :
		rl_a122_t8 = RG_rl_190 ;
	7'h3f :
		rl_a122_t8 = RG_rl_190 ;
	7'h40 :
		rl_a122_t8 = RG_rl_190 ;
	7'h41 :
		rl_a122_t8 = RG_rl_190 ;
	7'h42 :
		rl_a122_t8 = RG_rl_190 ;
	7'h43 :
		rl_a122_t8 = RG_rl_190 ;
	7'h44 :
		rl_a122_t8 = RG_rl_190 ;
	7'h45 :
		rl_a122_t8 = RG_rl_190 ;
	7'h46 :
		rl_a122_t8 = RG_rl_190 ;
	7'h47 :
		rl_a122_t8 = RG_rl_190 ;
	7'h48 :
		rl_a122_t8 = RG_rl_190 ;
	7'h49 :
		rl_a122_t8 = RG_rl_190 ;
	7'h4a :
		rl_a122_t8 = RG_rl_190 ;
	7'h4b :
		rl_a122_t8 = RG_rl_190 ;
	7'h4c :
		rl_a122_t8 = RG_rl_190 ;
	7'h4d :
		rl_a122_t8 = RG_rl_190 ;
	7'h4e :
		rl_a122_t8 = RG_rl_190 ;
	7'h4f :
		rl_a122_t8 = RG_rl_190 ;
	7'h50 :
		rl_a122_t8 = RG_rl_190 ;
	7'h51 :
		rl_a122_t8 = RG_rl_190 ;
	7'h52 :
		rl_a122_t8 = RG_rl_190 ;
	7'h53 :
		rl_a122_t8 = RG_rl_190 ;
	7'h54 :
		rl_a122_t8 = RG_rl_190 ;
	7'h55 :
		rl_a122_t8 = RG_rl_190 ;
	7'h56 :
		rl_a122_t8 = RG_rl_190 ;
	7'h57 :
		rl_a122_t8 = RG_rl_190 ;
	7'h58 :
		rl_a122_t8 = RG_rl_190 ;
	7'h59 :
		rl_a122_t8 = RG_rl_190 ;
	7'h5a :
		rl_a122_t8 = RG_rl_190 ;
	7'h5b :
		rl_a122_t8 = RG_rl_190 ;
	7'h5c :
		rl_a122_t8 = RG_rl_190 ;
	7'h5d :
		rl_a122_t8 = RG_rl_190 ;
	7'h5e :
		rl_a122_t8 = RG_rl_190 ;
	7'h5f :
		rl_a122_t8 = RG_rl_190 ;
	7'h60 :
		rl_a122_t8 = RG_rl_190 ;
	7'h61 :
		rl_a122_t8 = RG_rl_190 ;
	7'h62 :
		rl_a122_t8 = RG_rl_190 ;
	7'h63 :
		rl_a122_t8 = RG_rl_190 ;
	7'h64 :
		rl_a122_t8 = RG_rl_190 ;
	7'h65 :
		rl_a122_t8 = RG_rl_190 ;
	7'h66 :
		rl_a122_t8 = RG_rl_190 ;
	7'h67 :
		rl_a122_t8 = RG_rl_190 ;
	7'h68 :
		rl_a122_t8 = RG_rl_190 ;
	7'h69 :
		rl_a122_t8 = RG_rl_190 ;
	7'h6a :
		rl_a122_t8 = RG_rl_190 ;
	7'h6b :
		rl_a122_t8 = RG_rl_190 ;
	7'h6c :
		rl_a122_t8 = RG_rl_190 ;
	7'h6d :
		rl_a122_t8 = RG_rl_190 ;
	7'h6e :
		rl_a122_t8 = RG_rl_190 ;
	7'h6f :
		rl_a122_t8 = RG_rl_190 ;
	7'h70 :
		rl_a122_t8 = RG_rl_190 ;
	7'h71 :
		rl_a122_t8 = RG_rl_190 ;
	7'h72 :
		rl_a122_t8 = RG_rl_190 ;
	7'h73 :
		rl_a122_t8 = RG_rl_190 ;
	7'h74 :
		rl_a122_t8 = RG_rl_190 ;
	7'h75 :
		rl_a122_t8 = RG_rl_190 ;
	7'h76 :
		rl_a122_t8 = RG_rl_190 ;
	7'h77 :
		rl_a122_t8 = RG_rl_190 ;
	7'h78 :
		rl_a122_t8 = RG_rl_190 ;
	7'h79 :
		rl_a122_t8 = RG_rl_190 ;
	7'h7a :
		rl_a122_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h7b :
		rl_a122_t8 = RG_rl_190 ;
	7'h7c :
		rl_a122_t8 = RG_rl_190 ;
	7'h7d :
		rl_a122_t8 = RG_rl_190 ;
	7'h7e :
		rl_a122_t8 = RG_rl_190 ;
	7'h7f :
		rl_a122_t8 = RG_rl_190 ;
	default :
		rl_a122_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_59 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h01 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h02 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h03 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h04 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h05 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h06 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h07 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h08 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h09 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h0a :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h0b :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h0c :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h0d :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h0e :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h0f :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h10 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h11 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h12 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h13 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h14 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h15 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h16 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h17 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h18 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h19 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h1a :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h1b :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h1c :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h1d :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h1e :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h1f :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h20 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h21 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h22 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h23 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h24 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h25 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h26 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h27 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h28 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h29 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h2a :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h2b :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h2c :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h2d :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h2e :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h2f :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h30 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h31 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h32 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h33 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h34 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h35 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h36 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h37 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h38 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h39 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h3a :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h3b :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h3c :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h3d :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h3e :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h3f :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h40 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h41 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h42 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h43 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h44 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h45 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h46 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h47 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h48 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h49 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h4a :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h4b :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h4c :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h4d :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h4e :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h4f :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h50 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h51 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h52 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h53 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h54 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h55 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h56 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h57 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h58 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h59 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h5a :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h5b :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h5c :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h5d :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h5e :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h5f :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h60 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h61 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h62 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h63 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h64 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h65 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h66 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h67 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h68 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h69 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h6a :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h6b :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h6c :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h6d :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h6e :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h6f :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h70 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h71 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h72 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h73 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h74 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h75 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h76 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h77 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h78 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h79 :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h7a :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h7b :
		rl_a123_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h7c :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h7d :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h7e :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	7'h7f :
		rl_a123_t8 = RG_quantized_block_rl_59 ;
	default :
		rl_a123_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_191 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a124_t8 = RG_rl_191 ;
	7'h01 :
		rl_a124_t8 = RG_rl_191 ;
	7'h02 :
		rl_a124_t8 = RG_rl_191 ;
	7'h03 :
		rl_a124_t8 = RG_rl_191 ;
	7'h04 :
		rl_a124_t8 = RG_rl_191 ;
	7'h05 :
		rl_a124_t8 = RG_rl_191 ;
	7'h06 :
		rl_a124_t8 = RG_rl_191 ;
	7'h07 :
		rl_a124_t8 = RG_rl_191 ;
	7'h08 :
		rl_a124_t8 = RG_rl_191 ;
	7'h09 :
		rl_a124_t8 = RG_rl_191 ;
	7'h0a :
		rl_a124_t8 = RG_rl_191 ;
	7'h0b :
		rl_a124_t8 = RG_rl_191 ;
	7'h0c :
		rl_a124_t8 = RG_rl_191 ;
	7'h0d :
		rl_a124_t8 = RG_rl_191 ;
	7'h0e :
		rl_a124_t8 = RG_rl_191 ;
	7'h0f :
		rl_a124_t8 = RG_rl_191 ;
	7'h10 :
		rl_a124_t8 = RG_rl_191 ;
	7'h11 :
		rl_a124_t8 = RG_rl_191 ;
	7'h12 :
		rl_a124_t8 = RG_rl_191 ;
	7'h13 :
		rl_a124_t8 = RG_rl_191 ;
	7'h14 :
		rl_a124_t8 = RG_rl_191 ;
	7'h15 :
		rl_a124_t8 = RG_rl_191 ;
	7'h16 :
		rl_a124_t8 = RG_rl_191 ;
	7'h17 :
		rl_a124_t8 = RG_rl_191 ;
	7'h18 :
		rl_a124_t8 = RG_rl_191 ;
	7'h19 :
		rl_a124_t8 = RG_rl_191 ;
	7'h1a :
		rl_a124_t8 = RG_rl_191 ;
	7'h1b :
		rl_a124_t8 = RG_rl_191 ;
	7'h1c :
		rl_a124_t8 = RG_rl_191 ;
	7'h1d :
		rl_a124_t8 = RG_rl_191 ;
	7'h1e :
		rl_a124_t8 = RG_rl_191 ;
	7'h1f :
		rl_a124_t8 = RG_rl_191 ;
	7'h20 :
		rl_a124_t8 = RG_rl_191 ;
	7'h21 :
		rl_a124_t8 = RG_rl_191 ;
	7'h22 :
		rl_a124_t8 = RG_rl_191 ;
	7'h23 :
		rl_a124_t8 = RG_rl_191 ;
	7'h24 :
		rl_a124_t8 = RG_rl_191 ;
	7'h25 :
		rl_a124_t8 = RG_rl_191 ;
	7'h26 :
		rl_a124_t8 = RG_rl_191 ;
	7'h27 :
		rl_a124_t8 = RG_rl_191 ;
	7'h28 :
		rl_a124_t8 = RG_rl_191 ;
	7'h29 :
		rl_a124_t8 = RG_rl_191 ;
	7'h2a :
		rl_a124_t8 = RG_rl_191 ;
	7'h2b :
		rl_a124_t8 = RG_rl_191 ;
	7'h2c :
		rl_a124_t8 = RG_rl_191 ;
	7'h2d :
		rl_a124_t8 = RG_rl_191 ;
	7'h2e :
		rl_a124_t8 = RG_rl_191 ;
	7'h2f :
		rl_a124_t8 = RG_rl_191 ;
	7'h30 :
		rl_a124_t8 = RG_rl_191 ;
	7'h31 :
		rl_a124_t8 = RG_rl_191 ;
	7'h32 :
		rl_a124_t8 = RG_rl_191 ;
	7'h33 :
		rl_a124_t8 = RG_rl_191 ;
	7'h34 :
		rl_a124_t8 = RG_rl_191 ;
	7'h35 :
		rl_a124_t8 = RG_rl_191 ;
	7'h36 :
		rl_a124_t8 = RG_rl_191 ;
	7'h37 :
		rl_a124_t8 = RG_rl_191 ;
	7'h38 :
		rl_a124_t8 = RG_rl_191 ;
	7'h39 :
		rl_a124_t8 = RG_rl_191 ;
	7'h3a :
		rl_a124_t8 = RG_rl_191 ;
	7'h3b :
		rl_a124_t8 = RG_rl_191 ;
	7'h3c :
		rl_a124_t8 = RG_rl_191 ;
	7'h3d :
		rl_a124_t8 = RG_rl_191 ;
	7'h3e :
		rl_a124_t8 = RG_rl_191 ;
	7'h3f :
		rl_a124_t8 = RG_rl_191 ;
	7'h40 :
		rl_a124_t8 = RG_rl_191 ;
	7'h41 :
		rl_a124_t8 = RG_rl_191 ;
	7'h42 :
		rl_a124_t8 = RG_rl_191 ;
	7'h43 :
		rl_a124_t8 = RG_rl_191 ;
	7'h44 :
		rl_a124_t8 = RG_rl_191 ;
	7'h45 :
		rl_a124_t8 = RG_rl_191 ;
	7'h46 :
		rl_a124_t8 = RG_rl_191 ;
	7'h47 :
		rl_a124_t8 = RG_rl_191 ;
	7'h48 :
		rl_a124_t8 = RG_rl_191 ;
	7'h49 :
		rl_a124_t8 = RG_rl_191 ;
	7'h4a :
		rl_a124_t8 = RG_rl_191 ;
	7'h4b :
		rl_a124_t8 = RG_rl_191 ;
	7'h4c :
		rl_a124_t8 = RG_rl_191 ;
	7'h4d :
		rl_a124_t8 = RG_rl_191 ;
	7'h4e :
		rl_a124_t8 = RG_rl_191 ;
	7'h4f :
		rl_a124_t8 = RG_rl_191 ;
	7'h50 :
		rl_a124_t8 = RG_rl_191 ;
	7'h51 :
		rl_a124_t8 = RG_rl_191 ;
	7'h52 :
		rl_a124_t8 = RG_rl_191 ;
	7'h53 :
		rl_a124_t8 = RG_rl_191 ;
	7'h54 :
		rl_a124_t8 = RG_rl_191 ;
	7'h55 :
		rl_a124_t8 = RG_rl_191 ;
	7'h56 :
		rl_a124_t8 = RG_rl_191 ;
	7'h57 :
		rl_a124_t8 = RG_rl_191 ;
	7'h58 :
		rl_a124_t8 = RG_rl_191 ;
	7'h59 :
		rl_a124_t8 = RG_rl_191 ;
	7'h5a :
		rl_a124_t8 = RG_rl_191 ;
	7'h5b :
		rl_a124_t8 = RG_rl_191 ;
	7'h5c :
		rl_a124_t8 = RG_rl_191 ;
	7'h5d :
		rl_a124_t8 = RG_rl_191 ;
	7'h5e :
		rl_a124_t8 = RG_rl_191 ;
	7'h5f :
		rl_a124_t8 = RG_rl_191 ;
	7'h60 :
		rl_a124_t8 = RG_rl_191 ;
	7'h61 :
		rl_a124_t8 = RG_rl_191 ;
	7'h62 :
		rl_a124_t8 = RG_rl_191 ;
	7'h63 :
		rl_a124_t8 = RG_rl_191 ;
	7'h64 :
		rl_a124_t8 = RG_rl_191 ;
	7'h65 :
		rl_a124_t8 = RG_rl_191 ;
	7'h66 :
		rl_a124_t8 = RG_rl_191 ;
	7'h67 :
		rl_a124_t8 = RG_rl_191 ;
	7'h68 :
		rl_a124_t8 = RG_rl_191 ;
	7'h69 :
		rl_a124_t8 = RG_rl_191 ;
	7'h6a :
		rl_a124_t8 = RG_rl_191 ;
	7'h6b :
		rl_a124_t8 = RG_rl_191 ;
	7'h6c :
		rl_a124_t8 = RG_rl_191 ;
	7'h6d :
		rl_a124_t8 = RG_rl_191 ;
	7'h6e :
		rl_a124_t8 = RG_rl_191 ;
	7'h6f :
		rl_a124_t8 = RG_rl_191 ;
	7'h70 :
		rl_a124_t8 = RG_rl_191 ;
	7'h71 :
		rl_a124_t8 = RG_rl_191 ;
	7'h72 :
		rl_a124_t8 = RG_rl_191 ;
	7'h73 :
		rl_a124_t8 = RG_rl_191 ;
	7'h74 :
		rl_a124_t8 = RG_rl_191 ;
	7'h75 :
		rl_a124_t8 = RG_rl_191 ;
	7'h76 :
		rl_a124_t8 = RG_rl_191 ;
	7'h77 :
		rl_a124_t8 = RG_rl_191 ;
	7'h78 :
		rl_a124_t8 = RG_rl_191 ;
	7'h79 :
		rl_a124_t8 = RG_rl_191 ;
	7'h7a :
		rl_a124_t8 = RG_rl_191 ;
	7'h7b :
		rl_a124_t8 = RG_rl_191 ;
	7'h7c :
		rl_a124_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h7d :
		rl_a124_t8 = RG_rl_191 ;
	7'h7e :
		rl_a124_t8 = RG_rl_191 ;
	7'h7f :
		rl_a124_t8 = RG_rl_191 ;
	default :
		rl_a124_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_60 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h01 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h02 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h03 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h04 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h05 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h06 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h07 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h08 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h09 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h0a :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h0b :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h0c :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h0d :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h0e :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h0f :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h10 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h11 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h12 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h13 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h14 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h15 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h16 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h17 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h18 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h19 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h1a :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h1b :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h1c :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h1d :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h1e :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h1f :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h20 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h21 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h22 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h23 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h24 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h25 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h26 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h27 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h28 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h29 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h2a :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h2b :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h2c :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h2d :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h2e :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h2f :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h30 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h31 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h32 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h33 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h34 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h35 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h36 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h37 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h38 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h39 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h3a :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h3b :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h3c :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h3d :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h3e :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h3f :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h40 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h41 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h42 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h43 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h44 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h45 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h46 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h47 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h48 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h49 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h4a :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h4b :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h4c :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h4d :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h4e :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h4f :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h50 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h51 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h52 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h53 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h54 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h55 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h56 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h57 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h58 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h59 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h5a :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h5b :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h5c :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h5d :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h5e :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h5f :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h60 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h61 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h62 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h63 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h64 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h65 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h66 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h67 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h68 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h69 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h6a :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h6b :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h6c :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h6d :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h6e :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h6f :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h70 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h71 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h72 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h73 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h74 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h75 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h76 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h77 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h78 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h79 :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h7a :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h7b :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h7c :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h7d :
		rl_a125_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h7e :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	7'h7f :
		rl_a125_t8 = RG_quantized_block_rl_60 ;
	default :
		rl_a125_t8 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_quantized_block_rl_61 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h01 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h02 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h03 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h04 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h05 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h06 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h07 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h08 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h09 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h0a :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h0b :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h0c :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h0d :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h0e :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h0f :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h10 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h11 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h12 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h13 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h14 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h15 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h16 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h17 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h18 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h19 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h1a :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h1b :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h1c :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h1d :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h1e :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h1f :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h20 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h21 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h22 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h23 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h24 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h25 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h26 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h27 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h28 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h29 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h2a :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h2b :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h2c :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h2d :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h2e :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h2f :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h30 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h31 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h32 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h33 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h34 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h35 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h36 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h37 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h38 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h39 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h3a :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h3b :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h3c :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h3d :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h3e :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h3f :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h40 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h41 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h42 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h43 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h44 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h45 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h46 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h47 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h48 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h49 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h4a :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h4b :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h4c :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h4d :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h4e :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h4f :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h50 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h51 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h52 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h53 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h54 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h55 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h56 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h57 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h58 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h59 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h5a :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h5b :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h5c :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h5d :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h5e :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h5f :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h60 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h61 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h62 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h63 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h64 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h65 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h66 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h67 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h68 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h69 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h6a :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h6b :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h6c :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h6d :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h6e :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h6f :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h70 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h71 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h72 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h73 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h74 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h75 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h76 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h77 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h78 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h79 :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h7a :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h7b :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h7c :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h7d :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	7'h7e :
		rl_a126_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	7'h7f :
		rl_a126_t8 = RG_quantized_block_rl_61 ;
	default :
		rl_a126_t8 = 9'hx ;
	endcase
always @ ( RG_rl_127 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		rl_a127_t7 = RG_rl_127 ;
	7'h01 :
		rl_a127_t7 = RG_rl_127 ;
	7'h02 :
		rl_a127_t7 = RG_rl_127 ;
	7'h03 :
		rl_a127_t7 = RG_rl_127 ;
	7'h04 :
		rl_a127_t7 = RG_rl_127 ;
	7'h05 :
		rl_a127_t7 = RG_rl_127 ;
	7'h06 :
		rl_a127_t7 = RG_rl_127 ;
	7'h07 :
		rl_a127_t7 = RG_rl_127 ;
	7'h08 :
		rl_a127_t7 = RG_rl_127 ;
	7'h09 :
		rl_a127_t7 = RG_rl_127 ;
	7'h0a :
		rl_a127_t7 = RG_rl_127 ;
	7'h0b :
		rl_a127_t7 = RG_rl_127 ;
	7'h0c :
		rl_a127_t7 = RG_rl_127 ;
	7'h0d :
		rl_a127_t7 = RG_rl_127 ;
	7'h0e :
		rl_a127_t7 = RG_rl_127 ;
	7'h0f :
		rl_a127_t7 = RG_rl_127 ;
	7'h10 :
		rl_a127_t7 = RG_rl_127 ;
	7'h11 :
		rl_a127_t7 = RG_rl_127 ;
	7'h12 :
		rl_a127_t7 = RG_rl_127 ;
	7'h13 :
		rl_a127_t7 = RG_rl_127 ;
	7'h14 :
		rl_a127_t7 = RG_rl_127 ;
	7'h15 :
		rl_a127_t7 = RG_rl_127 ;
	7'h16 :
		rl_a127_t7 = RG_rl_127 ;
	7'h17 :
		rl_a127_t7 = RG_rl_127 ;
	7'h18 :
		rl_a127_t7 = RG_rl_127 ;
	7'h19 :
		rl_a127_t7 = RG_rl_127 ;
	7'h1a :
		rl_a127_t7 = RG_rl_127 ;
	7'h1b :
		rl_a127_t7 = RG_rl_127 ;
	7'h1c :
		rl_a127_t7 = RG_rl_127 ;
	7'h1d :
		rl_a127_t7 = RG_rl_127 ;
	7'h1e :
		rl_a127_t7 = RG_rl_127 ;
	7'h1f :
		rl_a127_t7 = RG_rl_127 ;
	7'h20 :
		rl_a127_t7 = RG_rl_127 ;
	7'h21 :
		rl_a127_t7 = RG_rl_127 ;
	7'h22 :
		rl_a127_t7 = RG_rl_127 ;
	7'h23 :
		rl_a127_t7 = RG_rl_127 ;
	7'h24 :
		rl_a127_t7 = RG_rl_127 ;
	7'h25 :
		rl_a127_t7 = RG_rl_127 ;
	7'h26 :
		rl_a127_t7 = RG_rl_127 ;
	7'h27 :
		rl_a127_t7 = RG_rl_127 ;
	7'h28 :
		rl_a127_t7 = RG_rl_127 ;
	7'h29 :
		rl_a127_t7 = RG_rl_127 ;
	7'h2a :
		rl_a127_t7 = RG_rl_127 ;
	7'h2b :
		rl_a127_t7 = RG_rl_127 ;
	7'h2c :
		rl_a127_t7 = RG_rl_127 ;
	7'h2d :
		rl_a127_t7 = RG_rl_127 ;
	7'h2e :
		rl_a127_t7 = RG_rl_127 ;
	7'h2f :
		rl_a127_t7 = RG_rl_127 ;
	7'h30 :
		rl_a127_t7 = RG_rl_127 ;
	7'h31 :
		rl_a127_t7 = RG_rl_127 ;
	7'h32 :
		rl_a127_t7 = RG_rl_127 ;
	7'h33 :
		rl_a127_t7 = RG_rl_127 ;
	7'h34 :
		rl_a127_t7 = RG_rl_127 ;
	7'h35 :
		rl_a127_t7 = RG_rl_127 ;
	7'h36 :
		rl_a127_t7 = RG_rl_127 ;
	7'h37 :
		rl_a127_t7 = RG_rl_127 ;
	7'h38 :
		rl_a127_t7 = RG_rl_127 ;
	7'h39 :
		rl_a127_t7 = RG_rl_127 ;
	7'h3a :
		rl_a127_t7 = RG_rl_127 ;
	7'h3b :
		rl_a127_t7 = RG_rl_127 ;
	7'h3c :
		rl_a127_t7 = RG_rl_127 ;
	7'h3d :
		rl_a127_t7 = RG_rl_127 ;
	7'h3e :
		rl_a127_t7 = RG_rl_127 ;
	7'h3f :
		rl_a127_t7 = RG_rl_127 ;
	7'h40 :
		rl_a127_t7 = RG_rl_127 ;
	7'h41 :
		rl_a127_t7 = RG_rl_127 ;
	7'h42 :
		rl_a127_t7 = RG_rl_127 ;
	7'h43 :
		rl_a127_t7 = RG_rl_127 ;
	7'h44 :
		rl_a127_t7 = RG_rl_127 ;
	7'h45 :
		rl_a127_t7 = RG_rl_127 ;
	7'h46 :
		rl_a127_t7 = RG_rl_127 ;
	7'h47 :
		rl_a127_t7 = RG_rl_127 ;
	7'h48 :
		rl_a127_t7 = RG_rl_127 ;
	7'h49 :
		rl_a127_t7 = RG_rl_127 ;
	7'h4a :
		rl_a127_t7 = RG_rl_127 ;
	7'h4b :
		rl_a127_t7 = RG_rl_127 ;
	7'h4c :
		rl_a127_t7 = RG_rl_127 ;
	7'h4d :
		rl_a127_t7 = RG_rl_127 ;
	7'h4e :
		rl_a127_t7 = RG_rl_127 ;
	7'h4f :
		rl_a127_t7 = RG_rl_127 ;
	7'h50 :
		rl_a127_t7 = RG_rl_127 ;
	7'h51 :
		rl_a127_t7 = RG_rl_127 ;
	7'h52 :
		rl_a127_t7 = RG_rl_127 ;
	7'h53 :
		rl_a127_t7 = RG_rl_127 ;
	7'h54 :
		rl_a127_t7 = RG_rl_127 ;
	7'h55 :
		rl_a127_t7 = RG_rl_127 ;
	7'h56 :
		rl_a127_t7 = RG_rl_127 ;
	7'h57 :
		rl_a127_t7 = RG_rl_127 ;
	7'h58 :
		rl_a127_t7 = RG_rl_127 ;
	7'h59 :
		rl_a127_t7 = RG_rl_127 ;
	7'h5a :
		rl_a127_t7 = RG_rl_127 ;
	7'h5b :
		rl_a127_t7 = RG_rl_127 ;
	7'h5c :
		rl_a127_t7 = RG_rl_127 ;
	7'h5d :
		rl_a127_t7 = RG_rl_127 ;
	7'h5e :
		rl_a127_t7 = RG_rl_127 ;
	7'h5f :
		rl_a127_t7 = RG_rl_127 ;
	7'h60 :
		rl_a127_t7 = RG_rl_127 ;
	7'h61 :
		rl_a127_t7 = RG_rl_127 ;
	7'h62 :
		rl_a127_t7 = RG_rl_127 ;
	7'h63 :
		rl_a127_t7 = RG_rl_127 ;
	7'h64 :
		rl_a127_t7 = RG_rl_127 ;
	7'h65 :
		rl_a127_t7 = RG_rl_127 ;
	7'h66 :
		rl_a127_t7 = RG_rl_127 ;
	7'h67 :
		rl_a127_t7 = RG_rl_127 ;
	7'h68 :
		rl_a127_t7 = RG_rl_127 ;
	7'h69 :
		rl_a127_t7 = RG_rl_127 ;
	7'h6a :
		rl_a127_t7 = RG_rl_127 ;
	7'h6b :
		rl_a127_t7 = RG_rl_127 ;
	7'h6c :
		rl_a127_t7 = RG_rl_127 ;
	7'h6d :
		rl_a127_t7 = RG_rl_127 ;
	7'h6e :
		rl_a127_t7 = RG_rl_127 ;
	7'h6f :
		rl_a127_t7 = RG_rl_127 ;
	7'h70 :
		rl_a127_t7 = RG_rl_127 ;
	7'h71 :
		rl_a127_t7 = RG_rl_127 ;
	7'h72 :
		rl_a127_t7 = RG_rl_127 ;
	7'h73 :
		rl_a127_t7 = RG_rl_127 ;
	7'h74 :
		rl_a127_t7 = RG_rl_127 ;
	7'h75 :
		rl_a127_t7 = RG_rl_127 ;
	7'h76 :
		rl_a127_t7 = RG_rl_127 ;
	7'h77 :
		rl_a127_t7 = RG_rl_127 ;
	7'h78 :
		rl_a127_t7 = RG_rl_127 ;
	7'h79 :
		rl_a127_t7 = RG_rl_127 ;
	7'h7a :
		rl_a127_t7 = RG_rl_127 ;
	7'h7b :
		rl_a127_t7 = RG_rl_127 ;
	7'h7c :
		rl_a127_t7 = RG_rl_127 ;
	7'h7d :
		rl_a127_t7 = RG_rl_127 ;
	7'h7e :
		rl_a127_t7 = RG_rl_127 ;
	7'h7f :
		rl_a127_t7 = 9'h000 ;	// line#=../rle.cpp:68
	default :
		rl_a127_t7 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01 or RG_rl_127 or RG_len )	// line#=../rle.cpp:73
	case ( RG_len [6:0] )
	7'h00 :
		rl_a127_t8 = RG_rl_127 ;
	7'h01 :
		rl_a127_t8 = RG_rl_127 ;
	7'h02 :
		rl_a127_t8 = RG_rl_127 ;
	7'h03 :
		rl_a127_t8 = RG_rl_127 ;
	7'h04 :
		rl_a127_t8 = RG_rl_127 ;
	7'h05 :
		rl_a127_t8 = RG_rl_127 ;
	7'h06 :
		rl_a127_t8 = RG_rl_127 ;
	7'h07 :
		rl_a127_t8 = RG_rl_127 ;
	7'h08 :
		rl_a127_t8 = RG_rl_127 ;
	7'h09 :
		rl_a127_t8 = RG_rl_127 ;
	7'h0a :
		rl_a127_t8 = RG_rl_127 ;
	7'h0b :
		rl_a127_t8 = RG_rl_127 ;
	7'h0c :
		rl_a127_t8 = RG_rl_127 ;
	7'h0d :
		rl_a127_t8 = RG_rl_127 ;
	7'h0e :
		rl_a127_t8 = RG_rl_127 ;
	7'h0f :
		rl_a127_t8 = RG_rl_127 ;
	7'h10 :
		rl_a127_t8 = RG_rl_127 ;
	7'h11 :
		rl_a127_t8 = RG_rl_127 ;
	7'h12 :
		rl_a127_t8 = RG_rl_127 ;
	7'h13 :
		rl_a127_t8 = RG_rl_127 ;
	7'h14 :
		rl_a127_t8 = RG_rl_127 ;
	7'h15 :
		rl_a127_t8 = RG_rl_127 ;
	7'h16 :
		rl_a127_t8 = RG_rl_127 ;
	7'h17 :
		rl_a127_t8 = RG_rl_127 ;
	7'h18 :
		rl_a127_t8 = RG_rl_127 ;
	7'h19 :
		rl_a127_t8 = RG_rl_127 ;
	7'h1a :
		rl_a127_t8 = RG_rl_127 ;
	7'h1b :
		rl_a127_t8 = RG_rl_127 ;
	7'h1c :
		rl_a127_t8 = RG_rl_127 ;
	7'h1d :
		rl_a127_t8 = RG_rl_127 ;
	7'h1e :
		rl_a127_t8 = RG_rl_127 ;
	7'h1f :
		rl_a127_t8 = RG_rl_127 ;
	7'h20 :
		rl_a127_t8 = RG_rl_127 ;
	7'h21 :
		rl_a127_t8 = RG_rl_127 ;
	7'h22 :
		rl_a127_t8 = RG_rl_127 ;
	7'h23 :
		rl_a127_t8 = RG_rl_127 ;
	7'h24 :
		rl_a127_t8 = RG_rl_127 ;
	7'h25 :
		rl_a127_t8 = RG_rl_127 ;
	7'h26 :
		rl_a127_t8 = RG_rl_127 ;
	7'h27 :
		rl_a127_t8 = RG_rl_127 ;
	7'h28 :
		rl_a127_t8 = RG_rl_127 ;
	7'h29 :
		rl_a127_t8 = RG_rl_127 ;
	7'h2a :
		rl_a127_t8 = RG_rl_127 ;
	7'h2b :
		rl_a127_t8 = RG_rl_127 ;
	7'h2c :
		rl_a127_t8 = RG_rl_127 ;
	7'h2d :
		rl_a127_t8 = RG_rl_127 ;
	7'h2e :
		rl_a127_t8 = RG_rl_127 ;
	7'h2f :
		rl_a127_t8 = RG_rl_127 ;
	7'h30 :
		rl_a127_t8 = RG_rl_127 ;
	7'h31 :
		rl_a127_t8 = RG_rl_127 ;
	7'h32 :
		rl_a127_t8 = RG_rl_127 ;
	7'h33 :
		rl_a127_t8 = RG_rl_127 ;
	7'h34 :
		rl_a127_t8 = RG_rl_127 ;
	7'h35 :
		rl_a127_t8 = RG_rl_127 ;
	7'h36 :
		rl_a127_t8 = RG_rl_127 ;
	7'h37 :
		rl_a127_t8 = RG_rl_127 ;
	7'h38 :
		rl_a127_t8 = RG_rl_127 ;
	7'h39 :
		rl_a127_t8 = RG_rl_127 ;
	7'h3a :
		rl_a127_t8 = RG_rl_127 ;
	7'h3b :
		rl_a127_t8 = RG_rl_127 ;
	7'h3c :
		rl_a127_t8 = RG_rl_127 ;
	7'h3d :
		rl_a127_t8 = RG_rl_127 ;
	7'h3e :
		rl_a127_t8 = RG_rl_127 ;
	7'h3f :
		rl_a127_t8 = RG_rl_127 ;
	7'h40 :
		rl_a127_t8 = RG_rl_127 ;
	7'h41 :
		rl_a127_t8 = RG_rl_127 ;
	7'h42 :
		rl_a127_t8 = RG_rl_127 ;
	7'h43 :
		rl_a127_t8 = RG_rl_127 ;
	7'h44 :
		rl_a127_t8 = RG_rl_127 ;
	7'h45 :
		rl_a127_t8 = RG_rl_127 ;
	7'h46 :
		rl_a127_t8 = RG_rl_127 ;
	7'h47 :
		rl_a127_t8 = RG_rl_127 ;
	7'h48 :
		rl_a127_t8 = RG_rl_127 ;
	7'h49 :
		rl_a127_t8 = RG_rl_127 ;
	7'h4a :
		rl_a127_t8 = RG_rl_127 ;
	7'h4b :
		rl_a127_t8 = RG_rl_127 ;
	7'h4c :
		rl_a127_t8 = RG_rl_127 ;
	7'h4d :
		rl_a127_t8 = RG_rl_127 ;
	7'h4e :
		rl_a127_t8 = RG_rl_127 ;
	7'h4f :
		rl_a127_t8 = RG_rl_127 ;
	7'h50 :
		rl_a127_t8 = RG_rl_127 ;
	7'h51 :
		rl_a127_t8 = RG_rl_127 ;
	7'h52 :
		rl_a127_t8 = RG_rl_127 ;
	7'h53 :
		rl_a127_t8 = RG_rl_127 ;
	7'h54 :
		rl_a127_t8 = RG_rl_127 ;
	7'h55 :
		rl_a127_t8 = RG_rl_127 ;
	7'h56 :
		rl_a127_t8 = RG_rl_127 ;
	7'h57 :
		rl_a127_t8 = RG_rl_127 ;
	7'h58 :
		rl_a127_t8 = RG_rl_127 ;
	7'h59 :
		rl_a127_t8 = RG_rl_127 ;
	7'h5a :
		rl_a127_t8 = RG_rl_127 ;
	7'h5b :
		rl_a127_t8 = RG_rl_127 ;
	7'h5c :
		rl_a127_t8 = RG_rl_127 ;
	7'h5d :
		rl_a127_t8 = RG_rl_127 ;
	7'h5e :
		rl_a127_t8 = RG_rl_127 ;
	7'h5f :
		rl_a127_t8 = RG_rl_127 ;
	7'h60 :
		rl_a127_t8 = RG_rl_127 ;
	7'h61 :
		rl_a127_t8 = RG_rl_127 ;
	7'h62 :
		rl_a127_t8 = RG_rl_127 ;
	7'h63 :
		rl_a127_t8 = RG_rl_127 ;
	7'h64 :
		rl_a127_t8 = RG_rl_127 ;
	7'h65 :
		rl_a127_t8 = RG_rl_127 ;
	7'h66 :
		rl_a127_t8 = RG_rl_127 ;
	7'h67 :
		rl_a127_t8 = RG_rl_127 ;
	7'h68 :
		rl_a127_t8 = RG_rl_127 ;
	7'h69 :
		rl_a127_t8 = RG_rl_127 ;
	7'h6a :
		rl_a127_t8 = RG_rl_127 ;
	7'h6b :
		rl_a127_t8 = RG_rl_127 ;
	7'h6c :
		rl_a127_t8 = RG_rl_127 ;
	7'h6d :
		rl_a127_t8 = RG_rl_127 ;
	7'h6e :
		rl_a127_t8 = RG_rl_127 ;
	7'h6f :
		rl_a127_t8 = RG_rl_127 ;
	7'h70 :
		rl_a127_t8 = RG_rl_127 ;
	7'h71 :
		rl_a127_t8 = RG_rl_127 ;
	7'h72 :
		rl_a127_t8 = RG_rl_127 ;
	7'h73 :
		rl_a127_t8 = RG_rl_127 ;
	7'h74 :
		rl_a127_t8 = RG_rl_127 ;
	7'h75 :
		rl_a127_t8 = RG_rl_127 ;
	7'h76 :
		rl_a127_t8 = RG_rl_127 ;
	7'h77 :
		rl_a127_t8 = RG_rl_127 ;
	7'h78 :
		rl_a127_t8 = RG_rl_127 ;
	7'h79 :
		rl_a127_t8 = RG_rl_127 ;
	7'h7a :
		rl_a127_t8 = RG_rl_127 ;
	7'h7b :
		rl_a127_t8 = RG_rl_127 ;
	7'h7c :
		rl_a127_t8 = RG_rl_127 ;
	7'h7d :
		rl_a127_t8 = RG_rl_127 ;
	7'h7e :
		rl_a127_t8 = RG_rl_127 ;
	7'h7f :
		rl_a127_t8 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:73
	default :
		rl_a127_t8 = 9'hx ;
	endcase
assign	sub8u1i1 = RG_len_1 ;	// line#=../rle.cpp:86
assign	sub8u1i2 = 2'h2 ;	// line#=../rle.cpp:86
assign	sub12s_91i1 = RG_previous_dc_zz ;	// line#=../rle.cpp:52
assign	sub12s_91i2 = RG_previous_dc_rl ;	// line#=../rle.cpp:52
assign	lop8u_11i1 = RG_k ;	// line#=../rle.cpp:109,110
assign	lop8u_11i2 = 6'h24 ;	// line#=../rle.cpp:109,110
assign	incr4s1i1 = RG_j ;	// line#=../rle.cpp:34
assign	incr8u2i1 = RG_len ;	// line#=../rle.cpp:73
assign	decr8u_71i1 = RG_len [6:0] ;	// line#=../rle.cpp:77,78
assign	sub8u_71i1 = RG_len_1 [6:0] ;	// line#=../rle.cpp:83,84
assign	sub8u_71i2 = 3'h4 ;	// line#=../rle.cpp:83,84
assign	C_01 = ~|{ ~incr4s1ot [3] , incr4s1ot [2:0] } ;	// line#=../rle.cpp:34,35
assign	U_01 = ( ST1_02d & C_01 ) ;	// line#=../rle.cpp:35
assign	U_05 = ( ST1_03d & lop8u_11ot ) ;	// line#=../rle.cpp:109,110
assign	U_06 = ( ST1_03d & ( ~lop8u_11ot ) ) ;	// line#=../rle.cpp:109,110
assign	C_02 = ( ( ~|RG_i_k_01 ) & M_48 ) ;	// line#=../rle.cpp:112,113
assign	U_79 = ( U_05 & C_02 ) ;	// line#=../rle.cpp:112,113
assign	U_80 = ( U_05 & ( ~C_02 ) ) ;	// line#=../rle.cpp:112,113
assign	U_81 = ( U_80 & CT_03 ) ;	// line#=../rle.cpp:117,118
assign	U_82 = ( U_80 & ( ~CT_03 ) ) ;	// line#=../rle.cpp:117,118
assign	U_83 = ( U_82 & ( ~FF_d ) ) ;	// line#=../rle.cpp:122,123
assign	U_84 = ( U_82 & FF_d ) ;	// line#=../rle.cpp:122,123
assign	U_87 = ( ST1_04d & ( ~RG_k_1 [6] ) ) ;	// line#=../rle.cpp:140,141
assign	U_88 = ( ST1_04d & RG_k_1 [6] ) ;	// line#=../rle.cpp:140,141
assign	M_48 = ~|{ ( RG_i_j_01 [31] & RG_i_j_01 [0] ) , RG_i_j_01 [0] } ;	// line#=../rle.cpp:112,113,143,144
assign	C_05 = ( ( ~|{ RG_i_k_01 [31:3] , ~RG_i_k_01 [2:0] } ) & M_48 ) ;	// line#=../rle.cpp:143,144
assign	U_161 = ( U_87 & C_05 ) ;	// line#=../rle.cpp:143,144
assign	U_162 = ( U_87 & ( ~C_05 ) ) ;	// line#=../rle.cpp:143,144
assign	U_163 = ( U_162 & CT_18 ) ;	// line#=../rle.cpp:148,149
assign	U_164 = ( U_162 & ( ~CT_18 ) ) ;	// line#=../rle.cpp:148,149
assign	U_165 = ( U_164 & ( ~FF_d ) ) ;	// line#=../rle.cpp:153,154
assign	U_166 = ( U_164 & FF_d ) ;	// line#=../rle.cpp:153,154
assign	C_07 = ( RG_i_j_01 [31] | ( ~|RG_i_j_01 [30:6] ) ) ;	// line#=../rle.cpp:57,58,61,62
assign	C_07_port = C_07 ;
assign	U_170 = ( ST1_05d & ( ~C_07 ) ) ;	// line#=../rle.cpp:57,58
assign	U_173 = ( U_170 & ( ~M_02_t128 ) ) ;	// line#=../rle.cpp:77,78
assign	U_174 = ( U_170 & M_02_t128 ) ;	// line#=../rle.cpp:77,78
assign	C_08 = ( M_01_t64 & ( RG_i_k_01 [31] | ( ( ~|RG_i_k_01 [30:4] ) & ( ~&RG_i_k_01 [3:0] ) ) ) ) ;	// line#=../rle.cpp:61,62
assign	C_08_port = C_08 ;
assign	U_183 = ( ST1_07d & M_03_t128 ) ;	// line#=../rle.cpp:83,84
assign	U_184 = ( ST1_07d & ( ~M_03_t128 ) ) ;	// line#=../rle.cpp:83,84
assign	C_09 = ~|{ RG_i_j_01 [31:7] , ~RG_i_j_01 [6] , RG_i_j_01 [5:0] } ;	// line#=../rle.cpp:66,67
assign	U_317 = ( ST1_08d & C_09 ) ;	// line#=../rle.cpp:66,67
assign	U_318 = ( ST1_08d & ( ~C_09 ) ) ;	// line#=../rle.cpp:66,67
always @ ( TR_12 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_265 = 9'h000 ;	// line#=../rle.cpp:80
	7'h01 :
		TR_265 = TR_12 ;
	7'h02 :
		TR_265 = TR_12 ;
	7'h03 :
		TR_265 = TR_12 ;
	7'h04 :
		TR_265 = TR_12 ;
	7'h05 :
		TR_265 = TR_12 ;
	7'h06 :
		TR_265 = TR_12 ;
	7'h07 :
		TR_265 = TR_12 ;
	7'h08 :
		TR_265 = TR_12 ;
	7'h09 :
		TR_265 = TR_12 ;
	7'h0a :
		TR_265 = TR_12 ;
	7'h0b :
		TR_265 = TR_12 ;
	7'h0c :
		TR_265 = TR_12 ;
	7'h0d :
		TR_265 = TR_12 ;
	7'h0e :
		TR_265 = TR_12 ;
	7'h0f :
		TR_265 = TR_12 ;
	7'h10 :
		TR_265 = TR_12 ;
	7'h11 :
		TR_265 = TR_12 ;
	7'h12 :
		TR_265 = TR_12 ;
	7'h13 :
		TR_265 = TR_12 ;
	7'h14 :
		TR_265 = TR_12 ;
	7'h15 :
		TR_265 = TR_12 ;
	7'h16 :
		TR_265 = TR_12 ;
	7'h17 :
		TR_265 = TR_12 ;
	7'h18 :
		TR_265 = TR_12 ;
	7'h19 :
		TR_265 = TR_12 ;
	7'h1a :
		TR_265 = TR_12 ;
	7'h1b :
		TR_265 = TR_12 ;
	7'h1c :
		TR_265 = TR_12 ;
	7'h1d :
		TR_265 = TR_12 ;
	7'h1e :
		TR_265 = TR_12 ;
	7'h1f :
		TR_265 = TR_12 ;
	7'h20 :
		TR_265 = TR_12 ;
	7'h21 :
		TR_265 = TR_12 ;
	7'h22 :
		TR_265 = TR_12 ;
	7'h23 :
		TR_265 = TR_12 ;
	7'h24 :
		TR_265 = TR_12 ;
	7'h25 :
		TR_265 = TR_12 ;
	7'h26 :
		TR_265 = TR_12 ;
	7'h27 :
		TR_265 = TR_12 ;
	7'h28 :
		TR_265 = TR_12 ;
	7'h29 :
		TR_265 = TR_12 ;
	7'h2a :
		TR_265 = TR_12 ;
	7'h2b :
		TR_265 = TR_12 ;
	7'h2c :
		TR_265 = TR_12 ;
	7'h2d :
		TR_265 = TR_12 ;
	7'h2e :
		TR_265 = TR_12 ;
	7'h2f :
		TR_265 = TR_12 ;
	7'h30 :
		TR_265 = TR_12 ;
	7'h31 :
		TR_265 = TR_12 ;
	7'h32 :
		TR_265 = TR_12 ;
	7'h33 :
		TR_265 = TR_12 ;
	7'h34 :
		TR_265 = TR_12 ;
	7'h35 :
		TR_265 = TR_12 ;
	7'h36 :
		TR_265 = TR_12 ;
	7'h37 :
		TR_265 = TR_12 ;
	7'h38 :
		TR_265 = TR_12 ;
	7'h39 :
		TR_265 = TR_12 ;
	7'h3a :
		TR_265 = TR_12 ;
	7'h3b :
		TR_265 = TR_12 ;
	7'h3c :
		TR_265 = TR_12 ;
	7'h3d :
		TR_265 = TR_12 ;
	7'h3e :
		TR_265 = TR_12 ;
	7'h3f :
		TR_265 = TR_12 ;
	7'h40 :
		TR_265 = TR_12 ;
	7'h41 :
		TR_265 = TR_12 ;
	7'h42 :
		TR_265 = TR_12 ;
	7'h43 :
		TR_265 = TR_12 ;
	7'h44 :
		TR_265 = TR_12 ;
	7'h45 :
		TR_265 = TR_12 ;
	7'h46 :
		TR_265 = TR_12 ;
	7'h47 :
		TR_265 = TR_12 ;
	7'h48 :
		TR_265 = TR_12 ;
	7'h49 :
		TR_265 = TR_12 ;
	7'h4a :
		TR_265 = TR_12 ;
	7'h4b :
		TR_265 = TR_12 ;
	7'h4c :
		TR_265 = TR_12 ;
	7'h4d :
		TR_265 = TR_12 ;
	7'h4e :
		TR_265 = TR_12 ;
	7'h4f :
		TR_265 = TR_12 ;
	7'h50 :
		TR_265 = TR_12 ;
	7'h51 :
		TR_265 = TR_12 ;
	7'h52 :
		TR_265 = TR_12 ;
	7'h53 :
		TR_265 = TR_12 ;
	7'h54 :
		TR_265 = TR_12 ;
	7'h55 :
		TR_265 = TR_12 ;
	7'h56 :
		TR_265 = TR_12 ;
	7'h57 :
		TR_265 = TR_12 ;
	7'h58 :
		TR_265 = TR_12 ;
	7'h59 :
		TR_265 = TR_12 ;
	7'h5a :
		TR_265 = TR_12 ;
	7'h5b :
		TR_265 = TR_12 ;
	7'h5c :
		TR_265 = TR_12 ;
	7'h5d :
		TR_265 = TR_12 ;
	7'h5e :
		TR_265 = TR_12 ;
	7'h5f :
		TR_265 = TR_12 ;
	7'h60 :
		TR_265 = TR_12 ;
	7'h61 :
		TR_265 = TR_12 ;
	7'h62 :
		TR_265 = TR_12 ;
	7'h63 :
		TR_265 = TR_12 ;
	7'h64 :
		TR_265 = TR_12 ;
	7'h65 :
		TR_265 = TR_12 ;
	7'h66 :
		TR_265 = TR_12 ;
	7'h67 :
		TR_265 = TR_12 ;
	7'h68 :
		TR_265 = TR_12 ;
	7'h69 :
		TR_265 = TR_12 ;
	7'h6a :
		TR_265 = TR_12 ;
	7'h6b :
		TR_265 = TR_12 ;
	7'h6c :
		TR_265 = TR_12 ;
	7'h6d :
		TR_265 = TR_12 ;
	7'h6e :
		TR_265 = TR_12 ;
	7'h6f :
		TR_265 = TR_12 ;
	7'h70 :
		TR_265 = TR_12 ;
	7'h71 :
		TR_265 = TR_12 ;
	7'h72 :
		TR_265 = TR_12 ;
	7'h73 :
		TR_265 = TR_12 ;
	7'h74 :
		TR_265 = TR_12 ;
	7'h75 :
		TR_265 = TR_12 ;
	7'h76 :
		TR_265 = TR_12 ;
	7'h77 :
		TR_265 = TR_12 ;
	7'h78 :
		TR_265 = TR_12 ;
	7'h79 :
		TR_265 = TR_12 ;
	7'h7a :
		TR_265 = TR_12 ;
	7'h7b :
		TR_265 = TR_12 ;
	7'h7c :
		TR_265 = TR_12 ;
	7'h7d :
		TR_265 = TR_12 ;
	7'h7e :
		TR_265 = TR_12 ;
	7'h7f :
		TR_265 = TR_12 ;
	default :
		TR_265 = 9'hx ;
	endcase
always @ ( TR_265 or U_173 or sub8u_71ot or U_183 or RG_previous_dc_rl or U_174 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_t_c1 = ( U_183 & ( ~|sub8u_71ot ) ) ;	// line#=../rle.cpp:85
	RG_rl_t = ( ( { 9{ U_174 } } & RG_previous_dc_rl )
		| ( { 9{ U_173 } } & TR_265 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_en = ( U_174 | RG_rl_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_en )
		RG_rl <= RG_rl_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( RG_quantized_block_rl_zz or U_184 or RG_k_1 or U_87 or M_184 or RG_k or 
	U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_previous_dc_zz_t_c1 = ( U_05 & ( ~|RG_k ) ) ;	// line#=../rle.cpp:111
	RG_previous_dc_zz_t_c2 = ( U_87 & ( ~|RG_k_1 [5:0] ) ) ;	// line#=../rle.cpp:142
	RG_previous_dc_zz_t = ( ( { 9{ RG_previous_dc_zz_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_previous_dc_zz_t_c2 } } & M_184 )			// line#=../rle.cpp:142
		| ( { 9{ U_184 } } & RG_quantized_block_rl_zz ) ) ;
	end
assign	RG_previous_dc_zz_en = ( RG_previous_dc_zz_t_c1 | RG_previous_dc_zz_t_c2 | 
	U_184 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_previous_dc_zz_en )
		RG_previous_dc_zz <= RG_previous_dc_zz_t ;	// line#=../rle.cpp:111,142
always @ ( TR_13 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_264 = TR_13 ;
	7'h01 :
		TR_264 = 9'h000 ;	// line#=../rle.cpp:80
	7'h02 :
		TR_264 = TR_13 ;
	7'h03 :
		TR_264 = TR_13 ;
	7'h04 :
		TR_264 = TR_13 ;
	7'h05 :
		TR_264 = TR_13 ;
	7'h06 :
		TR_264 = TR_13 ;
	7'h07 :
		TR_264 = TR_13 ;
	7'h08 :
		TR_264 = TR_13 ;
	7'h09 :
		TR_264 = TR_13 ;
	7'h0a :
		TR_264 = TR_13 ;
	7'h0b :
		TR_264 = TR_13 ;
	7'h0c :
		TR_264 = TR_13 ;
	7'h0d :
		TR_264 = TR_13 ;
	7'h0e :
		TR_264 = TR_13 ;
	7'h0f :
		TR_264 = TR_13 ;
	7'h10 :
		TR_264 = TR_13 ;
	7'h11 :
		TR_264 = TR_13 ;
	7'h12 :
		TR_264 = TR_13 ;
	7'h13 :
		TR_264 = TR_13 ;
	7'h14 :
		TR_264 = TR_13 ;
	7'h15 :
		TR_264 = TR_13 ;
	7'h16 :
		TR_264 = TR_13 ;
	7'h17 :
		TR_264 = TR_13 ;
	7'h18 :
		TR_264 = TR_13 ;
	7'h19 :
		TR_264 = TR_13 ;
	7'h1a :
		TR_264 = TR_13 ;
	7'h1b :
		TR_264 = TR_13 ;
	7'h1c :
		TR_264 = TR_13 ;
	7'h1d :
		TR_264 = TR_13 ;
	7'h1e :
		TR_264 = TR_13 ;
	7'h1f :
		TR_264 = TR_13 ;
	7'h20 :
		TR_264 = TR_13 ;
	7'h21 :
		TR_264 = TR_13 ;
	7'h22 :
		TR_264 = TR_13 ;
	7'h23 :
		TR_264 = TR_13 ;
	7'h24 :
		TR_264 = TR_13 ;
	7'h25 :
		TR_264 = TR_13 ;
	7'h26 :
		TR_264 = TR_13 ;
	7'h27 :
		TR_264 = TR_13 ;
	7'h28 :
		TR_264 = TR_13 ;
	7'h29 :
		TR_264 = TR_13 ;
	7'h2a :
		TR_264 = TR_13 ;
	7'h2b :
		TR_264 = TR_13 ;
	7'h2c :
		TR_264 = TR_13 ;
	7'h2d :
		TR_264 = TR_13 ;
	7'h2e :
		TR_264 = TR_13 ;
	7'h2f :
		TR_264 = TR_13 ;
	7'h30 :
		TR_264 = TR_13 ;
	7'h31 :
		TR_264 = TR_13 ;
	7'h32 :
		TR_264 = TR_13 ;
	7'h33 :
		TR_264 = TR_13 ;
	7'h34 :
		TR_264 = TR_13 ;
	7'h35 :
		TR_264 = TR_13 ;
	7'h36 :
		TR_264 = TR_13 ;
	7'h37 :
		TR_264 = TR_13 ;
	7'h38 :
		TR_264 = TR_13 ;
	7'h39 :
		TR_264 = TR_13 ;
	7'h3a :
		TR_264 = TR_13 ;
	7'h3b :
		TR_264 = TR_13 ;
	7'h3c :
		TR_264 = TR_13 ;
	7'h3d :
		TR_264 = TR_13 ;
	7'h3e :
		TR_264 = TR_13 ;
	7'h3f :
		TR_264 = TR_13 ;
	7'h40 :
		TR_264 = TR_13 ;
	7'h41 :
		TR_264 = TR_13 ;
	7'h42 :
		TR_264 = TR_13 ;
	7'h43 :
		TR_264 = TR_13 ;
	7'h44 :
		TR_264 = TR_13 ;
	7'h45 :
		TR_264 = TR_13 ;
	7'h46 :
		TR_264 = TR_13 ;
	7'h47 :
		TR_264 = TR_13 ;
	7'h48 :
		TR_264 = TR_13 ;
	7'h49 :
		TR_264 = TR_13 ;
	7'h4a :
		TR_264 = TR_13 ;
	7'h4b :
		TR_264 = TR_13 ;
	7'h4c :
		TR_264 = TR_13 ;
	7'h4d :
		TR_264 = TR_13 ;
	7'h4e :
		TR_264 = TR_13 ;
	7'h4f :
		TR_264 = TR_13 ;
	7'h50 :
		TR_264 = TR_13 ;
	7'h51 :
		TR_264 = TR_13 ;
	7'h52 :
		TR_264 = TR_13 ;
	7'h53 :
		TR_264 = TR_13 ;
	7'h54 :
		TR_264 = TR_13 ;
	7'h55 :
		TR_264 = TR_13 ;
	7'h56 :
		TR_264 = TR_13 ;
	7'h57 :
		TR_264 = TR_13 ;
	7'h58 :
		TR_264 = TR_13 ;
	7'h59 :
		TR_264 = TR_13 ;
	7'h5a :
		TR_264 = TR_13 ;
	7'h5b :
		TR_264 = TR_13 ;
	7'h5c :
		TR_264 = TR_13 ;
	7'h5d :
		TR_264 = TR_13 ;
	7'h5e :
		TR_264 = TR_13 ;
	7'h5f :
		TR_264 = TR_13 ;
	7'h60 :
		TR_264 = TR_13 ;
	7'h61 :
		TR_264 = TR_13 ;
	7'h62 :
		TR_264 = TR_13 ;
	7'h63 :
		TR_264 = TR_13 ;
	7'h64 :
		TR_264 = TR_13 ;
	7'h65 :
		TR_264 = TR_13 ;
	7'h66 :
		TR_264 = TR_13 ;
	7'h67 :
		TR_264 = TR_13 ;
	7'h68 :
		TR_264 = TR_13 ;
	7'h69 :
		TR_264 = TR_13 ;
	7'h6a :
		TR_264 = TR_13 ;
	7'h6b :
		TR_264 = TR_13 ;
	7'h6c :
		TR_264 = TR_13 ;
	7'h6d :
		TR_264 = TR_13 ;
	7'h6e :
		TR_264 = TR_13 ;
	7'h6f :
		TR_264 = TR_13 ;
	7'h70 :
		TR_264 = TR_13 ;
	7'h71 :
		TR_264 = TR_13 ;
	7'h72 :
		TR_264 = TR_13 ;
	7'h73 :
		TR_264 = TR_13 ;
	7'h74 :
		TR_264 = TR_13 ;
	7'h75 :
		TR_264 = TR_13 ;
	7'h76 :
		TR_264 = TR_13 ;
	7'h77 :
		TR_264 = TR_13 ;
	7'h78 :
		TR_264 = TR_13 ;
	7'h79 :
		TR_264 = TR_13 ;
	7'h7a :
		TR_264 = TR_13 ;
	7'h7b :
		TR_264 = TR_13 ;
	7'h7c :
		TR_264 = TR_13 ;
	7'h7d :
		TR_264 = TR_13 ;
	7'h7e :
		TR_264 = TR_13 ;
	7'h7f :
		TR_264 = TR_13 ;
	default :
		TR_264 = 9'hx ;
	endcase
always @ ( TR_264 or U_173 or sub8u_71ot or U_183 or RG_rl_128 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_1_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h01 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_1_t = ( ( { 9{ M_180 } } & RG_rl_128 )
		| ( { 9{ U_173 } } & TR_264 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_1_en = ( M_180 | RG_rl_1_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_1_en )
		RG_rl_1 <= RG_rl_1_t ;	// line#=../rle.cpp:79,80,83,84,85
assign	M_180 = ( ST1_01d | U_174 ) ;	// line#=../rle.cpp:83,84,85
always @ ( TR_14 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_263 = TR_14 ;
	7'h01 :
		TR_263 = TR_14 ;
	7'h02 :
		TR_263 = 9'h000 ;	// line#=../rle.cpp:80
	7'h03 :
		TR_263 = TR_14 ;
	7'h04 :
		TR_263 = TR_14 ;
	7'h05 :
		TR_263 = TR_14 ;
	7'h06 :
		TR_263 = TR_14 ;
	7'h07 :
		TR_263 = TR_14 ;
	7'h08 :
		TR_263 = TR_14 ;
	7'h09 :
		TR_263 = TR_14 ;
	7'h0a :
		TR_263 = TR_14 ;
	7'h0b :
		TR_263 = TR_14 ;
	7'h0c :
		TR_263 = TR_14 ;
	7'h0d :
		TR_263 = TR_14 ;
	7'h0e :
		TR_263 = TR_14 ;
	7'h0f :
		TR_263 = TR_14 ;
	7'h10 :
		TR_263 = TR_14 ;
	7'h11 :
		TR_263 = TR_14 ;
	7'h12 :
		TR_263 = TR_14 ;
	7'h13 :
		TR_263 = TR_14 ;
	7'h14 :
		TR_263 = TR_14 ;
	7'h15 :
		TR_263 = TR_14 ;
	7'h16 :
		TR_263 = TR_14 ;
	7'h17 :
		TR_263 = TR_14 ;
	7'h18 :
		TR_263 = TR_14 ;
	7'h19 :
		TR_263 = TR_14 ;
	7'h1a :
		TR_263 = TR_14 ;
	7'h1b :
		TR_263 = TR_14 ;
	7'h1c :
		TR_263 = TR_14 ;
	7'h1d :
		TR_263 = TR_14 ;
	7'h1e :
		TR_263 = TR_14 ;
	7'h1f :
		TR_263 = TR_14 ;
	7'h20 :
		TR_263 = TR_14 ;
	7'h21 :
		TR_263 = TR_14 ;
	7'h22 :
		TR_263 = TR_14 ;
	7'h23 :
		TR_263 = TR_14 ;
	7'h24 :
		TR_263 = TR_14 ;
	7'h25 :
		TR_263 = TR_14 ;
	7'h26 :
		TR_263 = TR_14 ;
	7'h27 :
		TR_263 = TR_14 ;
	7'h28 :
		TR_263 = TR_14 ;
	7'h29 :
		TR_263 = TR_14 ;
	7'h2a :
		TR_263 = TR_14 ;
	7'h2b :
		TR_263 = TR_14 ;
	7'h2c :
		TR_263 = TR_14 ;
	7'h2d :
		TR_263 = TR_14 ;
	7'h2e :
		TR_263 = TR_14 ;
	7'h2f :
		TR_263 = TR_14 ;
	7'h30 :
		TR_263 = TR_14 ;
	7'h31 :
		TR_263 = TR_14 ;
	7'h32 :
		TR_263 = TR_14 ;
	7'h33 :
		TR_263 = TR_14 ;
	7'h34 :
		TR_263 = TR_14 ;
	7'h35 :
		TR_263 = TR_14 ;
	7'h36 :
		TR_263 = TR_14 ;
	7'h37 :
		TR_263 = TR_14 ;
	7'h38 :
		TR_263 = TR_14 ;
	7'h39 :
		TR_263 = TR_14 ;
	7'h3a :
		TR_263 = TR_14 ;
	7'h3b :
		TR_263 = TR_14 ;
	7'h3c :
		TR_263 = TR_14 ;
	7'h3d :
		TR_263 = TR_14 ;
	7'h3e :
		TR_263 = TR_14 ;
	7'h3f :
		TR_263 = TR_14 ;
	7'h40 :
		TR_263 = TR_14 ;
	7'h41 :
		TR_263 = TR_14 ;
	7'h42 :
		TR_263 = TR_14 ;
	7'h43 :
		TR_263 = TR_14 ;
	7'h44 :
		TR_263 = TR_14 ;
	7'h45 :
		TR_263 = TR_14 ;
	7'h46 :
		TR_263 = TR_14 ;
	7'h47 :
		TR_263 = TR_14 ;
	7'h48 :
		TR_263 = TR_14 ;
	7'h49 :
		TR_263 = TR_14 ;
	7'h4a :
		TR_263 = TR_14 ;
	7'h4b :
		TR_263 = TR_14 ;
	7'h4c :
		TR_263 = TR_14 ;
	7'h4d :
		TR_263 = TR_14 ;
	7'h4e :
		TR_263 = TR_14 ;
	7'h4f :
		TR_263 = TR_14 ;
	7'h50 :
		TR_263 = TR_14 ;
	7'h51 :
		TR_263 = TR_14 ;
	7'h52 :
		TR_263 = TR_14 ;
	7'h53 :
		TR_263 = TR_14 ;
	7'h54 :
		TR_263 = TR_14 ;
	7'h55 :
		TR_263 = TR_14 ;
	7'h56 :
		TR_263 = TR_14 ;
	7'h57 :
		TR_263 = TR_14 ;
	7'h58 :
		TR_263 = TR_14 ;
	7'h59 :
		TR_263 = TR_14 ;
	7'h5a :
		TR_263 = TR_14 ;
	7'h5b :
		TR_263 = TR_14 ;
	7'h5c :
		TR_263 = TR_14 ;
	7'h5d :
		TR_263 = TR_14 ;
	7'h5e :
		TR_263 = TR_14 ;
	7'h5f :
		TR_263 = TR_14 ;
	7'h60 :
		TR_263 = TR_14 ;
	7'h61 :
		TR_263 = TR_14 ;
	7'h62 :
		TR_263 = TR_14 ;
	7'h63 :
		TR_263 = TR_14 ;
	7'h64 :
		TR_263 = TR_14 ;
	7'h65 :
		TR_263 = TR_14 ;
	7'h66 :
		TR_263 = TR_14 ;
	7'h67 :
		TR_263 = TR_14 ;
	7'h68 :
		TR_263 = TR_14 ;
	7'h69 :
		TR_263 = TR_14 ;
	7'h6a :
		TR_263 = TR_14 ;
	7'h6b :
		TR_263 = TR_14 ;
	7'h6c :
		TR_263 = TR_14 ;
	7'h6d :
		TR_263 = TR_14 ;
	7'h6e :
		TR_263 = TR_14 ;
	7'h6f :
		TR_263 = TR_14 ;
	7'h70 :
		TR_263 = TR_14 ;
	7'h71 :
		TR_263 = TR_14 ;
	7'h72 :
		TR_263 = TR_14 ;
	7'h73 :
		TR_263 = TR_14 ;
	7'h74 :
		TR_263 = TR_14 ;
	7'h75 :
		TR_263 = TR_14 ;
	7'h76 :
		TR_263 = TR_14 ;
	7'h77 :
		TR_263 = TR_14 ;
	7'h78 :
		TR_263 = TR_14 ;
	7'h79 :
		TR_263 = TR_14 ;
	7'h7a :
		TR_263 = TR_14 ;
	7'h7b :
		TR_263 = TR_14 ;
	7'h7c :
		TR_263 = TR_14 ;
	7'h7d :
		TR_263 = TR_14 ;
	7'h7e :
		TR_263 = TR_14 ;
	7'h7f :
		TR_263 = TR_14 ;
	default :
		TR_263 = 9'hx ;
	endcase
always @ ( TR_263 or U_173 or sub8u_71ot or U_183 or RG_rl_129 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_2_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h02 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_2_t = ( ( { 9{ M_180 } } & RG_rl_129 )
		| ( { 9{ U_173 } } & TR_263 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_2_en = ( M_180 | RG_rl_2_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_2_en )
		RG_rl_2 <= RG_rl_2_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_15 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_262 = TR_15 ;
	7'h01 :
		TR_262 = TR_15 ;
	7'h02 :
		TR_262 = TR_15 ;
	7'h03 :
		TR_262 = 9'h000 ;	// line#=../rle.cpp:80
	7'h04 :
		TR_262 = TR_15 ;
	7'h05 :
		TR_262 = TR_15 ;
	7'h06 :
		TR_262 = TR_15 ;
	7'h07 :
		TR_262 = TR_15 ;
	7'h08 :
		TR_262 = TR_15 ;
	7'h09 :
		TR_262 = TR_15 ;
	7'h0a :
		TR_262 = TR_15 ;
	7'h0b :
		TR_262 = TR_15 ;
	7'h0c :
		TR_262 = TR_15 ;
	7'h0d :
		TR_262 = TR_15 ;
	7'h0e :
		TR_262 = TR_15 ;
	7'h0f :
		TR_262 = TR_15 ;
	7'h10 :
		TR_262 = TR_15 ;
	7'h11 :
		TR_262 = TR_15 ;
	7'h12 :
		TR_262 = TR_15 ;
	7'h13 :
		TR_262 = TR_15 ;
	7'h14 :
		TR_262 = TR_15 ;
	7'h15 :
		TR_262 = TR_15 ;
	7'h16 :
		TR_262 = TR_15 ;
	7'h17 :
		TR_262 = TR_15 ;
	7'h18 :
		TR_262 = TR_15 ;
	7'h19 :
		TR_262 = TR_15 ;
	7'h1a :
		TR_262 = TR_15 ;
	7'h1b :
		TR_262 = TR_15 ;
	7'h1c :
		TR_262 = TR_15 ;
	7'h1d :
		TR_262 = TR_15 ;
	7'h1e :
		TR_262 = TR_15 ;
	7'h1f :
		TR_262 = TR_15 ;
	7'h20 :
		TR_262 = TR_15 ;
	7'h21 :
		TR_262 = TR_15 ;
	7'h22 :
		TR_262 = TR_15 ;
	7'h23 :
		TR_262 = TR_15 ;
	7'h24 :
		TR_262 = TR_15 ;
	7'h25 :
		TR_262 = TR_15 ;
	7'h26 :
		TR_262 = TR_15 ;
	7'h27 :
		TR_262 = TR_15 ;
	7'h28 :
		TR_262 = TR_15 ;
	7'h29 :
		TR_262 = TR_15 ;
	7'h2a :
		TR_262 = TR_15 ;
	7'h2b :
		TR_262 = TR_15 ;
	7'h2c :
		TR_262 = TR_15 ;
	7'h2d :
		TR_262 = TR_15 ;
	7'h2e :
		TR_262 = TR_15 ;
	7'h2f :
		TR_262 = TR_15 ;
	7'h30 :
		TR_262 = TR_15 ;
	7'h31 :
		TR_262 = TR_15 ;
	7'h32 :
		TR_262 = TR_15 ;
	7'h33 :
		TR_262 = TR_15 ;
	7'h34 :
		TR_262 = TR_15 ;
	7'h35 :
		TR_262 = TR_15 ;
	7'h36 :
		TR_262 = TR_15 ;
	7'h37 :
		TR_262 = TR_15 ;
	7'h38 :
		TR_262 = TR_15 ;
	7'h39 :
		TR_262 = TR_15 ;
	7'h3a :
		TR_262 = TR_15 ;
	7'h3b :
		TR_262 = TR_15 ;
	7'h3c :
		TR_262 = TR_15 ;
	7'h3d :
		TR_262 = TR_15 ;
	7'h3e :
		TR_262 = TR_15 ;
	7'h3f :
		TR_262 = TR_15 ;
	7'h40 :
		TR_262 = TR_15 ;
	7'h41 :
		TR_262 = TR_15 ;
	7'h42 :
		TR_262 = TR_15 ;
	7'h43 :
		TR_262 = TR_15 ;
	7'h44 :
		TR_262 = TR_15 ;
	7'h45 :
		TR_262 = TR_15 ;
	7'h46 :
		TR_262 = TR_15 ;
	7'h47 :
		TR_262 = TR_15 ;
	7'h48 :
		TR_262 = TR_15 ;
	7'h49 :
		TR_262 = TR_15 ;
	7'h4a :
		TR_262 = TR_15 ;
	7'h4b :
		TR_262 = TR_15 ;
	7'h4c :
		TR_262 = TR_15 ;
	7'h4d :
		TR_262 = TR_15 ;
	7'h4e :
		TR_262 = TR_15 ;
	7'h4f :
		TR_262 = TR_15 ;
	7'h50 :
		TR_262 = TR_15 ;
	7'h51 :
		TR_262 = TR_15 ;
	7'h52 :
		TR_262 = TR_15 ;
	7'h53 :
		TR_262 = TR_15 ;
	7'h54 :
		TR_262 = TR_15 ;
	7'h55 :
		TR_262 = TR_15 ;
	7'h56 :
		TR_262 = TR_15 ;
	7'h57 :
		TR_262 = TR_15 ;
	7'h58 :
		TR_262 = TR_15 ;
	7'h59 :
		TR_262 = TR_15 ;
	7'h5a :
		TR_262 = TR_15 ;
	7'h5b :
		TR_262 = TR_15 ;
	7'h5c :
		TR_262 = TR_15 ;
	7'h5d :
		TR_262 = TR_15 ;
	7'h5e :
		TR_262 = TR_15 ;
	7'h5f :
		TR_262 = TR_15 ;
	7'h60 :
		TR_262 = TR_15 ;
	7'h61 :
		TR_262 = TR_15 ;
	7'h62 :
		TR_262 = TR_15 ;
	7'h63 :
		TR_262 = TR_15 ;
	7'h64 :
		TR_262 = TR_15 ;
	7'h65 :
		TR_262 = TR_15 ;
	7'h66 :
		TR_262 = TR_15 ;
	7'h67 :
		TR_262 = TR_15 ;
	7'h68 :
		TR_262 = TR_15 ;
	7'h69 :
		TR_262 = TR_15 ;
	7'h6a :
		TR_262 = TR_15 ;
	7'h6b :
		TR_262 = TR_15 ;
	7'h6c :
		TR_262 = TR_15 ;
	7'h6d :
		TR_262 = TR_15 ;
	7'h6e :
		TR_262 = TR_15 ;
	7'h6f :
		TR_262 = TR_15 ;
	7'h70 :
		TR_262 = TR_15 ;
	7'h71 :
		TR_262 = TR_15 ;
	7'h72 :
		TR_262 = TR_15 ;
	7'h73 :
		TR_262 = TR_15 ;
	7'h74 :
		TR_262 = TR_15 ;
	7'h75 :
		TR_262 = TR_15 ;
	7'h76 :
		TR_262 = TR_15 ;
	7'h77 :
		TR_262 = TR_15 ;
	7'h78 :
		TR_262 = TR_15 ;
	7'h79 :
		TR_262 = TR_15 ;
	7'h7a :
		TR_262 = TR_15 ;
	7'h7b :
		TR_262 = TR_15 ;
	7'h7c :
		TR_262 = TR_15 ;
	7'h7d :
		TR_262 = TR_15 ;
	7'h7e :
		TR_262 = TR_15 ;
	7'h7f :
		TR_262 = TR_15 ;
	default :
		TR_262 = 9'hx ;
	endcase
always @ ( TR_262 or U_173 or sub8u_71ot or U_183 or RG_rl_130 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_3_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h03 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_3_t = ( ( { 9{ M_180 } } & RG_rl_130 )
		| ( { 9{ U_173 } } & TR_262 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_3_en = ( M_180 | RG_rl_3_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_3_en )
		RG_rl_3 <= RG_rl_3_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_16 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_261 = TR_16 ;
	7'h01 :
		TR_261 = TR_16 ;
	7'h02 :
		TR_261 = TR_16 ;
	7'h03 :
		TR_261 = TR_16 ;
	7'h04 :
		TR_261 = 9'h000 ;	// line#=../rle.cpp:80
	7'h05 :
		TR_261 = TR_16 ;
	7'h06 :
		TR_261 = TR_16 ;
	7'h07 :
		TR_261 = TR_16 ;
	7'h08 :
		TR_261 = TR_16 ;
	7'h09 :
		TR_261 = TR_16 ;
	7'h0a :
		TR_261 = TR_16 ;
	7'h0b :
		TR_261 = TR_16 ;
	7'h0c :
		TR_261 = TR_16 ;
	7'h0d :
		TR_261 = TR_16 ;
	7'h0e :
		TR_261 = TR_16 ;
	7'h0f :
		TR_261 = TR_16 ;
	7'h10 :
		TR_261 = TR_16 ;
	7'h11 :
		TR_261 = TR_16 ;
	7'h12 :
		TR_261 = TR_16 ;
	7'h13 :
		TR_261 = TR_16 ;
	7'h14 :
		TR_261 = TR_16 ;
	7'h15 :
		TR_261 = TR_16 ;
	7'h16 :
		TR_261 = TR_16 ;
	7'h17 :
		TR_261 = TR_16 ;
	7'h18 :
		TR_261 = TR_16 ;
	7'h19 :
		TR_261 = TR_16 ;
	7'h1a :
		TR_261 = TR_16 ;
	7'h1b :
		TR_261 = TR_16 ;
	7'h1c :
		TR_261 = TR_16 ;
	7'h1d :
		TR_261 = TR_16 ;
	7'h1e :
		TR_261 = TR_16 ;
	7'h1f :
		TR_261 = TR_16 ;
	7'h20 :
		TR_261 = TR_16 ;
	7'h21 :
		TR_261 = TR_16 ;
	7'h22 :
		TR_261 = TR_16 ;
	7'h23 :
		TR_261 = TR_16 ;
	7'h24 :
		TR_261 = TR_16 ;
	7'h25 :
		TR_261 = TR_16 ;
	7'h26 :
		TR_261 = TR_16 ;
	7'h27 :
		TR_261 = TR_16 ;
	7'h28 :
		TR_261 = TR_16 ;
	7'h29 :
		TR_261 = TR_16 ;
	7'h2a :
		TR_261 = TR_16 ;
	7'h2b :
		TR_261 = TR_16 ;
	7'h2c :
		TR_261 = TR_16 ;
	7'h2d :
		TR_261 = TR_16 ;
	7'h2e :
		TR_261 = TR_16 ;
	7'h2f :
		TR_261 = TR_16 ;
	7'h30 :
		TR_261 = TR_16 ;
	7'h31 :
		TR_261 = TR_16 ;
	7'h32 :
		TR_261 = TR_16 ;
	7'h33 :
		TR_261 = TR_16 ;
	7'h34 :
		TR_261 = TR_16 ;
	7'h35 :
		TR_261 = TR_16 ;
	7'h36 :
		TR_261 = TR_16 ;
	7'h37 :
		TR_261 = TR_16 ;
	7'h38 :
		TR_261 = TR_16 ;
	7'h39 :
		TR_261 = TR_16 ;
	7'h3a :
		TR_261 = TR_16 ;
	7'h3b :
		TR_261 = TR_16 ;
	7'h3c :
		TR_261 = TR_16 ;
	7'h3d :
		TR_261 = TR_16 ;
	7'h3e :
		TR_261 = TR_16 ;
	7'h3f :
		TR_261 = TR_16 ;
	7'h40 :
		TR_261 = TR_16 ;
	7'h41 :
		TR_261 = TR_16 ;
	7'h42 :
		TR_261 = TR_16 ;
	7'h43 :
		TR_261 = TR_16 ;
	7'h44 :
		TR_261 = TR_16 ;
	7'h45 :
		TR_261 = TR_16 ;
	7'h46 :
		TR_261 = TR_16 ;
	7'h47 :
		TR_261 = TR_16 ;
	7'h48 :
		TR_261 = TR_16 ;
	7'h49 :
		TR_261 = TR_16 ;
	7'h4a :
		TR_261 = TR_16 ;
	7'h4b :
		TR_261 = TR_16 ;
	7'h4c :
		TR_261 = TR_16 ;
	7'h4d :
		TR_261 = TR_16 ;
	7'h4e :
		TR_261 = TR_16 ;
	7'h4f :
		TR_261 = TR_16 ;
	7'h50 :
		TR_261 = TR_16 ;
	7'h51 :
		TR_261 = TR_16 ;
	7'h52 :
		TR_261 = TR_16 ;
	7'h53 :
		TR_261 = TR_16 ;
	7'h54 :
		TR_261 = TR_16 ;
	7'h55 :
		TR_261 = TR_16 ;
	7'h56 :
		TR_261 = TR_16 ;
	7'h57 :
		TR_261 = TR_16 ;
	7'h58 :
		TR_261 = TR_16 ;
	7'h59 :
		TR_261 = TR_16 ;
	7'h5a :
		TR_261 = TR_16 ;
	7'h5b :
		TR_261 = TR_16 ;
	7'h5c :
		TR_261 = TR_16 ;
	7'h5d :
		TR_261 = TR_16 ;
	7'h5e :
		TR_261 = TR_16 ;
	7'h5f :
		TR_261 = TR_16 ;
	7'h60 :
		TR_261 = TR_16 ;
	7'h61 :
		TR_261 = TR_16 ;
	7'h62 :
		TR_261 = TR_16 ;
	7'h63 :
		TR_261 = TR_16 ;
	7'h64 :
		TR_261 = TR_16 ;
	7'h65 :
		TR_261 = TR_16 ;
	7'h66 :
		TR_261 = TR_16 ;
	7'h67 :
		TR_261 = TR_16 ;
	7'h68 :
		TR_261 = TR_16 ;
	7'h69 :
		TR_261 = TR_16 ;
	7'h6a :
		TR_261 = TR_16 ;
	7'h6b :
		TR_261 = TR_16 ;
	7'h6c :
		TR_261 = TR_16 ;
	7'h6d :
		TR_261 = TR_16 ;
	7'h6e :
		TR_261 = TR_16 ;
	7'h6f :
		TR_261 = TR_16 ;
	7'h70 :
		TR_261 = TR_16 ;
	7'h71 :
		TR_261 = TR_16 ;
	7'h72 :
		TR_261 = TR_16 ;
	7'h73 :
		TR_261 = TR_16 ;
	7'h74 :
		TR_261 = TR_16 ;
	7'h75 :
		TR_261 = TR_16 ;
	7'h76 :
		TR_261 = TR_16 ;
	7'h77 :
		TR_261 = TR_16 ;
	7'h78 :
		TR_261 = TR_16 ;
	7'h79 :
		TR_261 = TR_16 ;
	7'h7a :
		TR_261 = TR_16 ;
	7'h7b :
		TR_261 = TR_16 ;
	7'h7c :
		TR_261 = TR_16 ;
	7'h7d :
		TR_261 = TR_16 ;
	7'h7e :
		TR_261 = TR_16 ;
	7'h7f :
		TR_261 = TR_16 ;
	default :
		TR_261 = 9'hx ;
	endcase
always @ ( TR_261 or U_173 or sub8u_71ot or U_183 or RG_rl_131 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_4_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h04 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_4_t = ( ( { 9{ M_180 } } & RG_rl_131 )
		| ( { 9{ U_173 } } & TR_261 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_4_en = ( M_180 | RG_rl_4_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_4_en )
		RG_rl_4 <= RG_rl_4_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_17 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_260 = TR_17 ;
	7'h01 :
		TR_260 = TR_17 ;
	7'h02 :
		TR_260 = TR_17 ;
	7'h03 :
		TR_260 = TR_17 ;
	7'h04 :
		TR_260 = TR_17 ;
	7'h05 :
		TR_260 = 9'h000 ;	// line#=../rle.cpp:80
	7'h06 :
		TR_260 = TR_17 ;
	7'h07 :
		TR_260 = TR_17 ;
	7'h08 :
		TR_260 = TR_17 ;
	7'h09 :
		TR_260 = TR_17 ;
	7'h0a :
		TR_260 = TR_17 ;
	7'h0b :
		TR_260 = TR_17 ;
	7'h0c :
		TR_260 = TR_17 ;
	7'h0d :
		TR_260 = TR_17 ;
	7'h0e :
		TR_260 = TR_17 ;
	7'h0f :
		TR_260 = TR_17 ;
	7'h10 :
		TR_260 = TR_17 ;
	7'h11 :
		TR_260 = TR_17 ;
	7'h12 :
		TR_260 = TR_17 ;
	7'h13 :
		TR_260 = TR_17 ;
	7'h14 :
		TR_260 = TR_17 ;
	7'h15 :
		TR_260 = TR_17 ;
	7'h16 :
		TR_260 = TR_17 ;
	7'h17 :
		TR_260 = TR_17 ;
	7'h18 :
		TR_260 = TR_17 ;
	7'h19 :
		TR_260 = TR_17 ;
	7'h1a :
		TR_260 = TR_17 ;
	7'h1b :
		TR_260 = TR_17 ;
	7'h1c :
		TR_260 = TR_17 ;
	7'h1d :
		TR_260 = TR_17 ;
	7'h1e :
		TR_260 = TR_17 ;
	7'h1f :
		TR_260 = TR_17 ;
	7'h20 :
		TR_260 = TR_17 ;
	7'h21 :
		TR_260 = TR_17 ;
	7'h22 :
		TR_260 = TR_17 ;
	7'h23 :
		TR_260 = TR_17 ;
	7'h24 :
		TR_260 = TR_17 ;
	7'h25 :
		TR_260 = TR_17 ;
	7'h26 :
		TR_260 = TR_17 ;
	7'h27 :
		TR_260 = TR_17 ;
	7'h28 :
		TR_260 = TR_17 ;
	7'h29 :
		TR_260 = TR_17 ;
	7'h2a :
		TR_260 = TR_17 ;
	7'h2b :
		TR_260 = TR_17 ;
	7'h2c :
		TR_260 = TR_17 ;
	7'h2d :
		TR_260 = TR_17 ;
	7'h2e :
		TR_260 = TR_17 ;
	7'h2f :
		TR_260 = TR_17 ;
	7'h30 :
		TR_260 = TR_17 ;
	7'h31 :
		TR_260 = TR_17 ;
	7'h32 :
		TR_260 = TR_17 ;
	7'h33 :
		TR_260 = TR_17 ;
	7'h34 :
		TR_260 = TR_17 ;
	7'h35 :
		TR_260 = TR_17 ;
	7'h36 :
		TR_260 = TR_17 ;
	7'h37 :
		TR_260 = TR_17 ;
	7'h38 :
		TR_260 = TR_17 ;
	7'h39 :
		TR_260 = TR_17 ;
	7'h3a :
		TR_260 = TR_17 ;
	7'h3b :
		TR_260 = TR_17 ;
	7'h3c :
		TR_260 = TR_17 ;
	7'h3d :
		TR_260 = TR_17 ;
	7'h3e :
		TR_260 = TR_17 ;
	7'h3f :
		TR_260 = TR_17 ;
	7'h40 :
		TR_260 = TR_17 ;
	7'h41 :
		TR_260 = TR_17 ;
	7'h42 :
		TR_260 = TR_17 ;
	7'h43 :
		TR_260 = TR_17 ;
	7'h44 :
		TR_260 = TR_17 ;
	7'h45 :
		TR_260 = TR_17 ;
	7'h46 :
		TR_260 = TR_17 ;
	7'h47 :
		TR_260 = TR_17 ;
	7'h48 :
		TR_260 = TR_17 ;
	7'h49 :
		TR_260 = TR_17 ;
	7'h4a :
		TR_260 = TR_17 ;
	7'h4b :
		TR_260 = TR_17 ;
	7'h4c :
		TR_260 = TR_17 ;
	7'h4d :
		TR_260 = TR_17 ;
	7'h4e :
		TR_260 = TR_17 ;
	7'h4f :
		TR_260 = TR_17 ;
	7'h50 :
		TR_260 = TR_17 ;
	7'h51 :
		TR_260 = TR_17 ;
	7'h52 :
		TR_260 = TR_17 ;
	7'h53 :
		TR_260 = TR_17 ;
	7'h54 :
		TR_260 = TR_17 ;
	7'h55 :
		TR_260 = TR_17 ;
	7'h56 :
		TR_260 = TR_17 ;
	7'h57 :
		TR_260 = TR_17 ;
	7'h58 :
		TR_260 = TR_17 ;
	7'h59 :
		TR_260 = TR_17 ;
	7'h5a :
		TR_260 = TR_17 ;
	7'h5b :
		TR_260 = TR_17 ;
	7'h5c :
		TR_260 = TR_17 ;
	7'h5d :
		TR_260 = TR_17 ;
	7'h5e :
		TR_260 = TR_17 ;
	7'h5f :
		TR_260 = TR_17 ;
	7'h60 :
		TR_260 = TR_17 ;
	7'h61 :
		TR_260 = TR_17 ;
	7'h62 :
		TR_260 = TR_17 ;
	7'h63 :
		TR_260 = TR_17 ;
	7'h64 :
		TR_260 = TR_17 ;
	7'h65 :
		TR_260 = TR_17 ;
	7'h66 :
		TR_260 = TR_17 ;
	7'h67 :
		TR_260 = TR_17 ;
	7'h68 :
		TR_260 = TR_17 ;
	7'h69 :
		TR_260 = TR_17 ;
	7'h6a :
		TR_260 = TR_17 ;
	7'h6b :
		TR_260 = TR_17 ;
	7'h6c :
		TR_260 = TR_17 ;
	7'h6d :
		TR_260 = TR_17 ;
	7'h6e :
		TR_260 = TR_17 ;
	7'h6f :
		TR_260 = TR_17 ;
	7'h70 :
		TR_260 = TR_17 ;
	7'h71 :
		TR_260 = TR_17 ;
	7'h72 :
		TR_260 = TR_17 ;
	7'h73 :
		TR_260 = TR_17 ;
	7'h74 :
		TR_260 = TR_17 ;
	7'h75 :
		TR_260 = TR_17 ;
	7'h76 :
		TR_260 = TR_17 ;
	7'h77 :
		TR_260 = TR_17 ;
	7'h78 :
		TR_260 = TR_17 ;
	7'h79 :
		TR_260 = TR_17 ;
	7'h7a :
		TR_260 = TR_17 ;
	7'h7b :
		TR_260 = TR_17 ;
	7'h7c :
		TR_260 = TR_17 ;
	7'h7d :
		TR_260 = TR_17 ;
	7'h7e :
		TR_260 = TR_17 ;
	7'h7f :
		TR_260 = TR_17 ;
	default :
		TR_260 = 9'hx ;
	endcase
always @ ( TR_260 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl or U_174 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_5_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h05 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_5_t = ( ( { 9{ U_174 } } & RG_quantized_block_rl )
		| ( { 9{ U_173 } } & TR_260 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_5_en = ( U_174 | RG_rl_5_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_5_en )
		RG_rl_5 <= RG_rl_5_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_18 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_259 = TR_18 ;
	7'h01 :
		TR_259 = TR_18 ;
	7'h02 :
		TR_259 = TR_18 ;
	7'h03 :
		TR_259 = TR_18 ;
	7'h04 :
		TR_259 = TR_18 ;
	7'h05 :
		TR_259 = TR_18 ;
	7'h06 :
		TR_259 = 9'h000 ;	// line#=../rle.cpp:80
	7'h07 :
		TR_259 = TR_18 ;
	7'h08 :
		TR_259 = TR_18 ;
	7'h09 :
		TR_259 = TR_18 ;
	7'h0a :
		TR_259 = TR_18 ;
	7'h0b :
		TR_259 = TR_18 ;
	7'h0c :
		TR_259 = TR_18 ;
	7'h0d :
		TR_259 = TR_18 ;
	7'h0e :
		TR_259 = TR_18 ;
	7'h0f :
		TR_259 = TR_18 ;
	7'h10 :
		TR_259 = TR_18 ;
	7'h11 :
		TR_259 = TR_18 ;
	7'h12 :
		TR_259 = TR_18 ;
	7'h13 :
		TR_259 = TR_18 ;
	7'h14 :
		TR_259 = TR_18 ;
	7'h15 :
		TR_259 = TR_18 ;
	7'h16 :
		TR_259 = TR_18 ;
	7'h17 :
		TR_259 = TR_18 ;
	7'h18 :
		TR_259 = TR_18 ;
	7'h19 :
		TR_259 = TR_18 ;
	7'h1a :
		TR_259 = TR_18 ;
	7'h1b :
		TR_259 = TR_18 ;
	7'h1c :
		TR_259 = TR_18 ;
	7'h1d :
		TR_259 = TR_18 ;
	7'h1e :
		TR_259 = TR_18 ;
	7'h1f :
		TR_259 = TR_18 ;
	7'h20 :
		TR_259 = TR_18 ;
	7'h21 :
		TR_259 = TR_18 ;
	7'h22 :
		TR_259 = TR_18 ;
	7'h23 :
		TR_259 = TR_18 ;
	7'h24 :
		TR_259 = TR_18 ;
	7'h25 :
		TR_259 = TR_18 ;
	7'h26 :
		TR_259 = TR_18 ;
	7'h27 :
		TR_259 = TR_18 ;
	7'h28 :
		TR_259 = TR_18 ;
	7'h29 :
		TR_259 = TR_18 ;
	7'h2a :
		TR_259 = TR_18 ;
	7'h2b :
		TR_259 = TR_18 ;
	7'h2c :
		TR_259 = TR_18 ;
	7'h2d :
		TR_259 = TR_18 ;
	7'h2e :
		TR_259 = TR_18 ;
	7'h2f :
		TR_259 = TR_18 ;
	7'h30 :
		TR_259 = TR_18 ;
	7'h31 :
		TR_259 = TR_18 ;
	7'h32 :
		TR_259 = TR_18 ;
	7'h33 :
		TR_259 = TR_18 ;
	7'h34 :
		TR_259 = TR_18 ;
	7'h35 :
		TR_259 = TR_18 ;
	7'h36 :
		TR_259 = TR_18 ;
	7'h37 :
		TR_259 = TR_18 ;
	7'h38 :
		TR_259 = TR_18 ;
	7'h39 :
		TR_259 = TR_18 ;
	7'h3a :
		TR_259 = TR_18 ;
	7'h3b :
		TR_259 = TR_18 ;
	7'h3c :
		TR_259 = TR_18 ;
	7'h3d :
		TR_259 = TR_18 ;
	7'h3e :
		TR_259 = TR_18 ;
	7'h3f :
		TR_259 = TR_18 ;
	7'h40 :
		TR_259 = TR_18 ;
	7'h41 :
		TR_259 = TR_18 ;
	7'h42 :
		TR_259 = TR_18 ;
	7'h43 :
		TR_259 = TR_18 ;
	7'h44 :
		TR_259 = TR_18 ;
	7'h45 :
		TR_259 = TR_18 ;
	7'h46 :
		TR_259 = TR_18 ;
	7'h47 :
		TR_259 = TR_18 ;
	7'h48 :
		TR_259 = TR_18 ;
	7'h49 :
		TR_259 = TR_18 ;
	7'h4a :
		TR_259 = TR_18 ;
	7'h4b :
		TR_259 = TR_18 ;
	7'h4c :
		TR_259 = TR_18 ;
	7'h4d :
		TR_259 = TR_18 ;
	7'h4e :
		TR_259 = TR_18 ;
	7'h4f :
		TR_259 = TR_18 ;
	7'h50 :
		TR_259 = TR_18 ;
	7'h51 :
		TR_259 = TR_18 ;
	7'h52 :
		TR_259 = TR_18 ;
	7'h53 :
		TR_259 = TR_18 ;
	7'h54 :
		TR_259 = TR_18 ;
	7'h55 :
		TR_259 = TR_18 ;
	7'h56 :
		TR_259 = TR_18 ;
	7'h57 :
		TR_259 = TR_18 ;
	7'h58 :
		TR_259 = TR_18 ;
	7'h59 :
		TR_259 = TR_18 ;
	7'h5a :
		TR_259 = TR_18 ;
	7'h5b :
		TR_259 = TR_18 ;
	7'h5c :
		TR_259 = TR_18 ;
	7'h5d :
		TR_259 = TR_18 ;
	7'h5e :
		TR_259 = TR_18 ;
	7'h5f :
		TR_259 = TR_18 ;
	7'h60 :
		TR_259 = TR_18 ;
	7'h61 :
		TR_259 = TR_18 ;
	7'h62 :
		TR_259 = TR_18 ;
	7'h63 :
		TR_259 = TR_18 ;
	7'h64 :
		TR_259 = TR_18 ;
	7'h65 :
		TR_259 = TR_18 ;
	7'h66 :
		TR_259 = TR_18 ;
	7'h67 :
		TR_259 = TR_18 ;
	7'h68 :
		TR_259 = TR_18 ;
	7'h69 :
		TR_259 = TR_18 ;
	7'h6a :
		TR_259 = TR_18 ;
	7'h6b :
		TR_259 = TR_18 ;
	7'h6c :
		TR_259 = TR_18 ;
	7'h6d :
		TR_259 = TR_18 ;
	7'h6e :
		TR_259 = TR_18 ;
	7'h6f :
		TR_259 = TR_18 ;
	7'h70 :
		TR_259 = TR_18 ;
	7'h71 :
		TR_259 = TR_18 ;
	7'h72 :
		TR_259 = TR_18 ;
	7'h73 :
		TR_259 = TR_18 ;
	7'h74 :
		TR_259 = TR_18 ;
	7'h75 :
		TR_259 = TR_18 ;
	7'h76 :
		TR_259 = TR_18 ;
	7'h77 :
		TR_259 = TR_18 ;
	7'h78 :
		TR_259 = TR_18 ;
	7'h79 :
		TR_259 = TR_18 ;
	7'h7a :
		TR_259 = TR_18 ;
	7'h7b :
		TR_259 = TR_18 ;
	7'h7c :
		TR_259 = TR_18 ;
	7'h7d :
		TR_259 = TR_18 ;
	7'h7e :
		TR_259 = TR_18 ;
	7'h7f :
		TR_259 = TR_18 ;
	default :
		TR_259 = 9'hx ;
	endcase
always @ ( TR_259 or U_173 or sub8u_71ot or U_183 or RG_rl_132 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_6_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h06 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_6_t = ( ( { 9{ M_180 } } & RG_rl_132 )
		| ( { 9{ U_173 } } & TR_259 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_6_en = ( M_180 | RG_rl_6_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_6_en )
		RG_rl_6 <= RG_rl_6_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_19 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_258 = TR_19 ;
	7'h01 :
		TR_258 = TR_19 ;
	7'h02 :
		TR_258 = TR_19 ;
	7'h03 :
		TR_258 = TR_19 ;
	7'h04 :
		TR_258 = TR_19 ;
	7'h05 :
		TR_258 = TR_19 ;
	7'h06 :
		TR_258 = TR_19 ;
	7'h07 :
		TR_258 = 9'h000 ;	// line#=../rle.cpp:80
	7'h08 :
		TR_258 = TR_19 ;
	7'h09 :
		TR_258 = TR_19 ;
	7'h0a :
		TR_258 = TR_19 ;
	7'h0b :
		TR_258 = TR_19 ;
	7'h0c :
		TR_258 = TR_19 ;
	7'h0d :
		TR_258 = TR_19 ;
	7'h0e :
		TR_258 = TR_19 ;
	7'h0f :
		TR_258 = TR_19 ;
	7'h10 :
		TR_258 = TR_19 ;
	7'h11 :
		TR_258 = TR_19 ;
	7'h12 :
		TR_258 = TR_19 ;
	7'h13 :
		TR_258 = TR_19 ;
	7'h14 :
		TR_258 = TR_19 ;
	7'h15 :
		TR_258 = TR_19 ;
	7'h16 :
		TR_258 = TR_19 ;
	7'h17 :
		TR_258 = TR_19 ;
	7'h18 :
		TR_258 = TR_19 ;
	7'h19 :
		TR_258 = TR_19 ;
	7'h1a :
		TR_258 = TR_19 ;
	7'h1b :
		TR_258 = TR_19 ;
	7'h1c :
		TR_258 = TR_19 ;
	7'h1d :
		TR_258 = TR_19 ;
	7'h1e :
		TR_258 = TR_19 ;
	7'h1f :
		TR_258 = TR_19 ;
	7'h20 :
		TR_258 = TR_19 ;
	7'h21 :
		TR_258 = TR_19 ;
	7'h22 :
		TR_258 = TR_19 ;
	7'h23 :
		TR_258 = TR_19 ;
	7'h24 :
		TR_258 = TR_19 ;
	7'h25 :
		TR_258 = TR_19 ;
	7'h26 :
		TR_258 = TR_19 ;
	7'h27 :
		TR_258 = TR_19 ;
	7'h28 :
		TR_258 = TR_19 ;
	7'h29 :
		TR_258 = TR_19 ;
	7'h2a :
		TR_258 = TR_19 ;
	7'h2b :
		TR_258 = TR_19 ;
	7'h2c :
		TR_258 = TR_19 ;
	7'h2d :
		TR_258 = TR_19 ;
	7'h2e :
		TR_258 = TR_19 ;
	7'h2f :
		TR_258 = TR_19 ;
	7'h30 :
		TR_258 = TR_19 ;
	7'h31 :
		TR_258 = TR_19 ;
	7'h32 :
		TR_258 = TR_19 ;
	7'h33 :
		TR_258 = TR_19 ;
	7'h34 :
		TR_258 = TR_19 ;
	7'h35 :
		TR_258 = TR_19 ;
	7'h36 :
		TR_258 = TR_19 ;
	7'h37 :
		TR_258 = TR_19 ;
	7'h38 :
		TR_258 = TR_19 ;
	7'h39 :
		TR_258 = TR_19 ;
	7'h3a :
		TR_258 = TR_19 ;
	7'h3b :
		TR_258 = TR_19 ;
	7'h3c :
		TR_258 = TR_19 ;
	7'h3d :
		TR_258 = TR_19 ;
	7'h3e :
		TR_258 = TR_19 ;
	7'h3f :
		TR_258 = TR_19 ;
	7'h40 :
		TR_258 = TR_19 ;
	7'h41 :
		TR_258 = TR_19 ;
	7'h42 :
		TR_258 = TR_19 ;
	7'h43 :
		TR_258 = TR_19 ;
	7'h44 :
		TR_258 = TR_19 ;
	7'h45 :
		TR_258 = TR_19 ;
	7'h46 :
		TR_258 = TR_19 ;
	7'h47 :
		TR_258 = TR_19 ;
	7'h48 :
		TR_258 = TR_19 ;
	7'h49 :
		TR_258 = TR_19 ;
	7'h4a :
		TR_258 = TR_19 ;
	7'h4b :
		TR_258 = TR_19 ;
	7'h4c :
		TR_258 = TR_19 ;
	7'h4d :
		TR_258 = TR_19 ;
	7'h4e :
		TR_258 = TR_19 ;
	7'h4f :
		TR_258 = TR_19 ;
	7'h50 :
		TR_258 = TR_19 ;
	7'h51 :
		TR_258 = TR_19 ;
	7'h52 :
		TR_258 = TR_19 ;
	7'h53 :
		TR_258 = TR_19 ;
	7'h54 :
		TR_258 = TR_19 ;
	7'h55 :
		TR_258 = TR_19 ;
	7'h56 :
		TR_258 = TR_19 ;
	7'h57 :
		TR_258 = TR_19 ;
	7'h58 :
		TR_258 = TR_19 ;
	7'h59 :
		TR_258 = TR_19 ;
	7'h5a :
		TR_258 = TR_19 ;
	7'h5b :
		TR_258 = TR_19 ;
	7'h5c :
		TR_258 = TR_19 ;
	7'h5d :
		TR_258 = TR_19 ;
	7'h5e :
		TR_258 = TR_19 ;
	7'h5f :
		TR_258 = TR_19 ;
	7'h60 :
		TR_258 = TR_19 ;
	7'h61 :
		TR_258 = TR_19 ;
	7'h62 :
		TR_258 = TR_19 ;
	7'h63 :
		TR_258 = TR_19 ;
	7'h64 :
		TR_258 = TR_19 ;
	7'h65 :
		TR_258 = TR_19 ;
	7'h66 :
		TR_258 = TR_19 ;
	7'h67 :
		TR_258 = TR_19 ;
	7'h68 :
		TR_258 = TR_19 ;
	7'h69 :
		TR_258 = TR_19 ;
	7'h6a :
		TR_258 = TR_19 ;
	7'h6b :
		TR_258 = TR_19 ;
	7'h6c :
		TR_258 = TR_19 ;
	7'h6d :
		TR_258 = TR_19 ;
	7'h6e :
		TR_258 = TR_19 ;
	7'h6f :
		TR_258 = TR_19 ;
	7'h70 :
		TR_258 = TR_19 ;
	7'h71 :
		TR_258 = TR_19 ;
	7'h72 :
		TR_258 = TR_19 ;
	7'h73 :
		TR_258 = TR_19 ;
	7'h74 :
		TR_258 = TR_19 ;
	7'h75 :
		TR_258 = TR_19 ;
	7'h76 :
		TR_258 = TR_19 ;
	7'h77 :
		TR_258 = TR_19 ;
	7'h78 :
		TR_258 = TR_19 ;
	7'h79 :
		TR_258 = TR_19 ;
	7'h7a :
		TR_258 = TR_19 ;
	7'h7b :
		TR_258 = TR_19 ;
	7'h7c :
		TR_258 = TR_19 ;
	7'h7d :
		TR_258 = TR_19 ;
	7'h7e :
		TR_258 = TR_19 ;
	7'h7f :
		TR_258 = TR_19 ;
	default :
		TR_258 = 9'hx ;
	endcase
always @ ( TR_258 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_1 or 
	U_174 or RG_rl_132 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_7_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h07 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_7_t = ( ( { 9{ ST1_03d } } & RG_rl_132 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_1 )
		| ( { 9{ U_173 } } & TR_258 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_7_en = ( ST1_03d | U_174 | RG_rl_7_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_7_en )
		RG_rl_7 <= RG_rl_7_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_20 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_257 = TR_20 ;
	7'h01 :
		TR_257 = TR_20 ;
	7'h02 :
		TR_257 = TR_20 ;
	7'h03 :
		TR_257 = TR_20 ;
	7'h04 :
		TR_257 = TR_20 ;
	7'h05 :
		TR_257 = TR_20 ;
	7'h06 :
		TR_257 = TR_20 ;
	7'h07 :
		TR_257 = TR_20 ;
	7'h08 :
		TR_257 = 9'h000 ;	// line#=../rle.cpp:80
	7'h09 :
		TR_257 = TR_20 ;
	7'h0a :
		TR_257 = TR_20 ;
	7'h0b :
		TR_257 = TR_20 ;
	7'h0c :
		TR_257 = TR_20 ;
	7'h0d :
		TR_257 = TR_20 ;
	7'h0e :
		TR_257 = TR_20 ;
	7'h0f :
		TR_257 = TR_20 ;
	7'h10 :
		TR_257 = TR_20 ;
	7'h11 :
		TR_257 = TR_20 ;
	7'h12 :
		TR_257 = TR_20 ;
	7'h13 :
		TR_257 = TR_20 ;
	7'h14 :
		TR_257 = TR_20 ;
	7'h15 :
		TR_257 = TR_20 ;
	7'h16 :
		TR_257 = TR_20 ;
	7'h17 :
		TR_257 = TR_20 ;
	7'h18 :
		TR_257 = TR_20 ;
	7'h19 :
		TR_257 = TR_20 ;
	7'h1a :
		TR_257 = TR_20 ;
	7'h1b :
		TR_257 = TR_20 ;
	7'h1c :
		TR_257 = TR_20 ;
	7'h1d :
		TR_257 = TR_20 ;
	7'h1e :
		TR_257 = TR_20 ;
	7'h1f :
		TR_257 = TR_20 ;
	7'h20 :
		TR_257 = TR_20 ;
	7'h21 :
		TR_257 = TR_20 ;
	7'h22 :
		TR_257 = TR_20 ;
	7'h23 :
		TR_257 = TR_20 ;
	7'h24 :
		TR_257 = TR_20 ;
	7'h25 :
		TR_257 = TR_20 ;
	7'h26 :
		TR_257 = TR_20 ;
	7'h27 :
		TR_257 = TR_20 ;
	7'h28 :
		TR_257 = TR_20 ;
	7'h29 :
		TR_257 = TR_20 ;
	7'h2a :
		TR_257 = TR_20 ;
	7'h2b :
		TR_257 = TR_20 ;
	7'h2c :
		TR_257 = TR_20 ;
	7'h2d :
		TR_257 = TR_20 ;
	7'h2e :
		TR_257 = TR_20 ;
	7'h2f :
		TR_257 = TR_20 ;
	7'h30 :
		TR_257 = TR_20 ;
	7'h31 :
		TR_257 = TR_20 ;
	7'h32 :
		TR_257 = TR_20 ;
	7'h33 :
		TR_257 = TR_20 ;
	7'h34 :
		TR_257 = TR_20 ;
	7'h35 :
		TR_257 = TR_20 ;
	7'h36 :
		TR_257 = TR_20 ;
	7'h37 :
		TR_257 = TR_20 ;
	7'h38 :
		TR_257 = TR_20 ;
	7'h39 :
		TR_257 = TR_20 ;
	7'h3a :
		TR_257 = TR_20 ;
	7'h3b :
		TR_257 = TR_20 ;
	7'h3c :
		TR_257 = TR_20 ;
	7'h3d :
		TR_257 = TR_20 ;
	7'h3e :
		TR_257 = TR_20 ;
	7'h3f :
		TR_257 = TR_20 ;
	7'h40 :
		TR_257 = TR_20 ;
	7'h41 :
		TR_257 = TR_20 ;
	7'h42 :
		TR_257 = TR_20 ;
	7'h43 :
		TR_257 = TR_20 ;
	7'h44 :
		TR_257 = TR_20 ;
	7'h45 :
		TR_257 = TR_20 ;
	7'h46 :
		TR_257 = TR_20 ;
	7'h47 :
		TR_257 = TR_20 ;
	7'h48 :
		TR_257 = TR_20 ;
	7'h49 :
		TR_257 = TR_20 ;
	7'h4a :
		TR_257 = TR_20 ;
	7'h4b :
		TR_257 = TR_20 ;
	7'h4c :
		TR_257 = TR_20 ;
	7'h4d :
		TR_257 = TR_20 ;
	7'h4e :
		TR_257 = TR_20 ;
	7'h4f :
		TR_257 = TR_20 ;
	7'h50 :
		TR_257 = TR_20 ;
	7'h51 :
		TR_257 = TR_20 ;
	7'h52 :
		TR_257 = TR_20 ;
	7'h53 :
		TR_257 = TR_20 ;
	7'h54 :
		TR_257 = TR_20 ;
	7'h55 :
		TR_257 = TR_20 ;
	7'h56 :
		TR_257 = TR_20 ;
	7'h57 :
		TR_257 = TR_20 ;
	7'h58 :
		TR_257 = TR_20 ;
	7'h59 :
		TR_257 = TR_20 ;
	7'h5a :
		TR_257 = TR_20 ;
	7'h5b :
		TR_257 = TR_20 ;
	7'h5c :
		TR_257 = TR_20 ;
	7'h5d :
		TR_257 = TR_20 ;
	7'h5e :
		TR_257 = TR_20 ;
	7'h5f :
		TR_257 = TR_20 ;
	7'h60 :
		TR_257 = TR_20 ;
	7'h61 :
		TR_257 = TR_20 ;
	7'h62 :
		TR_257 = TR_20 ;
	7'h63 :
		TR_257 = TR_20 ;
	7'h64 :
		TR_257 = TR_20 ;
	7'h65 :
		TR_257 = TR_20 ;
	7'h66 :
		TR_257 = TR_20 ;
	7'h67 :
		TR_257 = TR_20 ;
	7'h68 :
		TR_257 = TR_20 ;
	7'h69 :
		TR_257 = TR_20 ;
	7'h6a :
		TR_257 = TR_20 ;
	7'h6b :
		TR_257 = TR_20 ;
	7'h6c :
		TR_257 = TR_20 ;
	7'h6d :
		TR_257 = TR_20 ;
	7'h6e :
		TR_257 = TR_20 ;
	7'h6f :
		TR_257 = TR_20 ;
	7'h70 :
		TR_257 = TR_20 ;
	7'h71 :
		TR_257 = TR_20 ;
	7'h72 :
		TR_257 = TR_20 ;
	7'h73 :
		TR_257 = TR_20 ;
	7'h74 :
		TR_257 = TR_20 ;
	7'h75 :
		TR_257 = TR_20 ;
	7'h76 :
		TR_257 = TR_20 ;
	7'h77 :
		TR_257 = TR_20 ;
	7'h78 :
		TR_257 = TR_20 ;
	7'h79 :
		TR_257 = TR_20 ;
	7'h7a :
		TR_257 = TR_20 ;
	7'h7b :
		TR_257 = TR_20 ;
	7'h7c :
		TR_257 = TR_20 ;
	7'h7d :
		TR_257 = TR_20 ;
	7'h7e :
		TR_257 = TR_20 ;
	7'h7f :
		TR_257 = TR_20 ;
	default :
		TR_257 = 9'hx ;
	endcase
always @ ( TR_257 or U_173 or sub8u_71ot or U_183 or RG_rl_133 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_8_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h08 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_8_t = ( ( { 9{ M_180 } } & RG_rl_133 )
		| ( { 9{ U_173 } } & TR_257 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_8_en = ( M_180 | RG_rl_8_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_8_en )
		RG_rl_8 <= RG_rl_8_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_21 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_256 = TR_21 ;
	7'h01 :
		TR_256 = TR_21 ;
	7'h02 :
		TR_256 = TR_21 ;
	7'h03 :
		TR_256 = TR_21 ;
	7'h04 :
		TR_256 = TR_21 ;
	7'h05 :
		TR_256 = TR_21 ;
	7'h06 :
		TR_256 = TR_21 ;
	7'h07 :
		TR_256 = TR_21 ;
	7'h08 :
		TR_256 = TR_21 ;
	7'h09 :
		TR_256 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0a :
		TR_256 = TR_21 ;
	7'h0b :
		TR_256 = TR_21 ;
	7'h0c :
		TR_256 = TR_21 ;
	7'h0d :
		TR_256 = TR_21 ;
	7'h0e :
		TR_256 = TR_21 ;
	7'h0f :
		TR_256 = TR_21 ;
	7'h10 :
		TR_256 = TR_21 ;
	7'h11 :
		TR_256 = TR_21 ;
	7'h12 :
		TR_256 = TR_21 ;
	7'h13 :
		TR_256 = TR_21 ;
	7'h14 :
		TR_256 = TR_21 ;
	7'h15 :
		TR_256 = TR_21 ;
	7'h16 :
		TR_256 = TR_21 ;
	7'h17 :
		TR_256 = TR_21 ;
	7'h18 :
		TR_256 = TR_21 ;
	7'h19 :
		TR_256 = TR_21 ;
	7'h1a :
		TR_256 = TR_21 ;
	7'h1b :
		TR_256 = TR_21 ;
	7'h1c :
		TR_256 = TR_21 ;
	7'h1d :
		TR_256 = TR_21 ;
	7'h1e :
		TR_256 = TR_21 ;
	7'h1f :
		TR_256 = TR_21 ;
	7'h20 :
		TR_256 = TR_21 ;
	7'h21 :
		TR_256 = TR_21 ;
	7'h22 :
		TR_256 = TR_21 ;
	7'h23 :
		TR_256 = TR_21 ;
	7'h24 :
		TR_256 = TR_21 ;
	7'h25 :
		TR_256 = TR_21 ;
	7'h26 :
		TR_256 = TR_21 ;
	7'h27 :
		TR_256 = TR_21 ;
	7'h28 :
		TR_256 = TR_21 ;
	7'h29 :
		TR_256 = TR_21 ;
	7'h2a :
		TR_256 = TR_21 ;
	7'h2b :
		TR_256 = TR_21 ;
	7'h2c :
		TR_256 = TR_21 ;
	7'h2d :
		TR_256 = TR_21 ;
	7'h2e :
		TR_256 = TR_21 ;
	7'h2f :
		TR_256 = TR_21 ;
	7'h30 :
		TR_256 = TR_21 ;
	7'h31 :
		TR_256 = TR_21 ;
	7'h32 :
		TR_256 = TR_21 ;
	7'h33 :
		TR_256 = TR_21 ;
	7'h34 :
		TR_256 = TR_21 ;
	7'h35 :
		TR_256 = TR_21 ;
	7'h36 :
		TR_256 = TR_21 ;
	7'h37 :
		TR_256 = TR_21 ;
	7'h38 :
		TR_256 = TR_21 ;
	7'h39 :
		TR_256 = TR_21 ;
	7'h3a :
		TR_256 = TR_21 ;
	7'h3b :
		TR_256 = TR_21 ;
	7'h3c :
		TR_256 = TR_21 ;
	7'h3d :
		TR_256 = TR_21 ;
	7'h3e :
		TR_256 = TR_21 ;
	7'h3f :
		TR_256 = TR_21 ;
	7'h40 :
		TR_256 = TR_21 ;
	7'h41 :
		TR_256 = TR_21 ;
	7'h42 :
		TR_256 = TR_21 ;
	7'h43 :
		TR_256 = TR_21 ;
	7'h44 :
		TR_256 = TR_21 ;
	7'h45 :
		TR_256 = TR_21 ;
	7'h46 :
		TR_256 = TR_21 ;
	7'h47 :
		TR_256 = TR_21 ;
	7'h48 :
		TR_256 = TR_21 ;
	7'h49 :
		TR_256 = TR_21 ;
	7'h4a :
		TR_256 = TR_21 ;
	7'h4b :
		TR_256 = TR_21 ;
	7'h4c :
		TR_256 = TR_21 ;
	7'h4d :
		TR_256 = TR_21 ;
	7'h4e :
		TR_256 = TR_21 ;
	7'h4f :
		TR_256 = TR_21 ;
	7'h50 :
		TR_256 = TR_21 ;
	7'h51 :
		TR_256 = TR_21 ;
	7'h52 :
		TR_256 = TR_21 ;
	7'h53 :
		TR_256 = TR_21 ;
	7'h54 :
		TR_256 = TR_21 ;
	7'h55 :
		TR_256 = TR_21 ;
	7'h56 :
		TR_256 = TR_21 ;
	7'h57 :
		TR_256 = TR_21 ;
	7'h58 :
		TR_256 = TR_21 ;
	7'h59 :
		TR_256 = TR_21 ;
	7'h5a :
		TR_256 = TR_21 ;
	7'h5b :
		TR_256 = TR_21 ;
	7'h5c :
		TR_256 = TR_21 ;
	7'h5d :
		TR_256 = TR_21 ;
	7'h5e :
		TR_256 = TR_21 ;
	7'h5f :
		TR_256 = TR_21 ;
	7'h60 :
		TR_256 = TR_21 ;
	7'h61 :
		TR_256 = TR_21 ;
	7'h62 :
		TR_256 = TR_21 ;
	7'h63 :
		TR_256 = TR_21 ;
	7'h64 :
		TR_256 = TR_21 ;
	7'h65 :
		TR_256 = TR_21 ;
	7'h66 :
		TR_256 = TR_21 ;
	7'h67 :
		TR_256 = TR_21 ;
	7'h68 :
		TR_256 = TR_21 ;
	7'h69 :
		TR_256 = TR_21 ;
	7'h6a :
		TR_256 = TR_21 ;
	7'h6b :
		TR_256 = TR_21 ;
	7'h6c :
		TR_256 = TR_21 ;
	7'h6d :
		TR_256 = TR_21 ;
	7'h6e :
		TR_256 = TR_21 ;
	7'h6f :
		TR_256 = TR_21 ;
	7'h70 :
		TR_256 = TR_21 ;
	7'h71 :
		TR_256 = TR_21 ;
	7'h72 :
		TR_256 = TR_21 ;
	7'h73 :
		TR_256 = TR_21 ;
	7'h74 :
		TR_256 = TR_21 ;
	7'h75 :
		TR_256 = TR_21 ;
	7'h76 :
		TR_256 = TR_21 ;
	7'h77 :
		TR_256 = TR_21 ;
	7'h78 :
		TR_256 = TR_21 ;
	7'h79 :
		TR_256 = TR_21 ;
	7'h7a :
		TR_256 = TR_21 ;
	7'h7b :
		TR_256 = TR_21 ;
	7'h7c :
		TR_256 = TR_21 ;
	7'h7d :
		TR_256 = TR_21 ;
	7'h7e :
		TR_256 = TR_21 ;
	7'h7f :
		TR_256 = TR_21 ;
	default :
		TR_256 = 9'hx ;
	endcase
always @ ( TR_256 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_2 or 
	U_174 or RG_rl_133 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_9_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h09 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_9_t = ( ( { 9{ ST1_03d } } & RG_rl_133 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_2 )
		| ( { 9{ U_173 } } & TR_256 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_9_en = ( ST1_03d | U_174 | RG_rl_9_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_9_en )
		RG_rl_9 <= RG_rl_9_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_22 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_255 = TR_22 ;
	7'h01 :
		TR_255 = TR_22 ;
	7'h02 :
		TR_255 = TR_22 ;
	7'h03 :
		TR_255 = TR_22 ;
	7'h04 :
		TR_255 = TR_22 ;
	7'h05 :
		TR_255 = TR_22 ;
	7'h06 :
		TR_255 = TR_22 ;
	7'h07 :
		TR_255 = TR_22 ;
	7'h08 :
		TR_255 = TR_22 ;
	7'h09 :
		TR_255 = TR_22 ;
	7'h0a :
		TR_255 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0b :
		TR_255 = TR_22 ;
	7'h0c :
		TR_255 = TR_22 ;
	7'h0d :
		TR_255 = TR_22 ;
	7'h0e :
		TR_255 = TR_22 ;
	7'h0f :
		TR_255 = TR_22 ;
	7'h10 :
		TR_255 = TR_22 ;
	7'h11 :
		TR_255 = TR_22 ;
	7'h12 :
		TR_255 = TR_22 ;
	7'h13 :
		TR_255 = TR_22 ;
	7'h14 :
		TR_255 = TR_22 ;
	7'h15 :
		TR_255 = TR_22 ;
	7'h16 :
		TR_255 = TR_22 ;
	7'h17 :
		TR_255 = TR_22 ;
	7'h18 :
		TR_255 = TR_22 ;
	7'h19 :
		TR_255 = TR_22 ;
	7'h1a :
		TR_255 = TR_22 ;
	7'h1b :
		TR_255 = TR_22 ;
	7'h1c :
		TR_255 = TR_22 ;
	7'h1d :
		TR_255 = TR_22 ;
	7'h1e :
		TR_255 = TR_22 ;
	7'h1f :
		TR_255 = TR_22 ;
	7'h20 :
		TR_255 = TR_22 ;
	7'h21 :
		TR_255 = TR_22 ;
	7'h22 :
		TR_255 = TR_22 ;
	7'h23 :
		TR_255 = TR_22 ;
	7'h24 :
		TR_255 = TR_22 ;
	7'h25 :
		TR_255 = TR_22 ;
	7'h26 :
		TR_255 = TR_22 ;
	7'h27 :
		TR_255 = TR_22 ;
	7'h28 :
		TR_255 = TR_22 ;
	7'h29 :
		TR_255 = TR_22 ;
	7'h2a :
		TR_255 = TR_22 ;
	7'h2b :
		TR_255 = TR_22 ;
	7'h2c :
		TR_255 = TR_22 ;
	7'h2d :
		TR_255 = TR_22 ;
	7'h2e :
		TR_255 = TR_22 ;
	7'h2f :
		TR_255 = TR_22 ;
	7'h30 :
		TR_255 = TR_22 ;
	7'h31 :
		TR_255 = TR_22 ;
	7'h32 :
		TR_255 = TR_22 ;
	7'h33 :
		TR_255 = TR_22 ;
	7'h34 :
		TR_255 = TR_22 ;
	7'h35 :
		TR_255 = TR_22 ;
	7'h36 :
		TR_255 = TR_22 ;
	7'h37 :
		TR_255 = TR_22 ;
	7'h38 :
		TR_255 = TR_22 ;
	7'h39 :
		TR_255 = TR_22 ;
	7'h3a :
		TR_255 = TR_22 ;
	7'h3b :
		TR_255 = TR_22 ;
	7'h3c :
		TR_255 = TR_22 ;
	7'h3d :
		TR_255 = TR_22 ;
	7'h3e :
		TR_255 = TR_22 ;
	7'h3f :
		TR_255 = TR_22 ;
	7'h40 :
		TR_255 = TR_22 ;
	7'h41 :
		TR_255 = TR_22 ;
	7'h42 :
		TR_255 = TR_22 ;
	7'h43 :
		TR_255 = TR_22 ;
	7'h44 :
		TR_255 = TR_22 ;
	7'h45 :
		TR_255 = TR_22 ;
	7'h46 :
		TR_255 = TR_22 ;
	7'h47 :
		TR_255 = TR_22 ;
	7'h48 :
		TR_255 = TR_22 ;
	7'h49 :
		TR_255 = TR_22 ;
	7'h4a :
		TR_255 = TR_22 ;
	7'h4b :
		TR_255 = TR_22 ;
	7'h4c :
		TR_255 = TR_22 ;
	7'h4d :
		TR_255 = TR_22 ;
	7'h4e :
		TR_255 = TR_22 ;
	7'h4f :
		TR_255 = TR_22 ;
	7'h50 :
		TR_255 = TR_22 ;
	7'h51 :
		TR_255 = TR_22 ;
	7'h52 :
		TR_255 = TR_22 ;
	7'h53 :
		TR_255 = TR_22 ;
	7'h54 :
		TR_255 = TR_22 ;
	7'h55 :
		TR_255 = TR_22 ;
	7'h56 :
		TR_255 = TR_22 ;
	7'h57 :
		TR_255 = TR_22 ;
	7'h58 :
		TR_255 = TR_22 ;
	7'h59 :
		TR_255 = TR_22 ;
	7'h5a :
		TR_255 = TR_22 ;
	7'h5b :
		TR_255 = TR_22 ;
	7'h5c :
		TR_255 = TR_22 ;
	7'h5d :
		TR_255 = TR_22 ;
	7'h5e :
		TR_255 = TR_22 ;
	7'h5f :
		TR_255 = TR_22 ;
	7'h60 :
		TR_255 = TR_22 ;
	7'h61 :
		TR_255 = TR_22 ;
	7'h62 :
		TR_255 = TR_22 ;
	7'h63 :
		TR_255 = TR_22 ;
	7'h64 :
		TR_255 = TR_22 ;
	7'h65 :
		TR_255 = TR_22 ;
	7'h66 :
		TR_255 = TR_22 ;
	7'h67 :
		TR_255 = TR_22 ;
	7'h68 :
		TR_255 = TR_22 ;
	7'h69 :
		TR_255 = TR_22 ;
	7'h6a :
		TR_255 = TR_22 ;
	7'h6b :
		TR_255 = TR_22 ;
	7'h6c :
		TR_255 = TR_22 ;
	7'h6d :
		TR_255 = TR_22 ;
	7'h6e :
		TR_255 = TR_22 ;
	7'h6f :
		TR_255 = TR_22 ;
	7'h70 :
		TR_255 = TR_22 ;
	7'h71 :
		TR_255 = TR_22 ;
	7'h72 :
		TR_255 = TR_22 ;
	7'h73 :
		TR_255 = TR_22 ;
	7'h74 :
		TR_255 = TR_22 ;
	7'h75 :
		TR_255 = TR_22 ;
	7'h76 :
		TR_255 = TR_22 ;
	7'h77 :
		TR_255 = TR_22 ;
	7'h78 :
		TR_255 = TR_22 ;
	7'h79 :
		TR_255 = TR_22 ;
	7'h7a :
		TR_255 = TR_22 ;
	7'h7b :
		TR_255 = TR_22 ;
	7'h7c :
		TR_255 = TR_22 ;
	7'h7d :
		TR_255 = TR_22 ;
	7'h7e :
		TR_255 = TR_22 ;
	7'h7f :
		TR_255 = TR_22 ;
	default :
		TR_255 = 9'hx ;
	endcase
always @ ( TR_255 or U_173 or sub8u_71ot or U_183 or RG_rl_134 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_10_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h0a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_10_t = ( ( { 9{ M_180 } } & RG_rl_134 )
		| ( { 9{ U_173 } } & TR_255 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_10_en = ( M_180 | RG_rl_10_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_10_en )
		RG_rl_10 <= RG_rl_10_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_23 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_254 = TR_23 ;
	7'h01 :
		TR_254 = TR_23 ;
	7'h02 :
		TR_254 = TR_23 ;
	7'h03 :
		TR_254 = TR_23 ;
	7'h04 :
		TR_254 = TR_23 ;
	7'h05 :
		TR_254 = TR_23 ;
	7'h06 :
		TR_254 = TR_23 ;
	7'h07 :
		TR_254 = TR_23 ;
	7'h08 :
		TR_254 = TR_23 ;
	7'h09 :
		TR_254 = TR_23 ;
	7'h0a :
		TR_254 = TR_23 ;
	7'h0b :
		TR_254 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0c :
		TR_254 = TR_23 ;
	7'h0d :
		TR_254 = TR_23 ;
	7'h0e :
		TR_254 = TR_23 ;
	7'h0f :
		TR_254 = TR_23 ;
	7'h10 :
		TR_254 = TR_23 ;
	7'h11 :
		TR_254 = TR_23 ;
	7'h12 :
		TR_254 = TR_23 ;
	7'h13 :
		TR_254 = TR_23 ;
	7'h14 :
		TR_254 = TR_23 ;
	7'h15 :
		TR_254 = TR_23 ;
	7'h16 :
		TR_254 = TR_23 ;
	7'h17 :
		TR_254 = TR_23 ;
	7'h18 :
		TR_254 = TR_23 ;
	7'h19 :
		TR_254 = TR_23 ;
	7'h1a :
		TR_254 = TR_23 ;
	7'h1b :
		TR_254 = TR_23 ;
	7'h1c :
		TR_254 = TR_23 ;
	7'h1d :
		TR_254 = TR_23 ;
	7'h1e :
		TR_254 = TR_23 ;
	7'h1f :
		TR_254 = TR_23 ;
	7'h20 :
		TR_254 = TR_23 ;
	7'h21 :
		TR_254 = TR_23 ;
	7'h22 :
		TR_254 = TR_23 ;
	7'h23 :
		TR_254 = TR_23 ;
	7'h24 :
		TR_254 = TR_23 ;
	7'h25 :
		TR_254 = TR_23 ;
	7'h26 :
		TR_254 = TR_23 ;
	7'h27 :
		TR_254 = TR_23 ;
	7'h28 :
		TR_254 = TR_23 ;
	7'h29 :
		TR_254 = TR_23 ;
	7'h2a :
		TR_254 = TR_23 ;
	7'h2b :
		TR_254 = TR_23 ;
	7'h2c :
		TR_254 = TR_23 ;
	7'h2d :
		TR_254 = TR_23 ;
	7'h2e :
		TR_254 = TR_23 ;
	7'h2f :
		TR_254 = TR_23 ;
	7'h30 :
		TR_254 = TR_23 ;
	7'h31 :
		TR_254 = TR_23 ;
	7'h32 :
		TR_254 = TR_23 ;
	7'h33 :
		TR_254 = TR_23 ;
	7'h34 :
		TR_254 = TR_23 ;
	7'h35 :
		TR_254 = TR_23 ;
	7'h36 :
		TR_254 = TR_23 ;
	7'h37 :
		TR_254 = TR_23 ;
	7'h38 :
		TR_254 = TR_23 ;
	7'h39 :
		TR_254 = TR_23 ;
	7'h3a :
		TR_254 = TR_23 ;
	7'h3b :
		TR_254 = TR_23 ;
	7'h3c :
		TR_254 = TR_23 ;
	7'h3d :
		TR_254 = TR_23 ;
	7'h3e :
		TR_254 = TR_23 ;
	7'h3f :
		TR_254 = TR_23 ;
	7'h40 :
		TR_254 = TR_23 ;
	7'h41 :
		TR_254 = TR_23 ;
	7'h42 :
		TR_254 = TR_23 ;
	7'h43 :
		TR_254 = TR_23 ;
	7'h44 :
		TR_254 = TR_23 ;
	7'h45 :
		TR_254 = TR_23 ;
	7'h46 :
		TR_254 = TR_23 ;
	7'h47 :
		TR_254 = TR_23 ;
	7'h48 :
		TR_254 = TR_23 ;
	7'h49 :
		TR_254 = TR_23 ;
	7'h4a :
		TR_254 = TR_23 ;
	7'h4b :
		TR_254 = TR_23 ;
	7'h4c :
		TR_254 = TR_23 ;
	7'h4d :
		TR_254 = TR_23 ;
	7'h4e :
		TR_254 = TR_23 ;
	7'h4f :
		TR_254 = TR_23 ;
	7'h50 :
		TR_254 = TR_23 ;
	7'h51 :
		TR_254 = TR_23 ;
	7'h52 :
		TR_254 = TR_23 ;
	7'h53 :
		TR_254 = TR_23 ;
	7'h54 :
		TR_254 = TR_23 ;
	7'h55 :
		TR_254 = TR_23 ;
	7'h56 :
		TR_254 = TR_23 ;
	7'h57 :
		TR_254 = TR_23 ;
	7'h58 :
		TR_254 = TR_23 ;
	7'h59 :
		TR_254 = TR_23 ;
	7'h5a :
		TR_254 = TR_23 ;
	7'h5b :
		TR_254 = TR_23 ;
	7'h5c :
		TR_254 = TR_23 ;
	7'h5d :
		TR_254 = TR_23 ;
	7'h5e :
		TR_254 = TR_23 ;
	7'h5f :
		TR_254 = TR_23 ;
	7'h60 :
		TR_254 = TR_23 ;
	7'h61 :
		TR_254 = TR_23 ;
	7'h62 :
		TR_254 = TR_23 ;
	7'h63 :
		TR_254 = TR_23 ;
	7'h64 :
		TR_254 = TR_23 ;
	7'h65 :
		TR_254 = TR_23 ;
	7'h66 :
		TR_254 = TR_23 ;
	7'h67 :
		TR_254 = TR_23 ;
	7'h68 :
		TR_254 = TR_23 ;
	7'h69 :
		TR_254 = TR_23 ;
	7'h6a :
		TR_254 = TR_23 ;
	7'h6b :
		TR_254 = TR_23 ;
	7'h6c :
		TR_254 = TR_23 ;
	7'h6d :
		TR_254 = TR_23 ;
	7'h6e :
		TR_254 = TR_23 ;
	7'h6f :
		TR_254 = TR_23 ;
	7'h70 :
		TR_254 = TR_23 ;
	7'h71 :
		TR_254 = TR_23 ;
	7'h72 :
		TR_254 = TR_23 ;
	7'h73 :
		TR_254 = TR_23 ;
	7'h74 :
		TR_254 = TR_23 ;
	7'h75 :
		TR_254 = TR_23 ;
	7'h76 :
		TR_254 = TR_23 ;
	7'h77 :
		TR_254 = TR_23 ;
	7'h78 :
		TR_254 = TR_23 ;
	7'h79 :
		TR_254 = TR_23 ;
	7'h7a :
		TR_254 = TR_23 ;
	7'h7b :
		TR_254 = TR_23 ;
	7'h7c :
		TR_254 = TR_23 ;
	7'h7d :
		TR_254 = TR_23 ;
	7'h7e :
		TR_254 = TR_23 ;
	7'h7f :
		TR_254 = TR_23 ;
	default :
		TR_254 = 9'hx ;
	endcase
always @ ( TR_254 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_3 or 
	U_174 or RG_rl_134 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_11_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h0b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_11_t = ( ( { 9{ ST1_03d } } & RG_rl_134 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_3 )
		| ( { 9{ U_173 } } & TR_254 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_11_en = ( ST1_03d | U_174 | RG_rl_11_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_11_en )
		RG_rl_11 <= RG_rl_11_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_24 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_253 = TR_24 ;
	7'h01 :
		TR_253 = TR_24 ;
	7'h02 :
		TR_253 = TR_24 ;
	7'h03 :
		TR_253 = TR_24 ;
	7'h04 :
		TR_253 = TR_24 ;
	7'h05 :
		TR_253 = TR_24 ;
	7'h06 :
		TR_253 = TR_24 ;
	7'h07 :
		TR_253 = TR_24 ;
	7'h08 :
		TR_253 = TR_24 ;
	7'h09 :
		TR_253 = TR_24 ;
	7'h0a :
		TR_253 = TR_24 ;
	7'h0b :
		TR_253 = TR_24 ;
	7'h0c :
		TR_253 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0d :
		TR_253 = TR_24 ;
	7'h0e :
		TR_253 = TR_24 ;
	7'h0f :
		TR_253 = TR_24 ;
	7'h10 :
		TR_253 = TR_24 ;
	7'h11 :
		TR_253 = TR_24 ;
	7'h12 :
		TR_253 = TR_24 ;
	7'h13 :
		TR_253 = TR_24 ;
	7'h14 :
		TR_253 = TR_24 ;
	7'h15 :
		TR_253 = TR_24 ;
	7'h16 :
		TR_253 = TR_24 ;
	7'h17 :
		TR_253 = TR_24 ;
	7'h18 :
		TR_253 = TR_24 ;
	7'h19 :
		TR_253 = TR_24 ;
	7'h1a :
		TR_253 = TR_24 ;
	7'h1b :
		TR_253 = TR_24 ;
	7'h1c :
		TR_253 = TR_24 ;
	7'h1d :
		TR_253 = TR_24 ;
	7'h1e :
		TR_253 = TR_24 ;
	7'h1f :
		TR_253 = TR_24 ;
	7'h20 :
		TR_253 = TR_24 ;
	7'h21 :
		TR_253 = TR_24 ;
	7'h22 :
		TR_253 = TR_24 ;
	7'h23 :
		TR_253 = TR_24 ;
	7'h24 :
		TR_253 = TR_24 ;
	7'h25 :
		TR_253 = TR_24 ;
	7'h26 :
		TR_253 = TR_24 ;
	7'h27 :
		TR_253 = TR_24 ;
	7'h28 :
		TR_253 = TR_24 ;
	7'h29 :
		TR_253 = TR_24 ;
	7'h2a :
		TR_253 = TR_24 ;
	7'h2b :
		TR_253 = TR_24 ;
	7'h2c :
		TR_253 = TR_24 ;
	7'h2d :
		TR_253 = TR_24 ;
	7'h2e :
		TR_253 = TR_24 ;
	7'h2f :
		TR_253 = TR_24 ;
	7'h30 :
		TR_253 = TR_24 ;
	7'h31 :
		TR_253 = TR_24 ;
	7'h32 :
		TR_253 = TR_24 ;
	7'h33 :
		TR_253 = TR_24 ;
	7'h34 :
		TR_253 = TR_24 ;
	7'h35 :
		TR_253 = TR_24 ;
	7'h36 :
		TR_253 = TR_24 ;
	7'h37 :
		TR_253 = TR_24 ;
	7'h38 :
		TR_253 = TR_24 ;
	7'h39 :
		TR_253 = TR_24 ;
	7'h3a :
		TR_253 = TR_24 ;
	7'h3b :
		TR_253 = TR_24 ;
	7'h3c :
		TR_253 = TR_24 ;
	7'h3d :
		TR_253 = TR_24 ;
	7'h3e :
		TR_253 = TR_24 ;
	7'h3f :
		TR_253 = TR_24 ;
	7'h40 :
		TR_253 = TR_24 ;
	7'h41 :
		TR_253 = TR_24 ;
	7'h42 :
		TR_253 = TR_24 ;
	7'h43 :
		TR_253 = TR_24 ;
	7'h44 :
		TR_253 = TR_24 ;
	7'h45 :
		TR_253 = TR_24 ;
	7'h46 :
		TR_253 = TR_24 ;
	7'h47 :
		TR_253 = TR_24 ;
	7'h48 :
		TR_253 = TR_24 ;
	7'h49 :
		TR_253 = TR_24 ;
	7'h4a :
		TR_253 = TR_24 ;
	7'h4b :
		TR_253 = TR_24 ;
	7'h4c :
		TR_253 = TR_24 ;
	7'h4d :
		TR_253 = TR_24 ;
	7'h4e :
		TR_253 = TR_24 ;
	7'h4f :
		TR_253 = TR_24 ;
	7'h50 :
		TR_253 = TR_24 ;
	7'h51 :
		TR_253 = TR_24 ;
	7'h52 :
		TR_253 = TR_24 ;
	7'h53 :
		TR_253 = TR_24 ;
	7'h54 :
		TR_253 = TR_24 ;
	7'h55 :
		TR_253 = TR_24 ;
	7'h56 :
		TR_253 = TR_24 ;
	7'h57 :
		TR_253 = TR_24 ;
	7'h58 :
		TR_253 = TR_24 ;
	7'h59 :
		TR_253 = TR_24 ;
	7'h5a :
		TR_253 = TR_24 ;
	7'h5b :
		TR_253 = TR_24 ;
	7'h5c :
		TR_253 = TR_24 ;
	7'h5d :
		TR_253 = TR_24 ;
	7'h5e :
		TR_253 = TR_24 ;
	7'h5f :
		TR_253 = TR_24 ;
	7'h60 :
		TR_253 = TR_24 ;
	7'h61 :
		TR_253 = TR_24 ;
	7'h62 :
		TR_253 = TR_24 ;
	7'h63 :
		TR_253 = TR_24 ;
	7'h64 :
		TR_253 = TR_24 ;
	7'h65 :
		TR_253 = TR_24 ;
	7'h66 :
		TR_253 = TR_24 ;
	7'h67 :
		TR_253 = TR_24 ;
	7'h68 :
		TR_253 = TR_24 ;
	7'h69 :
		TR_253 = TR_24 ;
	7'h6a :
		TR_253 = TR_24 ;
	7'h6b :
		TR_253 = TR_24 ;
	7'h6c :
		TR_253 = TR_24 ;
	7'h6d :
		TR_253 = TR_24 ;
	7'h6e :
		TR_253 = TR_24 ;
	7'h6f :
		TR_253 = TR_24 ;
	7'h70 :
		TR_253 = TR_24 ;
	7'h71 :
		TR_253 = TR_24 ;
	7'h72 :
		TR_253 = TR_24 ;
	7'h73 :
		TR_253 = TR_24 ;
	7'h74 :
		TR_253 = TR_24 ;
	7'h75 :
		TR_253 = TR_24 ;
	7'h76 :
		TR_253 = TR_24 ;
	7'h77 :
		TR_253 = TR_24 ;
	7'h78 :
		TR_253 = TR_24 ;
	7'h79 :
		TR_253 = TR_24 ;
	7'h7a :
		TR_253 = TR_24 ;
	7'h7b :
		TR_253 = TR_24 ;
	7'h7c :
		TR_253 = TR_24 ;
	7'h7d :
		TR_253 = TR_24 ;
	7'h7e :
		TR_253 = TR_24 ;
	7'h7f :
		TR_253 = TR_24 ;
	default :
		TR_253 = 9'hx ;
	endcase
always @ ( TR_253 or U_173 or sub8u_71ot or U_183 or RG_rl_135 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_12_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h0c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_12_t = ( ( { 9{ M_180 } } & RG_rl_135 )
		| ( { 9{ U_173 } } & TR_253 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_12_en = ( M_180 | RG_rl_12_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_12_en )
		RG_rl_12 <= RG_rl_12_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_25 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_252 = TR_25 ;
	7'h01 :
		TR_252 = TR_25 ;
	7'h02 :
		TR_252 = TR_25 ;
	7'h03 :
		TR_252 = TR_25 ;
	7'h04 :
		TR_252 = TR_25 ;
	7'h05 :
		TR_252 = TR_25 ;
	7'h06 :
		TR_252 = TR_25 ;
	7'h07 :
		TR_252 = TR_25 ;
	7'h08 :
		TR_252 = TR_25 ;
	7'h09 :
		TR_252 = TR_25 ;
	7'h0a :
		TR_252 = TR_25 ;
	7'h0b :
		TR_252 = TR_25 ;
	7'h0c :
		TR_252 = TR_25 ;
	7'h0d :
		TR_252 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0e :
		TR_252 = TR_25 ;
	7'h0f :
		TR_252 = TR_25 ;
	7'h10 :
		TR_252 = TR_25 ;
	7'h11 :
		TR_252 = TR_25 ;
	7'h12 :
		TR_252 = TR_25 ;
	7'h13 :
		TR_252 = TR_25 ;
	7'h14 :
		TR_252 = TR_25 ;
	7'h15 :
		TR_252 = TR_25 ;
	7'h16 :
		TR_252 = TR_25 ;
	7'h17 :
		TR_252 = TR_25 ;
	7'h18 :
		TR_252 = TR_25 ;
	7'h19 :
		TR_252 = TR_25 ;
	7'h1a :
		TR_252 = TR_25 ;
	7'h1b :
		TR_252 = TR_25 ;
	7'h1c :
		TR_252 = TR_25 ;
	7'h1d :
		TR_252 = TR_25 ;
	7'h1e :
		TR_252 = TR_25 ;
	7'h1f :
		TR_252 = TR_25 ;
	7'h20 :
		TR_252 = TR_25 ;
	7'h21 :
		TR_252 = TR_25 ;
	7'h22 :
		TR_252 = TR_25 ;
	7'h23 :
		TR_252 = TR_25 ;
	7'h24 :
		TR_252 = TR_25 ;
	7'h25 :
		TR_252 = TR_25 ;
	7'h26 :
		TR_252 = TR_25 ;
	7'h27 :
		TR_252 = TR_25 ;
	7'h28 :
		TR_252 = TR_25 ;
	7'h29 :
		TR_252 = TR_25 ;
	7'h2a :
		TR_252 = TR_25 ;
	7'h2b :
		TR_252 = TR_25 ;
	7'h2c :
		TR_252 = TR_25 ;
	7'h2d :
		TR_252 = TR_25 ;
	7'h2e :
		TR_252 = TR_25 ;
	7'h2f :
		TR_252 = TR_25 ;
	7'h30 :
		TR_252 = TR_25 ;
	7'h31 :
		TR_252 = TR_25 ;
	7'h32 :
		TR_252 = TR_25 ;
	7'h33 :
		TR_252 = TR_25 ;
	7'h34 :
		TR_252 = TR_25 ;
	7'h35 :
		TR_252 = TR_25 ;
	7'h36 :
		TR_252 = TR_25 ;
	7'h37 :
		TR_252 = TR_25 ;
	7'h38 :
		TR_252 = TR_25 ;
	7'h39 :
		TR_252 = TR_25 ;
	7'h3a :
		TR_252 = TR_25 ;
	7'h3b :
		TR_252 = TR_25 ;
	7'h3c :
		TR_252 = TR_25 ;
	7'h3d :
		TR_252 = TR_25 ;
	7'h3e :
		TR_252 = TR_25 ;
	7'h3f :
		TR_252 = TR_25 ;
	7'h40 :
		TR_252 = TR_25 ;
	7'h41 :
		TR_252 = TR_25 ;
	7'h42 :
		TR_252 = TR_25 ;
	7'h43 :
		TR_252 = TR_25 ;
	7'h44 :
		TR_252 = TR_25 ;
	7'h45 :
		TR_252 = TR_25 ;
	7'h46 :
		TR_252 = TR_25 ;
	7'h47 :
		TR_252 = TR_25 ;
	7'h48 :
		TR_252 = TR_25 ;
	7'h49 :
		TR_252 = TR_25 ;
	7'h4a :
		TR_252 = TR_25 ;
	7'h4b :
		TR_252 = TR_25 ;
	7'h4c :
		TR_252 = TR_25 ;
	7'h4d :
		TR_252 = TR_25 ;
	7'h4e :
		TR_252 = TR_25 ;
	7'h4f :
		TR_252 = TR_25 ;
	7'h50 :
		TR_252 = TR_25 ;
	7'h51 :
		TR_252 = TR_25 ;
	7'h52 :
		TR_252 = TR_25 ;
	7'h53 :
		TR_252 = TR_25 ;
	7'h54 :
		TR_252 = TR_25 ;
	7'h55 :
		TR_252 = TR_25 ;
	7'h56 :
		TR_252 = TR_25 ;
	7'h57 :
		TR_252 = TR_25 ;
	7'h58 :
		TR_252 = TR_25 ;
	7'h59 :
		TR_252 = TR_25 ;
	7'h5a :
		TR_252 = TR_25 ;
	7'h5b :
		TR_252 = TR_25 ;
	7'h5c :
		TR_252 = TR_25 ;
	7'h5d :
		TR_252 = TR_25 ;
	7'h5e :
		TR_252 = TR_25 ;
	7'h5f :
		TR_252 = TR_25 ;
	7'h60 :
		TR_252 = TR_25 ;
	7'h61 :
		TR_252 = TR_25 ;
	7'h62 :
		TR_252 = TR_25 ;
	7'h63 :
		TR_252 = TR_25 ;
	7'h64 :
		TR_252 = TR_25 ;
	7'h65 :
		TR_252 = TR_25 ;
	7'h66 :
		TR_252 = TR_25 ;
	7'h67 :
		TR_252 = TR_25 ;
	7'h68 :
		TR_252 = TR_25 ;
	7'h69 :
		TR_252 = TR_25 ;
	7'h6a :
		TR_252 = TR_25 ;
	7'h6b :
		TR_252 = TR_25 ;
	7'h6c :
		TR_252 = TR_25 ;
	7'h6d :
		TR_252 = TR_25 ;
	7'h6e :
		TR_252 = TR_25 ;
	7'h6f :
		TR_252 = TR_25 ;
	7'h70 :
		TR_252 = TR_25 ;
	7'h71 :
		TR_252 = TR_25 ;
	7'h72 :
		TR_252 = TR_25 ;
	7'h73 :
		TR_252 = TR_25 ;
	7'h74 :
		TR_252 = TR_25 ;
	7'h75 :
		TR_252 = TR_25 ;
	7'h76 :
		TR_252 = TR_25 ;
	7'h77 :
		TR_252 = TR_25 ;
	7'h78 :
		TR_252 = TR_25 ;
	7'h79 :
		TR_252 = TR_25 ;
	7'h7a :
		TR_252 = TR_25 ;
	7'h7b :
		TR_252 = TR_25 ;
	7'h7c :
		TR_252 = TR_25 ;
	7'h7d :
		TR_252 = TR_25 ;
	7'h7e :
		TR_252 = TR_25 ;
	7'h7f :
		TR_252 = TR_25 ;
	default :
		TR_252 = 9'hx ;
	endcase
always @ ( TR_252 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_4 or 
	U_174 or RG_rl_135 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_13_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h0d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_13_t = ( ( { 9{ ST1_03d } } & RG_rl_135 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_4 )
		| ( { 9{ U_173 } } & TR_252 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_13_en = ( ST1_03d | U_174 | RG_rl_13_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_13_en )
		RG_rl_13 <= RG_rl_13_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_26 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_251 = TR_26 ;
	7'h01 :
		TR_251 = TR_26 ;
	7'h02 :
		TR_251 = TR_26 ;
	7'h03 :
		TR_251 = TR_26 ;
	7'h04 :
		TR_251 = TR_26 ;
	7'h05 :
		TR_251 = TR_26 ;
	7'h06 :
		TR_251 = TR_26 ;
	7'h07 :
		TR_251 = TR_26 ;
	7'h08 :
		TR_251 = TR_26 ;
	7'h09 :
		TR_251 = TR_26 ;
	7'h0a :
		TR_251 = TR_26 ;
	7'h0b :
		TR_251 = TR_26 ;
	7'h0c :
		TR_251 = TR_26 ;
	7'h0d :
		TR_251 = TR_26 ;
	7'h0e :
		TR_251 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0f :
		TR_251 = TR_26 ;
	7'h10 :
		TR_251 = TR_26 ;
	7'h11 :
		TR_251 = TR_26 ;
	7'h12 :
		TR_251 = TR_26 ;
	7'h13 :
		TR_251 = TR_26 ;
	7'h14 :
		TR_251 = TR_26 ;
	7'h15 :
		TR_251 = TR_26 ;
	7'h16 :
		TR_251 = TR_26 ;
	7'h17 :
		TR_251 = TR_26 ;
	7'h18 :
		TR_251 = TR_26 ;
	7'h19 :
		TR_251 = TR_26 ;
	7'h1a :
		TR_251 = TR_26 ;
	7'h1b :
		TR_251 = TR_26 ;
	7'h1c :
		TR_251 = TR_26 ;
	7'h1d :
		TR_251 = TR_26 ;
	7'h1e :
		TR_251 = TR_26 ;
	7'h1f :
		TR_251 = TR_26 ;
	7'h20 :
		TR_251 = TR_26 ;
	7'h21 :
		TR_251 = TR_26 ;
	7'h22 :
		TR_251 = TR_26 ;
	7'h23 :
		TR_251 = TR_26 ;
	7'h24 :
		TR_251 = TR_26 ;
	7'h25 :
		TR_251 = TR_26 ;
	7'h26 :
		TR_251 = TR_26 ;
	7'h27 :
		TR_251 = TR_26 ;
	7'h28 :
		TR_251 = TR_26 ;
	7'h29 :
		TR_251 = TR_26 ;
	7'h2a :
		TR_251 = TR_26 ;
	7'h2b :
		TR_251 = TR_26 ;
	7'h2c :
		TR_251 = TR_26 ;
	7'h2d :
		TR_251 = TR_26 ;
	7'h2e :
		TR_251 = TR_26 ;
	7'h2f :
		TR_251 = TR_26 ;
	7'h30 :
		TR_251 = TR_26 ;
	7'h31 :
		TR_251 = TR_26 ;
	7'h32 :
		TR_251 = TR_26 ;
	7'h33 :
		TR_251 = TR_26 ;
	7'h34 :
		TR_251 = TR_26 ;
	7'h35 :
		TR_251 = TR_26 ;
	7'h36 :
		TR_251 = TR_26 ;
	7'h37 :
		TR_251 = TR_26 ;
	7'h38 :
		TR_251 = TR_26 ;
	7'h39 :
		TR_251 = TR_26 ;
	7'h3a :
		TR_251 = TR_26 ;
	7'h3b :
		TR_251 = TR_26 ;
	7'h3c :
		TR_251 = TR_26 ;
	7'h3d :
		TR_251 = TR_26 ;
	7'h3e :
		TR_251 = TR_26 ;
	7'h3f :
		TR_251 = TR_26 ;
	7'h40 :
		TR_251 = TR_26 ;
	7'h41 :
		TR_251 = TR_26 ;
	7'h42 :
		TR_251 = TR_26 ;
	7'h43 :
		TR_251 = TR_26 ;
	7'h44 :
		TR_251 = TR_26 ;
	7'h45 :
		TR_251 = TR_26 ;
	7'h46 :
		TR_251 = TR_26 ;
	7'h47 :
		TR_251 = TR_26 ;
	7'h48 :
		TR_251 = TR_26 ;
	7'h49 :
		TR_251 = TR_26 ;
	7'h4a :
		TR_251 = TR_26 ;
	7'h4b :
		TR_251 = TR_26 ;
	7'h4c :
		TR_251 = TR_26 ;
	7'h4d :
		TR_251 = TR_26 ;
	7'h4e :
		TR_251 = TR_26 ;
	7'h4f :
		TR_251 = TR_26 ;
	7'h50 :
		TR_251 = TR_26 ;
	7'h51 :
		TR_251 = TR_26 ;
	7'h52 :
		TR_251 = TR_26 ;
	7'h53 :
		TR_251 = TR_26 ;
	7'h54 :
		TR_251 = TR_26 ;
	7'h55 :
		TR_251 = TR_26 ;
	7'h56 :
		TR_251 = TR_26 ;
	7'h57 :
		TR_251 = TR_26 ;
	7'h58 :
		TR_251 = TR_26 ;
	7'h59 :
		TR_251 = TR_26 ;
	7'h5a :
		TR_251 = TR_26 ;
	7'h5b :
		TR_251 = TR_26 ;
	7'h5c :
		TR_251 = TR_26 ;
	7'h5d :
		TR_251 = TR_26 ;
	7'h5e :
		TR_251 = TR_26 ;
	7'h5f :
		TR_251 = TR_26 ;
	7'h60 :
		TR_251 = TR_26 ;
	7'h61 :
		TR_251 = TR_26 ;
	7'h62 :
		TR_251 = TR_26 ;
	7'h63 :
		TR_251 = TR_26 ;
	7'h64 :
		TR_251 = TR_26 ;
	7'h65 :
		TR_251 = TR_26 ;
	7'h66 :
		TR_251 = TR_26 ;
	7'h67 :
		TR_251 = TR_26 ;
	7'h68 :
		TR_251 = TR_26 ;
	7'h69 :
		TR_251 = TR_26 ;
	7'h6a :
		TR_251 = TR_26 ;
	7'h6b :
		TR_251 = TR_26 ;
	7'h6c :
		TR_251 = TR_26 ;
	7'h6d :
		TR_251 = TR_26 ;
	7'h6e :
		TR_251 = TR_26 ;
	7'h6f :
		TR_251 = TR_26 ;
	7'h70 :
		TR_251 = TR_26 ;
	7'h71 :
		TR_251 = TR_26 ;
	7'h72 :
		TR_251 = TR_26 ;
	7'h73 :
		TR_251 = TR_26 ;
	7'h74 :
		TR_251 = TR_26 ;
	7'h75 :
		TR_251 = TR_26 ;
	7'h76 :
		TR_251 = TR_26 ;
	7'h77 :
		TR_251 = TR_26 ;
	7'h78 :
		TR_251 = TR_26 ;
	7'h79 :
		TR_251 = TR_26 ;
	7'h7a :
		TR_251 = TR_26 ;
	7'h7b :
		TR_251 = TR_26 ;
	7'h7c :
		TR_251 = TR_26 ;
	7'h7d :
		TR_251 = TR_26 ;
	7'h7e :
		TR_251 = TR_26 ;
	7'h7f :
		TR_251 = TR_26 ;
	default :
		TR_251 = 9'hx ;
	endcase
always @ ( TR_251 or U_173 or sub8u_71ot or U_183 or RG_rl_136 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_14_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h0e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_14_t = ( ( { 9{ M_180 } } & RG_rl_136 )
		| ( { 9{ U_173 } } & TR_251 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_14_en = ( M_180 | RG_rl_14_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_14_en )
		RG_rl_14 <= RG_rl_14_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_27 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_250 = TR_27 ;
	7'h01 :
		TR_250 = TR_27 ;
	7'h02 :
		TR_250 = TR_27 ;
	7'h03 :
		TR_250 = TR_27 ;
	7'h04 :
		TR_250 = TR_27 ;
	7'h05 :
		TR_250 = TR_27 ;
	7'h06 :
		TR_250 = TR_27 ;
	7'h07 :
		TR_250 = TR_27 ;
	7'h08 :
		TR_250 = TR_27 ;
	7'h09 :
		TR_250 = TR_27 ;
	7'h0a :
		TR_250 = TR_27 ;
	7'h0b :
		TR_250 = TR_27 ;
	7'h0c :
		TR_250 = TR_27 ;
	7'h0d :
		TR_250 = TR_27 ;
	7'h0e :
		TR_250 = TR_27 ;
	7'h0f :
		TR_250 = 9'h000 ;	// line#=../rle.cpp:80
	7'h10 :
		TR_250 = TR_27 ;
	7'h11 :
		TR_250 = TR_27 ;
	7'h12 :
		TR_250 = TR_27 ;
	7'h13 :
		TR_250 = TR_27 ;
	7'h14 :
		TR_250 = TR_27 ;
	7'h15 :
		TR_250 = TR_27 ;
	7'h16 :
		TR_250 = TR_27 ;
	7'h17 :
		TR_250 = TR_27 ;
	7'h18 :
		TR_250 = TR_27 ;
	7'h19 :
		TR_250 = TR_27 ;
	7'h1a :
		TR_250 = TR_27 ;
	7'h1b :
		TR_250 = TR_27 ;
	7'h1c :
		TR_250 = TR_27 ;
	7'h1d :
		TR_250 = TR_27 ;
	7'h1e :
		TR_250 = TR_27 ;
	7'h1f :
		TR_250 = TR_27 ;
	7'h20 :
		TR_250 = TR_27 ;
	7'h21 :
		TR_250 = TR_27 ;
	7'h22 :
		TR_250 = TR_27 ;
	7'h23 :
		TR_250 = TR_27 ;
	7'h24 :
		TR_250 = TR_27 ;
	7'h25 :
		TR_250 = TR_27 ;
	7'h26 :
		TR_250 = TR_27 ;
	7'h27 :
		TR_250 = TR_27 ;
	7'h28 :
		TR_250 = TR_27 ;
	7'h29 :
		TR_250 = TR_27 ;
	7'h2a :
		TR_250 = TR_27 ;
	7'h2b :
		TR_250 = TR_27 ;
	7'h2c :
		TR_250 = TR_27 ;
	7'h2d :
		TR_250 = TR_27 ;
	7'h2e :
		TR_250 = TR_27 ;
	7'h2f :
		TR_250 = TR_27 ;
	7'h30 :
		TR_250 = TR_27 ;
	7'h31 :
		TR_250 = TR_27 ;
	7'h32 :
		TR_250 = TR_27 ;
	7'h33 :
		TR_250 = TR_27 ;
	7'h34 :
		TR_250 = TR_27 ;
	7'h35 :
		TR_250 = TR_27 ;
	7'h36 :
		TR_250 = TR_27 ;
	7'h37 :
		TR_250 = TR_27 ;
	7'h38 :
		TR_250 = TR_27 ;
	7'h39 :
		TR_250 = TR_27 ;
	7'h3a :
		TR_250 = TR_27 ;
	7'h3b :
		TR_250 = TR_27 ;
	7'h3c :
		TR_250 = TR_27 ;
	7'h3d :
		TR_250 = TR_27 ;
	7'h3e :
		TR_250 = TR_27 ;
	7'h3f :
		TR_250 = TR_27 ;
	7'h40 :
		TR_250 = TR_27 ;
	7'h41 :
		TR_250 = TR_27 ;
	7'h42 :
		TR_250 = TR_27 ;
	7'h43 :
		TR_250 = TR_27 ;
	7'h44 :
		TR_250 = TR_27 ;
	7'h45 :
		TR_250 = TR_27 ;
	7'h46 :
		TR_250 = TR_27 ;
	7'h47 :
		TR_250 = TR_27 ;
	7'h48 :
		TR_250 = TR_27 ;
	7'h49 :
		TR_250 = TR_27 ;
	7'h4a :
		TR_250 = TR_27 ;
	7'h4b :
		TR_250 = TR_27 ;
	7'h4c :
		TR_250 = TR_27 ;
	7'h4d :
		TR_250 = TR_27 ;
	7'h4e :
		TR_250 = TR_27 ;
	7'h4f :
		TR_250 = TR_27 ;
	7'h50 :
		TR_250 = TR_27 ;
	7'h51 :
		TR_250 = TR_27 ;
	7'h52 :
		TR_250 = TR_27 ;
	7'h53 :
		TR_250 = TR_27 ;
	7'h54 :
		TR_250 = TR_27 ;
	7'h55 :
		TR_250 = TR_27 ;
	7'h56 :
		TR_250 = TR_27 ;
	7'h57 :
		TR_250 = TR_27 ;
	7'h58 :
		TR_250 = TR_27 ;
	7'h59 :
		TR_250 = TR_27 ;
	7'h5a :
		TR_250 = TR_27 ;
	7'h5b :
		TR_250 = TR_27 ;
	7'h5c :
		TR_250 = TR_27 ;
	7'h5d :
		TR_250 = TR_27 ;
	7'h5e :
		TR_250 = TR_27 ;
	7'h5f :
		TR_250 = TR_27 ;
	7'h60 :
		TR_250 = TR_27 ;
	7'h61 :
		TR_250 = TR_27 ;
	7'h62 :
		TR_250 = TR_27 ;
	7'h63 :
		TR_250 = TR_27 ;
	7'h64 :
		TR_250 = TR_27 ;
	7'h65 :
		TR_250 = TR_27 ;
	7'h66 :
		TR_250 = TR_27 ;
	7'h67 :
		TR_250 = TR_27 ;
	7'h68 :
		TR_250 = TR_27 ;
	7'h69 :
		TR_250 = TR_27 ;
	7'h6a :
		TR_250 = TR_27 ;
	7'h6b :
		TR_250 = TR_27 ;
	7'h6c :
		TR_250 = TR_27 ;
	7'h6d :
		TR_250 = TR_27 ;
	7'h6e :
		TR_250 = TR_27 ;
	7'h6f :
		TR_250 = TR_27 ;
	7'h70 :
		TR_250 = TR_27 ;
	7'h71 :
		TR_250 = TR_27 ;
	7'h72 :
		TR_250 = TR_27 ;
	7'h73 :
		TR_250 = TR_27 ;
	7'h74 :
		TR_250 = TR_27 ;
	7'h75 :
		TR_250 = TR_27 ;
	7'h76 :
		TR_250 = TR_27 ;
	7'h77 :
		TR_250 = TR_27 ;
	7'h78 :
		TR_250 = TR_27 ;
	7'h79 :
		TR_250 = TR_27 ;
	7'h7a :
		TR_250 = TR_27 ;
	7'h7b :
		TR_250 = TR_27 ;
	7'h7c :
		TR_250 = TR_27 ;
	7'h7d :
		TR_250 = TR_27 ;
	7'h7e :
		TR_250 = TR_27 ;
	7'h7f :
		TR_250 = TR_27 ;
	default :
		TR_250 = 9'hx ;
	endcase
always @ ( TR_250 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_5 or 
	U_174 or RG_rl_136 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_15_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h0f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_15_t = ( ( { 9{ ST1_03d } } & RG_rl_136 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_5 )
		| ( { 9{ U_173 } } & TR_250 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_15_en = ( ST1_03d | U_174 | RG_rl_15_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_15_en )
		RG_rl_15 <= RG_rl_15_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_28 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_249 = TR_28 ;
	7'h01 :
		TR_249 = TR_28 ;
	7'h02 :
		TR_249 = TR_28 ;
	7'h03 :
		TR_249 = TR_28 ;
	7'h04 :
		TR_249 = TR_28 ;
	7'h05 :
		TR_249 = TR_28 ;
	7'h06 :
		TR_249 = TR_28 ;
	7'h07 :
		TR_249 = TR_28 ;
	7'h08 :
		TR_249 = TR_28 ;
	7'h09 :
		TR_249 = TR_28 ;
	7'h0a :
		TR_249 = TR_28 ;
	7'h0b :
		TR_249 = TR_28 ;
	7'h0c :
		TR_249 = TR_28 ;
	7'h0d :
		TR_249 = TR_28 ;
	7'h0e :
		TR_249 = TR_28 ;
	7'h0f :
		TR_249 = TR_28 ;
	7'h10 :
		TR_249 = 9'h000 ;	// line#=../rle.cpp:80
	7'h11 :
		TR_249 = TR_28 ;
	7'h12 :
		TR_249 = TR_28 ;
	7'h13 :
		TR_249 = TR_28 ;
	7'h14 :
		TR_249 = TR_28 ;
	7'h15 :
		TR_249 = TR_28 ;
	7'h16 :
		TR_249 = TR_28 ;
	7'h17 :
		TR_249 = TR_28 ;
	7'h18 :
		TR_249 = TR_28 ;
	7'h19 :
		TR_249 = TR_28 ;
	7'h1a :
		TR_249 = TR_28 ;
	7'h1b :
		TR_249 = TR_28 ;
	7'h1c :
		TR_249 = TR_28 ;
	7'h1d :
		TR_249 = TR_28 ;
	7'h1e :
		TR_249 = TR_28 ;
	7'h1f :
		TR_249 = TR_28 ;
	7'h20 :
		TR_249 = TR_28 ;
	7'h21 :
		TR_249 = TR_28 ;
	7'h22 :
		TR_249 = TR_28 ;
	7'h23 :
		TR_249 = TR_28 ;
	7'h24 :
		TR_249 = TR_28 ;
	7'h25 :
		TR_249 = TR_28 ;
	7'h26 :
		TR_249 = TR_28 ;
	7'h27 :
		TR_249 = TR_28 ;
	7'h28 :
		TR_249 = TR_28 ;
	7'h29 :
		TR_249 = TR_28 ;
	7'h2a :
		TR_249 = TR_28 ;
	7'h2b :
		TR_249 = TR_28 ;
	7'h2c :
		TR_249 = TR_28 ;
	7'h2d :
		TR_249 = TR_28 ;
	7'h2e :
		TR_249 = TR_28 ;
	7'h2f :
		TR_249 = TR_28 ;
	7'h30 :
		TR_249 = TR_28 ;
	7'h31 :
		TR_249 = TR_28 ;
	7'h32 :
		TR_249 = TR_28 ;
	7'h33 :
		TR_249 = TR_28 ;
	7'h34 :
		TR_249 = TR_28 ;
	7'h35 :
		TR_249 = TR_28 ;
	7'h36 :
		TR_249 = TR_28 ;
	7'h37 :
		TR_249 = TR_28 ;
	7'h38 :
		TR_249 = TR_28 ;
	7'h39 :
		TR_249 = TR_28 ;
	7'h3a :
		TR_249 = TR_28 ;
	7'h3b :
		TR_249 = TR_28 ;
	7'h3c :
		TR_249 = TR_28 ;
	7'h3d :
		TR_249 = TR_28 ;
	7'h3e :
		TR_249 = TR_28 ;
	7'h3f :
		TR_249 = TR_28 ;
	7'h40 :
		TR_249 = TR_28 ;
	7'h41 :
		TR_249 = TR_28 ;
	7'h42 :
		TR_249 = TR_28 ;
	7'h43 :
		TR_249 = TR_28 ;
	7'h44 :
		TR_249 = TR_28 ;
	7'h45 :
		TR_249 = TR_28 ;
	7'h46 :
		TR_249 = TR_28 ;
	7'h47 :
		TR_249 = TR_28 ;
	7'h48 :
		TR_249 = TR_28 ;
	7'h49 :
		TR_249 = TR_28 ;
	7'h4a :
		TR_249 = TR_28 ;
	7'h4b :
		TR_249 = TR_28 ;
	7'h4c :
		TR_249 = TR_28 ;
	7'h4d :
		TR_249 = TR_28 ;
	7'h4e :
		TR_249 = TR_28 ;
	7'h4f :
		TR_249 = TR_28 ;
	7'h50 :
		TR_249 = TR_28 ;
	7'h51 :
		TR_249 = TR_28 ;
	7'h52 :
		TR_249 = TR_28 ;
	7'h53 :
		TR_249 = TR_28 ;
	7'h54 :
		TR_249 = TR_28 ;
	7'h55 :
		TR_249 = TR_28 ;
	7'h56 :
		TR_249 = TR_28 ;
	7'h57 :
		TR_249 = TR_28 ;
	7'h58 :
		TR_249 = TR_28 ;
	7'h59 :
		TR_249 = TR_28 ;
	7'h5a :
		TR_249 = TR_28 ;
	7'h5b :
		TR_249 = TR_28 ;
	7'h5c :
		TR_249 = TR_28 ;
	7'h5d :
		TR_249 = TR_28 ;
	7'h5e :
		TR_249 = TR_28 ;
	7'h5f :
		TR_249 = TR_28 ;
	7'h60 :
		TR_249 = TR_28 ;
	7'h61 :
		TR_249 = TR_28 ;
	7'h62 :
		TR_249 = TR_28 ;
	7'h63 :
		TR_249 = TR_28 ;
	7'h64 :
		TR_249 = TR_28 ;
	7'h65 :
		TR_249 = TR_28 ;
	7'h66 :
		TR_249 = TR_28 ;
	7'h67 :
		TR_249 = TR_28 ;
	7'h68 :
		TR_249 = TR_28 ;
	7'h69 :
		TR_249 = TR_28 ;
	7'h6a :
		TR_249 = TR_28 ;
	7'h6b :
		TR_249 = TR_28 ;
	7'h6c :
		TR_249 = TR_28 ;
	7'h6d :
		TR_249 = TR_28 ;
	7'h6e :
		TR_249 = TR_28 ;
	7'h6f :
		TR_249 = TR_28 ;
	7'h70 :
		TR_249 = TR_28 ;
	7'h71 :
		TR_249 = TR_28 ;
	7'h72 :
		TR_249 = TR_28 ;
	7'h73 :
		TR_249 = TR_28 ;
	7'h74 :
		TR_249 = TR_28 ;
	7'h75 :
		TR_249 = TR_28 ;
	7'h76 :
		TR_249 = TR_28 ;
	7'h77 :
		TR_249 = TR_28 ;
	7'h78 :
		TR_249 = TR_28 ;
	7'h79 :
		TR_249 = TR_28 ;
	7'h7a :
		TR_249 = TR_28 ;
	7'h7b :
		TR_249 = TR_28 ;
	7'h7c :
		TR_249 = TR_28 ;
	7'h7d :
		TR_249 = TR_28 ;
	7'h7e :
		TR_249 = TR_28 ;
	7'h7f :
		TR_249 = TR_28 ;
	default :
		TR_249 = 9'hx ;
	endcase
always @ ( TR_249 or U_173 or sub8u_71ot or U_183 or RG_rl_137 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_16_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h10 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_16_t = ( ( { 9{ M_180 } } & RG_rl_137 )
		| ( { 9{ U_173 } } & TR_249 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_16_en = ( M_180 | RG_rl_16_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_16_en )
		RG_rl_16 <= RG_rl_16_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_29 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_248 = TR_29 ;
	7'h01 :
		TR_248 = TR_29 ;
	7'h02 :
		TR_248 = TR_29 ;
	7'h03 :
		TR_248 = TR_29 ;
	7'h04 :
		TR_248 = TR_29 ;
	7'h05 :
		TR_248 = TR_29 ;
	7'h06 :
		TR_248 = TR_29 ;
	7'h07 :
		TR_248 = TR_29 ;
	7'h08 :
		TR_248 = TR_29 ;
	7'h09 :
		TR_248 = TR_29 ;
	7'h0a :
		TR_248 = TR_29 ;
	7'h0b :
		TR_248 = TR_29 ;
	7'h0c :
		TR_248 = TR_29 ;
	7'h0d :
		TR_248 = TR_29 ;
	7'h0e :
		TR_248 = TR_29 ;
	7'h0f :
		TR_248 = TR_29 ;
	7'h10 :
		TR_248 = TR_29 ;
	7'h11 :
		TR_248 = 9'h000 ;	// line#=../rle.cpp:80
	7'h12 :
		TR_248 = TR_29 ;
	7'h13 :
		TR_248 = TR_29 ;
	7'h14 :
		TR_248 = TR_29 ;
	7'h15 :
		TR_248 = TR_29 ;
	7'h16 :
		TR_248 = TR_29 ;
	7'h17 :
		TR_248 = TR_29 ;
	7'h18 :
		TR_248 = TR_29 ;
	7'h19 :
		TR_248 = TR_29 ;
	7'h1a :
		TR_248 = TR_29 ;
	7'h1b :
		TR_248 = TR_29 ;
	7'h1c :
		TR_248 = TR_29 ;
	7'h1d :
		TR_248 = TR_29 ;
	7'h1e :
		TR_248 = TR_29 ;
	7'h1f :
		TR_248 = TR_29 ;
	7'h20 :
		TR_248 = TR_29 ;
	7'h21 :
		TR_248 = TR_29 ;
	7'h22 :
		TR_248 = TR_29 ;
	7'h23 :
		TR_248 = TR_29 ;
	7'h24 :
		TR_248 = TR_29 ;
	7'h25 :
		TR_248 = TR_29 ;
	7'h26 :
		TR_248 = TR_29 ;
	7'h27 :
		TR_248 = TR_29 ;
	7'h28 :
		TR_248 = TR_29 ;
	7'h29 :
		TR_248 = TR_29 ;
	7'h2a :
		TR_248 = TR_29 ;
	7'h2b :
		TR_248 = TR_29 ;
	7'h2c :
		TR_248 = TR_29 ;
	7'h2d :
		TR_248 = TR_29 ;
	7'h2e :
		TR_248 = TR_29 ;
	7'h2f :
		TR_248 = TR_29 ;
	7'h30 :
		TR_248 = TR_29 ;
	7'h31 :
		TR_248 = TR_29 ;
	7'h32 :
		TR_248 = TR_29 ;
	7'h33 :
		TR_248 = TR_29 ;
	7'h34 :
		TR_248 = TR_29 ;
	7'h35 :
		TR_248 = TR_29 ;
	7'h36 :
		TR_248 = TR_29 ;
	7'h37 :
		TR_248 = TR_29 ;
	7'h38 :
		TR_248 = TR_29 ;
	7'h39 :
		TR_248 = TR_29 ;
	7'h3a :
		TR_248 = TR_29 ;
	7'h3b :
		TR_248 = TR_29 ;
	7'h3c :
		TR_248 = TR_29 ;
	7'h3d :
		TR_248 = TR_29 ;
	7'h3e :
		TR_248 = TR_29 ;
	7'h3f :
		TR_248 = TR_29 ;
	7'h40 :
		TR_248 = TR_29 ;
	7'h41 :
		TR_248 = TR_29 ;
	7'h42 :
		TR_248 = TR_29 ;
	7'h43 :
		TR_248 = TR_29 ;
	7'h44 :
		TR_248 = TR_29 ;
	7'h45 :
		TR_248 = TR_29 ;
	7'h46 :
		TR_248 = TR_29 ;
	7'h47 :
		TR_248 = TR_29 ;
	7'h48 :
		TR_248 = TR_29 ;
	7'h49 :
		TR_248 = TR_29 ;
	7'h4a :
		TR_248 = TR_29 ;
	7'h4b :
		TR_248 = TR_29 ;
	7'h4c :
		TR_248 = TR_29 ;
	7'h4d :
		TR_248 = TR_29 ;
	7'h4e :
		TR_248 = TR_29 ;
	7'h4f :
		TR_248 = TR_29 ;
	7'h50 :
		TR_248 = TR_29 ;
	7'h51 :
		TR_248 = TR_29 ;
	7'h52 :
		TR_248 = TR_29 ;
	7'h53 :
		TR_248 = TR_29 ;
	7'h54 :
		TR_248 = TR_29 ;
	7'h55 :
		TR_248 = TR_29 ;
	7'h56 :
		TR_248 = TR_29 ;
	7'h57 :
		TR_248 = TR_29 ;
	7'h58 :
		TR_248 = TR_29 ;
	7'h59 :
		TR_248 = TR_29 ;
	7'h5a :
		TR_248 = TR_29 ;
	7'h5b :
		TR_248 = TR_29 ;
	7'h5c :
		TR_248 = TR_29 ;
	7'h5d :
		TR_248 = TR_29 ;
	7'h5e :
		TR_248 = TR_29 ;
	7'h5f :
		TR_248 = TR_29 ;
	7'h60 :
		TR_248 = TR_29 ;
	7'h61 :
		TR_248 = TR_29 ;
	7'h62 :
		TR_248 = TR_29 ;
	7'h63 :
		TR_248 = TR_29 ;
	7'h64 :
		TR_248 = TR_29 ;
	7'h65 :
		TR_248 = TR_29 ;
	7'h66 :
		TR_248 = TR_29 ;
	7'h67 :
		TR_248 = TR_29 ;
	7'h68 :
		TR_248 = TR_29 ;
	7'h69 :
		TR_248 = TR_29 ;
	7'h6a :
		TR_248 = TR_29 ;
	7'h6b :
		TR_248 = TR_29 ;
	7'h6c :
		TR_248 = TR_29 ;
	7'h6d :
		TR_248 = TR_29 ;
	7'h6e :
		TR_248 = TR_29 ;
	7'h6f :
		TR_248 = TR_29 ;
	7'h70 :
		TR_248 = TR_29 ;
	7'h71 :
		TR_248 = TR_29 ;
	7'h72 :
		TR_248 = TR_29 ;
	7'h73 :
		TR_248 = TR_29 ;
	7'h74 :
		TR_248 = TR_29 ;
	7'h75 :
		TR_248 = TR_29 ;
	7'h76 :
		TR_248 = TR_29 ;
	7'h77 :
		TR_248 = TR_29 ;
	7'h78 :
		TR_248 = TR_29 ;
	7'h79 :
		TR_248 = TR_29 ;
	7'h7a :
		TR_248 = TR_29 ;
	7'h7b :
		TR_248 = TR_29 ;
	7'h7c :
		TR_248 = TR_29 ;
	7'h7d :
		TR_248 = TR_29 ;
	7'h7e :
		TR_248 = TR_29 ;
	7'h7f :
		TR_248 = TR_29 ;
	default :
		TR_248 = 9'hx ;
	endcase
always @ ( TR_248 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_6 or 
	U_174 or RG_rl_137 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_17_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h11 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_17_t = ( ( { 9{ ST1_03d } } & RG_rl_137 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_6 )
		| ( { 9{ U_173 } } & TR_248 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_17_en = ( ST1_03d | U_174 | RG_rl_17_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_17_en )
		RG_rl_17 <= RG_rl_17_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_30 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_247 = TR_30 ;
	7'h01 :
		TR_247 = TR_30 ;
	7'h02 :
		TR_247 = TR_30 ;
	7'h03 :
		TR_247 = TR_30 ;
	7'h04 :
		TR_247 = TR_30 ;
	7'h05 :
		TR_247 = TR_30 ;
	7'h06 :
		TR_247 = TR_30 ;
	7'h07 :
		TR_247 = TR_30 ;
	7'h08 :
		TR_247 = TR_30 ;
	7'h09 :
		TR_247 = TR_30 ;
	7'h0a :
		TR_247 = TR_30 ;
	7'h0b :
		TR_247 = TR_30 ;
	7'h0c :
		TR_247 = TR_30 ;
	7'h0d :
		TR_247 = TR_30 ;
	7'h0e :
		TR_247 = TR_30 ;
	7'h0f :
		TR_247 = TR_30 ;
	7'h10 :
		TR_247 = TR_30 ;
	7'h11 :
		TR_247 = TR_30 ;
	7'h12 :
		TR_247 = 9'h000 ;	// line#=../rle.cpp:80
	7'h13 :
		TR_247 = TR_30 ;
	7'h14 :
		TR_247 = TR_30 ;
	7'h15 :
		TR_247 = TR_30 ;
	7'h16 :
		TR_247 = TR_30 ;
	7'h17 :
		TR_247 = TR_30 ;
	7'h18 :
		TR_247 = TR_30 ;
	7'h19 :
		TR_247 = TR_30 ;
	7'h1a :
		TR_247 = TR_30 ;
	7'h1b :
		TR_247 = TR_30 ;
	7'h1c :
		TR_247 = TR_30 ;
	7'h1d :
		TR_247 = TR_30 ;
	7'h1e :
		TR_247 = TR_30 ;
	7'h1f :
		TR_247 = TR_30 ;
	7'h20 :
		TR_247 = TR_30 ;
	7'h21 :
		TR_247 = TR_30 ;
	7'h22 :
		TR_247 = TR_30 ;
	7'h23 :
		TR_247 = TR_30 ;
	7'h24 :
		TR_247 = TR_30 ;
	7'h25 :
		TR_247 = TR_30 ;
	7'h26 :
		TR_247 = TR_30 ;
	7'h27 :
		TR_247 = TR_30 ;
	7'h28 :
		TR_247 = TR_30 ;
	7'h29 :
		TR_247 = TR_30 ;
	7'h2a :
		TR_247 = TR_30 ;
	7'h2b :
		TR_247 = TR_30 ;
	7'h2c :
		TR_247 = TR_30 ;
	7'h2d :
		TR_247 = TR_30 ;
	7'h2e :
		TR_247 = TR_30 ;
	7'h2f :
		TR_247 = TR_30 ;
	7'h30 :
		TR_247 = TR_30 ;
	7'h31 :
		TR_247 = TR_30 ;
	7'h32 :
		TR_247 = TR_30 ;
	7'h33 :
		TR_247 = TR_30 ;
	7'h34 :
		TR_247 = TR_30 ;
	7'h35 :
		TR_247 = TR_30 ;
	7'h36 :
		TR_247 = TR_30 ;
	7'h37 :
		TR_247 = TR_30 ;
	7'h38 :
		TR_247 = TR_30 ;
	7'h39 :
		TR_247 = TR_30 ;
	7'h3a :
		TR_247 = TR_30 ;
	7'h3b :
		TR_247 = TR_30 ;
	7'h3c :
		TR_247 = TR_30 ;
	7'h3d :
		TR_247 = TR_30 ;
	7'h3e :
		TR_247 = TR_30 ;
	7'h3f :
		TR_247 = TR_30 ;
	7'h40 :
		TR_247 = TR_30 ;
	7'h41 :
		TR_247 = TR_30 ;
	7'h42 :
		TR_247 = TR_30 ;
	7'h43 :
		TR_247 = TR_30 ;
	7'h44 :
		TR_247 = TR_30 ;
	7'h45 :
		TR_247 = TR_30 ;
	7'h46 :
		TR_247 = TR_30 ;
	7'h47 :
		TR_247 = TR_30 ;
	7'h48 :
		TR_247 = TR_30 ;
	7'h49 :
		TR_247 = TR_30 ;
	7'h4a :
		TR_247 = TR_30 ;
	7'h4b :
		TR_247 = TR_30 ;
	7'h4c :
		TR_247 = TR_30 ;
	7'h4d :
		TR_247 = TR_30 ;
	7'h4e :
		TR_247 = TR_30 ;
	7'h4f :
		TR_247 = TR_30 ;
	7'h50 :
		TR_247 = TR_30 ;
	7'h51 :
		TR_247 = TR_30 ;
	7'h52 :
		TR_247 = TR_30 ;
	7'h53 :
		TR_247 = TR_30 ;
	7'h54 :
		TR_247 = TR_30 ;
	7'h55 :
		TR_247 = TR_30 ;
	7'h56 :
		TR_247 = TR_30 ;
	7'h57 :
		TR_247 = TR_30 ;
	7'h58 :
		TR_247 = TR_30 ;
	7'h59 :
		TR_247 = TR_30 ;
	7'h5a :
		TR_247 = TR_30 ;
	7'h5b :
		TR_247 = TR_30 ;
	7'h5c :
		TR_247 = TR_30 ;
	7'h5d :
		TR_247 = TR_30 ;
	7'h5e :
		TR_247 = TR_30 ;
	7'h5f :
		TR_247 = TR_30 ;
	7'h60 :
		TR_247 = TR_30 ;
	7'h61 :
		TR_247 = TR_30 ;
	7'h62 :
		TR_247 = TR_30 ;
	7'h63 :
		TR_247 = TR_30 ;
	7'h64 :
		TR_247 = TR_30 ;
	7'h65 :
		TR_247 = TR_30 ;
	7'h66 :
		TR_247 = TR_30 ;
	7'h67 :
		TR_247 = TR_30 ;
	7'h68 :
		TR_247 = TR_30 ;
	7'h69 :
		TR_247 = TR_30 ;
	7'h6a :
		TR_247 = TR_30 ;
	7'h6b :
		TR_247 = TR_30 ;
	7'h6c :
		TR_247 = TR_30 ;
	7'h6d :
		TR_247 = TR_30 ;
	7'h6e :
		TR_247 = TR_30 ;
	7'h6f :
		TR_247 = TR_30 ;
	7'h70 :
		TR_247 = TR_30 ;
	7'h71 :
		TR_247 = TR_30 ;
	7'h72 :
		TR_247 = TR_30 ;
	7'h73 :
		TR_247 = TR_30 ;
	7'h74 :
		TR_247 = TR_30 ;
	7'h75 :
		TR_247 = TR_30 ;
	7'h76 :
		TR_247 = TR_30 ;
	7'h77 :
		TR_247 = TR_30 ;
	7'h78 :
		TR_247 = TR_30 ;
	7'h79 :
		TR_247 = TR_30 ;
	7'h7a :
		TR_247 = TR_30 ;
	7'h7b :
		TR_247 = TR_30 ;
	7'h7c :
		TR_247 = TR_30 ;
	7'h7d :
		TR_247 = TR_30 ;
	7'h7e :
		TR_247 = TR_30 ;
	7'h7f :
		TR_247 = TR_30 ;
	default :
		TR_247 = 9'hx ;
	endcase
always @ ( TR_247 or U_173 or sub8u_71ot or U_183 or RG_rl_138 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_18_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h12 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_18_t = ( ( { 9{ M_180 } } & RG_rl_138 )
		| ( { 9{ U_173 } } & TR_247 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_18_en = ( M_180 | RG_rl_18_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_18_en )
		RG_rl_18 <= RG_rl_18_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_31 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_246 = TR_31 ;
	7'h01 :
		TR_246 = TR_31 ;
	7'h02 :
		TR_246 = TR_31 ;
	7'h03 :
		TR_246 = TR_31 ;
	7'h04 :
		TR_246 = TR_31 ;
	7'h05 :
		TR_246 = TR_31 ;
	7'h06 :
		TR_246 = TR_31 ;
	7'h07 :
		TR_246 = TR_31 ;
	7'h08 :
		TR_246 = TR_31 ;
	7'h09 :
		TR_246 = TR_31 ;
	7'h0a :
		TR_246 = TR_31 ;
	7'h0b :
		TR_246 = TR_31 ;
	7'h0c :
		TR_246 = TR_31 ;
	7'h0d :
		TR_246 = TR_31 ;
	7'h0e :
		TR_246 = TR_31 ;
	7'h0f :
		TR_246 = TR_31 ;
	7'h10 :
		TR_246 = TR_31 ;
	7'h11 :
		TR_246 = TR_31 ;
	7'h12 :
		TR_246 = TR_31 ;
	7'h13 :
		TR_246 = 9'h000 ;	// line#=../rle.cpp:80
	7'h14 :
		TR_246 = TR_31 ;
	7'h15 :
		TR_246 = TR_31 ;
	7'h16 :
		TR_246 = TR_31 ;
	7'h17 :
		TR_246 = TR_31 ;
	7'h18 :
		TR_246 = TR_31 ;
	7'h19 :
		TR_246 = TR_31 ;
	7'h1a :
		TR_246 = TR_31 ;
	7'h1b :
		TR_246 = TR_31 ;
	7'h1c :
		TR_246 = TR_31 ;
	7'h1d :
		TR_246 = TR_31 ;
	7'h1e :
		TR_246 = TR_31 ;
	7'h1f :
		TR_246 = TR_31 ;
	7'h20 :
		TR_246 = TR_31 ;
	7'h21 :
		TR_246 = TR_31 ;
	7'h22 :
		TR_246 = TR_31 ;
	7'h23 :
		TR_246 = TR_31 ;
	7'h24 :
		TR_246 = TR_31 ;
	7'h25 :
		TR_246 = TR_31 ;
	7'h26 :
		TR_246 = TR_31 ;
	7'h27 :
		TR_246 = TR_31 ;
	7'h28 :
		TR_246 = TR_31 ;
	7'h29 :
		TR_246 = TR_31 ;
	7'h2a :
		TR_246 = TR_31 ;
	7'h2b :
		TR_246 = TR_31 ;
	7'h2c :
		TR_246 = TR_31 ;
	7'h2d :
		TR_246 = TR_31 ;
	7'h2e :
		TR_246 = TR_31 ;
	7'h2f :
		TR_246 = TR_31 ;
	7'h30 :
		TR_246 = TR_31 ;
	7'h31 :
		TR_246 = TR_31 ;
	7'h32 :
		TR_246 = TR_31 ;
	7'h33 :
		TR_246 = TR_31 ;
	7'h34 :
		TR_246 = TR_31 ;
	7'h35 :
		TR_246 = TR_31 ;
	7'h36 :
		TR_246 = TR_31 ;
	7'h37 :
		TR_246 = TR_31 ;
	7'h38 :
		TR_246 = TR_31 ;
	7'h39 :
		TR_246 = TR_31 ;
	7'h3a :
		TR_246 = TR_31 ;
	7'h3b :
		TR_246 = TR_31 ;
	7'h3c :
		TR_246 = TR_31 ;
	7'h3d :
		TR_246 = TR_31 ;
	7'h3e :
		TR_246 = TR_31 ;
	7'h3f :
		TR_246 = TR_31 ;
	7'h40 :
		TR_246 = TR_31 ;
	7'h41 :
		TR_246 = TR_31 ;
	7'h42 :
		TR_246 = TR_31 ;
	7'h43 :
		TR_246 = TR_31 ;
	7'h44 :
		TR_246 = TR_31 ;
	7'h45 :
		TR_246 = TR_31 ;
	7'h46 :
		TR_246 = TR_31 ;
	7'h47 :
		TR_246 = TR_31 ;
	7'h48 :
		TR_246 = TR_31 ;
	7'h49 :
		TR_246 = TR_31 ;
	7'h4a :
		TR_246 = TR_31 ;
	7'h4b :
		TR_246 = TR_31 ;
	7'h4c :
		TR_246 = TR_31 ;
	7'h4d :
		TR_246 = TR_31 ;
	7'h4e :
		TR_246 = TR_31 ;
	7'h4f :
		TR_246 = TR_31 ;
	7'h50 :
		TR_246 = TR_31 ;
	7'h51 :
		TR_246 = TR_31 ;
	7'h52 :
		TR_246 = TR_31 ;
	7'h53 :
		TR_246 = TR_31 ;
	7'h54 :
		TR_246 = TR_31 ;
	7'h55 :
		TR_246 = TR_31 ;
	7'h56 :
		TR_246 = TR_31 ;
	7'h57 :
		TR_246 = TR_31 ;
	7'h58 :
		TR_246 = TR_31 ;
	7'h59 :
		TR_246 = TR_31 ;
	7'h5a :
		TR_246 = TR_31 ;
	7'h5b :
		TR_246 = TR_31 ;
	7'h5c :
		TR_246 = TR_31 ;
	7'h5d :
		TR_246 = TR_31 ;
	7'h5e :
		TR_246 = TR_31 ;
	7'h5f :
		TR_246 = TR_31 ;
	7'h60 :
		TR_246 = TR_31 ;
	7'h61 :
		TR_246 = TR_31 ;
	7'h62 :
		TR_246 = TR_31 ;
	7'h63 :
		TR_246 = TR_31 ;
	7'h64 :
		TR_246 = TR_31 ;
	7'h65 :
		TR_246 = TR_31 ;
	7'h66 :
		TR_246 = TR_31 ;
	7'h67 :
		TR_246 = TR_31 ;
	7'h68 :
		TR_246 = TR_31 ;
	7'h69 :
		TR_246 = TR_31 ;
	7'h6a :
		TR_246 = TR_31 ;
	7'h6b :
		TR_246 = TR_31 ;
	7'h6c :
		TR_246 = TR_31 ;
	7'h6d :
		TR_246 = TR_31 ;
	7'h6e :
		TR_246 = TR_31 ;
	7'h6f :
		TR_246 = TR_31 ;
	7'h70 :
		TR_246 = TR_31 ;
	7'h71 :
		TR_246 = TR_31 ;
	7'h72 :
		TR_246 = TR_31 ;
	7'h73 :
		TR_246 = TR_31 ;
	7'h74 :
		TR_246 = TR_31 ;
	7'h75 :
		TR_246 = TR_31 ;
	7'h76 :
		TR_246 = TR_31 ;
	7'h77 :
		TR_246 = TR_31 ;
	7'h78 :
		TR_246 = TR_31 ;
	7'h79 :
		TR_246 = TR_31 ;
	7'h7a :
		TR_246 = TR_31 ;
	7'h7b :
		TR_246 = TR_31 ;
	7'h7c :
		TR_246 = TR_31 ;
	7'h7d :
		TR_246 = TR_31 ;
	7'h7e :
		TR_246 = TR_31 ;
	7'h7f :
		TR_246 = TR_31 ;
	default :
		TR_246 = 9'hx ;
	endcase
always @ ( TR_246 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_7 or 
	U_174 or RG_rl_138 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_19_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h13 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_19_t = ( ( { 9{ ST1_03d } } & RG_rl_138 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_7 )
		| ( { 9{ U_173 } } & TR_246 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_19_en = ( ST1_03d | U_174 | RG_rl_19_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_19_en )
		RG_rl_19 <= RG_rl_19_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_32 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_245 = TR_32 ;
	7'h01 :
		TR_245 = TR_32 ;
	7'h02 :
		TR_245 = TR_32 ;
	7'h03 :
		TR_245 = TR_32 ;
	7'h04 :
		TR_245 = TR_32 ;
	7'h05 :
		TR_245 = TR_32 ;
	7'h06 :
		TR_245 = TR_32 ;
	7'h07 :
		TR_245 = TR_32 ;
	7'h08 :
		TR_245 = TR_32 ;
	7'h09 :
		TR_245 = TR_32 ;
	7'h0a :
		TR_245 = TR_32 ;
	7'h0b :
		TR_245 = TR_32 ;
	7'h0c :
		TR_245 = TR_32 ;
	7'h0d :
		TR_245 = TR_32 ;
	7'h0e :
		TR_245 = TR_32 ;
	7'h0f :
		TR_245 = TR_32 ;
	7'h10 :
		TR_245 = TR_32 ;
	7'h11 :
		TR_245 = TR_32 ;
	7'h12 :
		TR_245 = TR_32 ;
	7'h13 :
		TR_245 = TR_32 ;
	7'h14 :
		TR_245 = 9'h000 ;	// line#=../rle.cpp:80
	7'h15 :
		TR_245 = TR_32 ;
	7'h16 :
		TR_245 = TR_32 ;
	7'h17 :
		TR_245 = TR_32 ;
	7'h18 :
		TR_245 = TR_32 ;
	7'h19 :
		TR_245 = TR_32 ;
	7'h1a :
		TR_245 = TR_32 ;
	7'h1b :
		TR_245 = TR_32 ;
	7'h1c :
		TR_245 = TR_32 ;
	7'h1d :
		TR_245 = TR_32 ;
	7'h1e :
		TR_245 = TR_32 ;
	7'h1f :
		TR_245 = TR_32 ;
	7'h20 :
		TR_245 = TR_32 ;
	7'h21 :
		TR_245 = TR_32 ;
	7'h22 :
		TR_245 = TR_32 ;
	7'h23 :
		TR_245 = TR_32 ;
	7'h24 :
		TR_245 = TR_32 ;
	7'h25 :
		TR_245 = TR_32 ;
	7'h26 :
		TR_245 = TR_32 ;
	7'h27 :
		TR_245 = TR_32 ;
	7'h28 :
		TR_245 = TR_32 ;
	7'h29 :
		TR_245 = TR_32 ;
	7'h2a :
		TR_245 = TR_32 ;
	7'h2b :
		TR_245 = TR_32 ;
	7'h2c :
		TR_245 = TR_32 ;
	7'h2d :
		TR_245 = TR_32 ;
	7'h2e :
		TR_245 = TR_32 ;
	7'h2f :
		TR_245 = TR_32 ;
	7'h30 :
		TR_245 = TR_32 ;
	7'h31 :
		TR_245 = TR_32 ;
	7'h32 :
		TR_245 = TR_32 ;
	7'h33 :
		TR_245 = TR_32 ;
	7'h34 :
		TR_245 = TR_32 ;
	7'h35 :
		TR_245 = TR_32 ;
	7'h36 :
		TR_245 = TR_32 ;
	7'h37 :
		TR_245 = TR_32 ;
	7'h38 :
		TR_245 = TR_32 ;
	7'h39 :
		TR_245 = TR_32 ;
	7'h3a :
		TR_245 = TR_32 ;
	7'h3b :
		TR_245 = TR_32 ;
	7'h3c :
		TR_245 = TR_32 ;
	7'h3d :
		TR_245 = TR_32 ;
	7'h3e :
		TR_245 = TR_32 ;
	7'h3f :
		TR_245 = TR_32 ;
	7'h40 :
		TR_245 = TR_32 ;
	7'h41 :
		TR_245 = TR_32 ;
	7'h42 :
		TR_245 = TR_32 ;
	7'h43 :
		TR_245 = TR_32 ;
	7'h44 :
		TR_245 = TR_32 ;
	7'h45 :
		TR_245 = TR_32 ;
	7'h46 :
		TR_245 = TR_32 ;
	7'h47 :
		TR_245 = TR_32 ;
	7'h48 :
		TR_245 = TR_32 ;
	7'h49 :
		TR_245 = TR_32 ;
	7'h4a :
		TR_245 = TR_32 ;
	7'h4b :
		TR_245 = TR_32 ;
	7'h4c :
		TR_245 = TR_32 ;
	7'h4d :
		TR_245 = TR_32 ;
	7'h4e :
		TR_245 = TR_32 ;
	7'h4f :
		TR_245 = TR_32 ;
	7'h50 :
		TR_245 = TR_32 ;
	7'h51 :
		TR_245 = TR_32 ;
	7'h52 :
		TR_245 = TR_32 ;
	7'h53 :
		TR_245 = TR_32 ;
	7'h54 :
		TR_245 = TR_32 ;
	7'h55 :
		TR_245 = TR_32 ;
	7'h56 :
		TR_245 = TR_32 ;
	7'h57 :
		TR_245 = TR_32 ;
	7'h58 :
		TR_245 = TR_32 ;
	7'h59 :
		TR_245 = TR_32 ;
	7'h5a :
		TR_245 = TR_32 ;
	7'h5b :
		TR_245 = TR_32 ;
	7'h5c :
		TR_245 = TR_32 ;
	7'h5d :
		TR_245 = TR_32 ;
	7'h5e :
		TR_245 = TR_32 ;
	7'h5f :
		TR_245 = TR_32 ;
	7'h60 :
		TR_245 = TR_32 ;
	7'h61 :
		TR_245 = TR_32 ;
	7'h62 :
		TR_245 = TR_32 ;
	7'h63 :
		TR_245 = TR_32 ;
	7'h64 :
		TR_245 = TR_32 ;
	7'h65 :
		TR_245 = TR_32 ;
	7'h66 :
		TR_245 = TR_32 ;
	7'h67 :
		TR_245 = TR_32 ;
	7'h68 :
		TR_245 = TR_32 ;
	7'h69 :
		TR_245 = TR_32 ;
	7'h6a :
		TR_245 = TR_32 ;
	7'h6b :
		TR_245 = TR_32 ;
	7'h6c :
		TR_245 = TR_32 ;
	7'h6d :
		TR_245 = TR_32 ;
	7'h6e :
		TR_245 = TR_32 ;
	7'h6f :
		TR_245 = TR_32 ;
	7'h70 :
		TR_245 = TR_32 ;
	7'h71 :
		TR_245 = TR_32 ;
	7'h72 :
		TR_245 = TR_32 ;
	7'h73 :
		TR_245 = TR_32 ;
	7'h74 :
		TR_245 = TR_32 ;
	7'h75 :
		TR_245 = TR_32 ;
	7'h76 :
		TR_245 = TR_32 ;
	7'h77 :
		TR_245 = TR_32 ;
	7'h78 :
		TR_245 = TR_32 ;
	7'h79 :
		TR_245 = TR_32 ;
	7'h7a :
		TR_245 = TR_32 ;
	7'h7b :
		TR_245 = TR_32 ;
	7'h7c :
		TR_245 = TR_32 ;
	7'h7d :
		TR_245 = TR_32 ;
	7'h7e :
		TR_245 = TR_32 ;
	7'h7f :
		TR_245 = TR_32 ;
	default :
		TR_245 = 9'hx ;
	endcase
always @ ( TR_245 or U_173 or sub8u_71ot or U_183 or RG_rl_139 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_20_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h14 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_20_t = ( ( { 9{ M_180 } } & RG_rl_139 )
		| ( { 9{ U_173 } } & TR_245 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_20_en = ( M_180 | RG_rl_20_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_20_en )
		RG_rl_20 <= RG_rl_20_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_33 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_244 = TR_33 ;
	7'h01 :
		TR_244 = TR_33 ;
	7'h02 :
		TR_244 = TR_33 ;
	7'h03 :
		TR_244 = TR_33 ;
	7'h04 :
		TR_244 = TR_33 ;
	7'h05 :
		TR_244 = TR_33 ;
	7'h06 :
		TR_244 = TR_33 ;
	7'h07 :
		TR_244 = TR_33 ;
	7'h08 :
		TR_244 = TR_33 ;
	7'h09 :
		TR_244 = TR_33 ;
	7'h0a :
		TR_244 = TR_33 ;
	7'h0b :
		TR_244 = TR_33 ;
	7'h0c :
		TR_244 = TR_33 ;
	7'h0d :
		TR_244 = TR_33 ;
	7'h0e :
		TR_244 = TR_33 ;
	7'h0f :
		TR_244 = TR_33 ;
	7'h10 :
		TR_244 = TR_33 ;
	7'h11 :
		TR_244 = TR_33 ;
	7'h12 :
		TR_244 = TR_33 ;
	7'h13 :
		TR_244 = TR_33 ;
	7'h14 :
		TR_244 = TR_33 ;
	7'h15 :
		TR_244 = 9'h000 ;	// line#=../rle.cpp:80
	7'h16 :
		TR_244 = TR_33 ;
	7'h17 :
		TR_244 = TR_33 ;
	7'h18 :
		TR_244 = TR_33 ;
	7'h19 :
		TR_244 = TR_33 ;
	7'h1a :
		TR_244 = TR_33 ;
	7'h1b :
		TR_244 = TR_33 ;
	7'h1c :
		TR_244 = TR_33 ;
	7'h1d :
		TR_244 = TR_33 ;
	7'h1e :
		TR_244 = TR_33 ;
	7'h1f :
		TR_244 = TR_33 ;
	7'h20 :
		TR_244 = TR_33 ;
	7'h21 :
		TR_244 = TR_33 ;
	7'h22 :
		TR_244 = TR_33 ;
	7'h23 :
		TR_244 = TR_33 ;
	7'h24 :
		TR_244 = TR_33 ;
	7'h25 :
		TR_244 = TR_33 ;
	7'h26 :
		TR_244 = TR_33 ;
	7'h27 :
		TR_244 = TR_33 ;
	7'h28 :
		TR_244 = TR_33 ;
	7'h29 :
		TR_244 = TR_33 ;
	7'h2a :
		TR_244 = TR_33 ;
	7'h2b :
		TR_244 = TR_33 ;
	7'h2c :
		TR_244 = TR_33 ;
	7'h2d :
		TR_244 = TR_33 ;
	7'h2e :
		TR_244 = TR_33 ;
	7'h2f :
		TR_244 = TR_33 ;
	7'h30 :
		TR_244 = TR_33 ;
	7'h31 :
		TR_244 = TR_33 ;
	7'h32 :
		TR_244 = TR_33 ;
	7'h33 :
		TR_244 = TR_33 ;
	7'h34 :
		TR_244 = TR_33 ;
	7'h35 :
		TR_244 = TR_33 ;
	7'h36 :
		TR_244 = TR_33 ;
	7'h37 :
		TR_244 = TR_33 ;
	7'h38 :
		TR_244 = TR_33 ;
	7'h39 :
		TR_244 = TR_33 ;
	7'h3a :
		TR_244 = TR_33 ;
	7'h3b :
		TR_244 = TR_33 ;
	7'h3c :
		TR_244 = TR_33 ;
	7'h3d :
		TR_244 = TR_33 ;
	7'h3e :
		TR_244 = TR_33 ;
	7'h3f :
		TR_244 = TR_33 ;
	7'h40 :
		TR_244 = TR_33 ;
	7'h41 :
		TR_244 = TR_33 ;
	7'h42 :
		TR_244 = TR_33 ;
	7'h43 :
		TR_244 = TR_33 ;
	7'h44 :
		TR_244 = TR_33 ;
	7'h45 :
		TR_244 = TR_33 ;
	7'h46 :
		TR_244 = TR_33 ;
	7'h47 :
		TR_244 = TR_33 ;
	7'h48 :
		TR_244 = TR_33 ;
	7'h49 :
		TR_244 = TR_33 ;
	7'h4a :
		TR_244 = TR_33 ;
	7'h4b :
		TR_244 = TR_33 ;
	7'h4c :
		TR_244 = TR_33 ;
	7'h4d :
		TR_244 = TR_33 ;
	7'h4e :
		TR_244 = TR_33 ;
	7'h4f :
		TR_244 = TR_33 ;
	7'h50 :
		TR_244 = TR_33 ;
	7'h51 :
		TR_244 = TR_33 ;
	7'h52 :
		TR_244 = TR_33 ;
	7'h53 :
		TR_244 = TR_33 ;
	7'h54 :
		TR_244 = TR_33 ;
	7'h55 :
		TR_244 = TR_33 ;
	7'h56 :
		TR_244 = TR_33 ;
	7'h57 :
		TR_244 = TR_33 ;
	7'h58 :
		TR_244 = TR_33 ;
	7'h59 :
		TR_244 = TR_33 ;
	7'h5a :
		TR_244 = TR_33 ;
	7'h5b :
		TR_244 = TR_33 ;
	7'h5c :
		TR_244 = TR_33 ;
	7'h5d :
		TR_244 = TR_33 ;
	7'h5e :
		TR_244 = TR_33 ;
	7'h5f :
		TR_244 = TR_33 ;
	7'h60 :
		TR_244 = TR_33 ;
	7'h61 :
		TR_244 = TR_33 ;
	7'h62 :
		TR_244 = TR_33 ;
	7'h63 :
		TR_244 = TR_33 ;
	7'h64 :
		TR_244 = TR_33 ;
	7'h65 :
		TR_244 = TR_33 ;
	7'h66 :
		TR_244 = TR_33 ;
	7'h67 :
		TR_244 = TR_33 ;
	7'h68 :
		TR_244 = TR_33 ;
	7'h69 :
		TR_244 = TR_33 ;
	7'h6a :
		TR_244 = TR_33 ;
	7'h6b :
		TR_244 = TR_33 ;
	7'h6c :
		TR_244 = TR_33 ;
	7'h6d :
		TR_244 = TR_33 ;
	7'h6e :
		TR_244 = TR_33 ;
	7'h6f :
		TR_244 = TR_33 ;
	7'h70 :
		TR_244 = TR_33 ;
	7'h71 :
		TR_244 = TR_33 ;
	7'h72 :
		TR_244 = TR_33 ;
	7'h73 :
		TR_244 = TR_33 ;
	7'h74 :
		TR_244 = TR_33 ;
	7'h75 :
		TR_244 = TR_33 ;
	7'h76 :
		TR_244 = TR_33 ;
	7'h77 :
		TR_244 = TR_33 ;
	7'h78 :
		TR_244 = TR_33 ;
	7'h79 :
		TR_244 = TR_33 ;
	7'h7a :
		TR_244 = TR_33 ;
	7'h7b :
		TR_244 = TR_33 ;
	7'h7c :
		TR_244 = TR_33 ;
	7'h7d :
		TR_244 = TR_33 ;
	7'h7e :
		TR_244 = TR_33 ;
	7'h7f :
		TR_244 = TR_33 ;
	default :
		TR_244 = 9'hx ;
	endcase
always @ ( TR_244 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_8 or 
	U_174 or RG_rl_139 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_21_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h15 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_21_t = ( ( { 9{ ST1_03d } } & RG_rl_139 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_8 )
		| ( { 9{ U_173 } } & TR_244 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_21_en = ( ST1_03d | U_174 | RG_rl_21_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_21_en )
		RG_rl_21 <= RG_rl_21_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_34 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_243 = TR_34 ;
	7'h01 :
		TR_243 = TR_34 ;
	7'h02 :
		TR_243 = TR_34 ;
	7'h03 :
		TR_243 = TR_34 ;
	7'h04 :
		TR_243 = TR_34 ;
	7'h05 :
		TR_243 = TR_34 ;
	7'h06 :
		TR_243 = TR_34 ;
	7'h07 :
		TR_243 = TR_34 ;
	7'h08 :
		TR_243 = TR_34 ;
	7'h09 :
		TR_243 = TR_34 ;
	7'h0a :
		TR_243 = TR_34 ;
	7'h0b :
		TR_243 = TR_34 ;
	7'h0c :
		TR_243 = TR_34 ;
	7'h0d :
		TR_243 = TR_34 ;
	7'h0e :
		TR_243 = TR_34 ;
	7'h0f :
		TR_243 = TR_34 ;
	7'h10 :
		TR_243 = TR_34 ;
	7'h11 :
		TR_243 = TR_34 ;
	7'h12 :
		TR_243 = TR_34 ;
	7'h13 :
		TR_243 = TR_34 ;
	7'h14 :
		TR_243 = TR_34 ;
	7'h15 :
		TR_243 = TR_34 ;
	7'h16 :
		TR_243 = 9'h000 ;	// line#=../rle.cpp:80
	7'h17 :
		TR_243 = TR_34 ;
	7'h18 :
		TR_243 = TR_34 ;
	7'h19 :
		TR_243 = TR_34 ;
	7'h1a :
		TR_243 = TR_34 ;
	7'h1b :
		TR_243 = TR_34 ;
	7'h1c :
		TR_243 = TR_34 ;
	7'h1d :
		TR_243 = TR_34 ;
	7'h1e :
		TR_243 = TR_34 ;
	7'h1f :
		TR_243 = TR_34 ;
	7'h20 :
		TR_243 = TR_34 ;
	7'h21 :
		TR_243 = TR_34 ;
	7'h22 :
		TR_243 = TR_34 ;
	7'h23 :
		TR_243 = TR_34 ;
	7'h24 :
		TR_243 = TR_34 ;
	7'h25 :
		TR_243 = TR_34 ;
	7'h26 :
		TR_243 = TR_34 ;
	7'h27 :
		TR_243 = TR_34 ;
	7'h28 :
		TR_243 = TR_34 ;
	7'h29 :
		TR_243 = TR_34 ;
	7'h2a :
		TR_243 = TR_34 ;
	7'h2b :
		TR_243 = TR_34 ;
	7'h2c :
		TR_243 = TR_34 ;
	7'h2d :
		TR_243 = TR_34 ;
	7'h2e :
		TR_243 = TR_34 ;
	7'h2f :
		TR_243 = TR_34 ;
	7'h30 :
		TR_243 = TR_34 ;
	7'h31 :
		TR_243 = TR_34 ;
	7'h32 :
		TR_243 = TR_34 ;
	7'h33 :
		TR_243 = TR_34 ;
	7'h34 :
		TR_243 = TR_34 ;
	7'h35 :
		TR_243 = TR_34 ;
	7'h36 :
		TR_243 = TR_34 ;
	7'h37 :
		TR_243 = TR_34 ;
	7'h38 :
		TR_243 = TR_34 ;
	7'h39 :
		TR_243 = TR_34 ;
	7'h3a :
		TR_243 = TR_34 ;
	7'h3b :
		TR_243 = TR_34 ;
	7'h3c :
		TR_243 = TR_34 ;
	7'h3d :
		TR_243 = TR_34 ;
	7'h3e :
		TR_243 = TR_34 ;
	7'h3f :
		TR_243 = TR_34 ;
	7'h40 :
		TR_243 = TR_34 ;
	7'h41 :
		TR_243 = TR_34 ;
	7'h42 :
		TR_243 = TR_34 ;
	7'h43 :
		TR_243 = TR_34 ;
	7'h44 :
		TR_243 = TR_34 ;
	7'h45 :
		TR_243 = TR_34 ;
	7'h46 :
		TR_243 = TR_34 ;
	7'h47 :
		TR_243 = TR_34 ;
	7'h48 :
		TR_243 = TR_34 ;
	7'h49 :
		TR_243 = TR_34 ;
	7'h4a :
		TR_243 = TR_34 ;
	7'h4b :
		TR_243 = TR_34 ;
	7'h4c :
		TR_243 = TR_34 ;
	7'h4d :
		TR_243 = TR_34 ;
	7'h4e :
		TR_243 = TR_34 ;
	7'h4f :
		TR_243 = TR_34 ;
	7'h50 :
		TR_243 = TR_34 ;
	7'h51 :
		TR_243 = TR_34 ;
	7'h52 :
		TR_243 = TR_34 ;
	7'h53 :
		TR_243 = TR_34 ;
	7'h54 :
		TR_243 = TR_34 ;
	7'h55 :
		TR_243 = TR_34 ;
	7'h56 :
		TR_243 = TR_34 ;
	7'h57 :
		TR_243 = TR_34 ;
	7'h58 :
		TR_243 = TR_34 ;
	7'h59 :
		TR_243 = TR_34 ;
	7'h5a :
		TR_243 = TR_34 ;
	7'h5b :
		TR_243 = TR_34 ;
	7'h5c :
		TR_243 = TR_34 ;
	7'h5d :
		TR_243 = TR_34 ;
	7'h5e :
		TR_243 = TR_34 ;
	7'h5f :
		TR_243 = TR_34 ;
	7'h60 :
		TR_243 = TR_34 ;
	7'h61 :
		TR_243 = TR_34 ;
	7'h62 :
		TR_243 = TR_34 ;
	7'h63 :
		TR_243 = TR_34 ;
	7'h64 :
		TR_243 = TR_34 ;
	7'h65 :
		TR_243 = TR_34 ;
	7'h66 :
		TR_243 = TR_34 ;
	7'h67 :
		TR_243 = TR_34 ;
	7'h68 :
		TR_243 = TR_34 ;
	7'h69 :
		TR_243 = TR_34 ;
	7'h6a :
		TR_243 = TR_34 ;
	7'h6b :
		TR_243 = TR_34 ;
	7'h6c :
		TR_243 = TR_34 ;
	7'h6d :
		TR_243 = TR_34 ;
	7'h6e :
		TR_243 = TR_34 ;
	7'h6f :
		TR_243 = TR_34 ;
	7'h70 :
		TR_243 = TR_34 ;
	7'h71 :
		TR_243 = TR_34 ;
	7'h72 :
		TR_243 = TR_34 ;
	7'h73 :
		TR_243 = TR_34 ;
	7'h74 :
		TR_243 = TR_34 ;
	7'h75 :
		TR_243 = TR_34 ;
	7'h76 :
		TR_243 = TR_34 ;
	7'h77 :
		TR_243 = TR_34 ;
	7'h78 :
		TR_243 = TR_34 ;
	7'h79 :
		TR_243 = TR_34 ;
	7'h7a :
		TR_243 = TR_34 ;
	7'h7b :
		TR_243 = TR_34 ;
	7'h7c :
		TR_243 = TR_34 ;
	7'h7d :
		TR_243 = TR_34 ;
	7'h7e :
		TR_243 = TR_34 ;
	7'h7f :
		TR_243 = TR_34 ;
	default :
		TR_243 = 9'hx ;
	endcase
always @ ( TR_243 or U_173 or sub8u_71ot or U_183 or RG_rl_140 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_22_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h16 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_22_t = ( ( { 9{ M_180 } } & RG_rl_140 )
		| ( { 9{ U_173 } } & TR_243 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_22_en = ( M_180 | RG_rl_22_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_22_en )
		RG_rl_22 <= RG_rl_22_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_35 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_242 = TR_35 ;
	7'h01 :
		TR_242 = TR_35 ;
	7'h02 :
		TR_242 = TR_35 ;
	7'h03 :
		TR_242 = TR_35 ;
	7'h04 :
		TR_242 = TR_35 ;
	7'h05 :
		TR_242 = TR_35 ;
	7'h06 :
		TR_242 = TR_35 ;
	7'h07 :
		TR_242 = TR_35 ;
	7'h08 :
		TR_242 = TR_35 ;
	7'h09 :
		TR_242 = TR_35 ;
	7'h0a :
		TR_242 = TR_35 ;
	7'h0b :
		TR_242 = TR_35 ;
	7'h0c :
		TR_242 = TR_35 ;
	7'h0d :
		TR_242 = TR_35 ;
	7'h0e :
		TR_242 = TR_35 ;
	7'h0f :
		TR_242 = TR_35 ;
	7'h10 :
		TR_242 = TR_35 ;
	7'h11 :
		TR_242 = TR_35 ;
	7'h12 :
		TR_242 = TR_35 ;
	7'h13 :
		TR_242 = TR_35 ;
	7'h14 :
		TR_242 = TR_35 ;
	7'h15 :
		TR_242 = TR_35 ;
	7'h16 :
		TR_242 = TR_35 ;
	7'h17 :
		TR_242 = 9'h000 ;	// line#=../rle.cpp:80
	7'h18 :
		TR_242 = TR_35 ;
	7'h19 :
		TR_242 = TR_35 ;
	7'h1a :
		TR_242 = TR_35 ;
	7'h1b :
		TR_242 = TR_35 ;
	7'h1c :
		TR_242 = TR_35 ;
	7'h1d :
		TR_242 = TR_35 ;
	7'h1e :
		TR_242 = TR_35 ;
	7'h1f :
		TR_242 = TR_35 ;
	7'h20 :
		TR_242 = TR_35 ;
	7'h21 :
		TR_242 = TR_35 ;
	7'h22 :
		TR_242 = TR_35 ;
	7'h23 :
		TR_242 = TR_35 ;
	7'h24 :
		TR_242 = TR_35 ;
	7'h25 :
		TR_242 = TR_35 ;
	7'h26 :
		TR_242 = TR_35 ;
	7'h27 :
		TR_242 = TR_35 ;
	7'h28 :
		TR_242 = TR_35 ;
	7'h29 :
		TR_242 = TR_35 ;
	7'h2a :
		TR_242 = TR_35 ;
	7'h2b :
		TR_242 = TR_35 ;
	7'h2c :
		TR_242 = TR_35 ;
	7'h2d :
		TR_242 = TR_35 ;
	7'h2e :
		TR_242 = TR_35 ;
	7'h2f :
		TR_242 = TR_35 ;
	7'h30 :
		TR_242 = TR_35 ;
	7'h31 :
		TR_242 = TR_35 ;
	7'h32 :
		TR_242 = TR_35 ;
	7'h33 :
		TR_242 = TR_35 ;
	7'h34 :
		TR_242 = TR_35 ;
	7'h35 :
		TR_242 = TR_35 ;
	7'h36 :
		TR_242 = TR_35 ;
	7'h37 :
		TR_242 = TR_35 ;
	7'h38 :
		TR_242 = TR_35 ;
	7'h39 :
		TR_242 = TR_35 ;
	7'h3a :
		TR_242 = TR_35 ;
	7'h3b :
		TR_242 = TR_35 ;
	7'h3c :
		TR_242 = TR_35 ;
	7'h3d :
		TR_242 = TR_35 ;
	7'h3e :
		TR_242 = TR_35 ;
	7'h3f :
		TR_242 = TR_35 ;
	7'h40 :
		TR_242 = TR_35 ;
	7'h41 :
		TR_242 = TR_35 ;
	7'h42 :
		TR_242 = TR_35 ;
	7'h43 :
		TR_242 = TR_35 ;
	7'h44 :
		TR_242 = TR_35 ;
	7'h45 :
		TR_242 = TR_35 ;
	7'h46 :
		TR_242 = TR_35 ;
	7'h47 :
		TR_242 = TR_35 ;
	7'h48 :
		TR_242 = TR_35 ;
	7'h49 :
		TR_242 = TR_35 ;
	7'h4a :
		TR_242 = TR_35 ;
	7'h4b :
		TR_242 = TR_35 ;
	7'h4c :
		TR_242 = TR_35 ;
	7'h4d :
		TR_242 = TR_35 ;
	7'h4e :
		TR_242 = TR_35 ;
	7'h4f :
		TR_242 = TR_35 ;
	7'h50 :
		TR_242 = TR_35 ;
	7'h51 :
		TR_242 = TR_35 ;
	7'h52 :
		TR_242 = TR_35 ;
	7'h53 :
		TR_242 = TR_35 ;
	7'h54 :
		TR_242 = TR_35 ;
	7'h55 :
		TR_242 = TR_35 ;
	7'h56 :
		TR_242 = TR_35 ;
	7'h57 :
		TR_242 = TR_35 ;
	7'h58 :
		TR_242 = TR_35 ;
	7'h59 :
		TR_242 = TR_35 ;
	7'h5a :
		TR_242 = TR_35 ;
	7'h5b :
		TR_242 = TR_35 ;
	7'h5c :
		TR_242 = TR_35 ;
	7'h5d :
		TR_242 = TR_35 ;
	7'h5e :
		TR_242 = TR_35 ;
	7'h5f :
		TR_242 = TR_35 ;
	7'h60 :
		TR_242 = TR_35 ;
	7'h61 :
		TR_242 = TR_35 ;
	7'h62 :
		TR_242 = TR_35 ;
	7'h63 :
		TR_242 = TR_35 ;
	7'h64 :
		TR_242 = TR_35 ;
	7'h65 :
		TR_242 = TR_35 ;
	7'h66 :
		TR_242 = TR_35 ;
	7'h67 :
		TR_242 = TR_35 ;
	7'h68 :
		TR_242 = TR_35 ;
	7'h69 :
		TR_242 = TR_35 ;
	7'h6a :
		TR_242 = TR_35 ;
	7'h6b :
		TR_242 = TR_35 ;
	7'h6c :
		TR_242 = TR_35 ;
	7'h6d :
		TR_242 = TR_35 ;
	7'h6e :
		TR_242 = TR_35 ;
	7'h6f :
		TR_242 = TR_35 ;
	7'h70 :
		TR_242 = TR_35 ;
	7'h71 :
		TR_242 = TR_35 ;
	7'h72 :
		TR_242 = TR_35 ;
	7'h73 :
		TR_242 = TR_35 ;
	7'h74 :
		TR_242 = TR_35 ;
	7'h75 :
		TR_242 = TR_35 ;
	7'h76 :
		TR_242 = TR_35 ;
	7'h77 :
		TR_242 = TR_35 ;
	7'h78 :
		TR_242 = TR_35 ;
	7'h79 :
		TR_242 = TR_35 ;
	7'h7a :
		TR_242 = TR_35 ;
	7'h7b :
		TR_242 = TR_35 ;
	7'h7c :
		TR_242 = TR_35 ;
	7'h7d :
		TR_242 = TR_35 ;
	7'h7e :
		TR_242 = TR_35 ;
	7'h7f :
		TR_242 = TR_35 ;
	default :
		TR_242 = 9'hx ;
	endcase
always @ ( TR_242 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_9 or 
	U_174 or RG_rl_140 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_23_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h17 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_23_t = ( ( { 9{ ST1_03d } } & RG_rl_140 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_9 )
		| ( { 9{ U_173 } } & TR_242 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_23_en = ( ST1_03d | U_174 | RG_rl_23_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_23_en )
		RG_rl_23 <= RG_rl_23_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_36 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_241 = TR_36 ;
	7'h01 :
		TR_241 = TR_36 ;
	7'h02 :
		TR_241 = TR_36 ;
	7'h03 :
		TR_241 = TR_36 ;
	7'h04 :
		TR_241 = TR_36 ;
	7'h05 :
		TR_241 = TR_36 ;
	7'h06 :
		TR_241 = TR_36 ;
	7'h07 :
		TR_241 = TR_36 ;
	7'h08 :
		TR_241 = TR_36 ;
	7'h09 :
		TR_241 = TR_36 ;
	7'h0a :
		TR_241 = TR_36 ;
	7'h0b :
		TR_241 = TR_36 ;
	7'h0c :
		TR_241 = TR_36 ;
	7'h0d :
		TR_241 = TR_36 ;
	7'h0e :
		TR_241 = TR_36 ;
	7'h0f :
		TR_241 = TR_36 ;
	7'h10 :
		TR_241 = TR_36 ;
	7'h11 :
		TR_241 = TR_36 ;
	7'h12 :
		TR_241 = TR_36 ;
	7'h13 :
		TR_241 = TR_36 ;
	7'h14 :
		TR_241 = TR_36 ;
	7'h15 :
		TR_241 = TR_36 ;
	7'h16 :
		TR_241 = TR_36 ;
	7'h17 :
		TR_241 = TR_36 ;
	7'h18 :
		TR_241 = 9'h000 ;	// line#=../rle.cpp:80
	7'h19 :
		TR_241 = TR_36 ;
	7'h1a :
		TR_241 = TR_36 ;
	7'h1b :
		TR_241 = TR_36 ;
	7'h1c :
		TR_241 = TR_36 ;
	7'h1d :
		TR_241 = TR_36 ;
	7'h1e :
		TR_241 = TR_36 ;
	7'h1f :
		TR_241 = TR_36 ;
	7'h20 :
		TR_241 = TR_36 ;
	7'h21 :
		TR_241 = TR_36 ;
	7'h22 :
		TR_241 = TR_36 ;
	7'h23 :
		TR_241 = TR_36 ;
	7'h24 :
		TR_241 = TR_36 ;
	7'h25 :
		TR_241 = TR_36 ;
	7'h26 :
		TR_241 = TR_36 ;
	7'h27 :
		TR_241 = TR_36 ;
	7'h28 :
		TR_241 = TR_36 ;
	7'h29 :
		TR_241 = TR_36 ;
	7'h2a :
		TR_241 = TR_36 ;
	7'h2b :
		TR_241 = TR_36 ;
	7'h2c :
		TR_241 = TR_36 ;
	7'h2d :
		TR_241 = TR_36 ;
	7'h2e :
		TR_241 = TR_36 ;
	7'h2f :
		TR_241 = TR_36 ;
	7'h30 :
		TR_241 = TR_36 ;
	7'h31 :
		TR_241 = TR_36 ;
	7'h32 :
		TR_241 = TR_36 ;
	7'h33 :
		TR_241 = TR_36 ;
	7'h34 :
		TR_241 = TR_36 ;
	7'h35 :
		TR_241 = TR_36 ;
	7'h36 :
		TR_241 = TR_36 ;
	7'h37 :
		TR_241 = TR_36 ;
	7'h38 :
		TR_241 = TR_36 ;
	7'h39 :
		TR_241 = TR_36 ;
	7'h3a :
		TR_241 = TR_36 ;
	7'h3b :
		TR_241 = TR_36 ;
	7'h3c :
		TR_241 = TR_36 ;
	7'h3d :
		TR_241 = TR_36 ;
	7'h3e :
		TR_241 = TR_36 ;
	7'h3f :
		TR_241 = TR_36 ;
	7'h40 :
		TR_241 = TR_36 ;
	7'h41 :
		TR_241 = TR_36 ;
	7'h42 :
		TR_241 = TR_36 ;
	7'h43 :
		TR_241 = TR_36 ;
	7'h44 :
		TR_241 = TR_36 ;
	7'h45 :
		TR_241 = TR_36 ;
	7'h46 :
		TR_241 = TR_36 ;
	7'h47 :
		TR_241 = TR_36 ;
	7'h48 :
		TR_241 = TR_36 ;
	7'h49 :
		TR_241 = TR_36 ;
	7'h4a :
		TR_241 = TR_36 ;
	7'h4b :
		TR_241 = TR_36 ;
	7'h4c :
		TR_241 = TR_36 ;
	7'h4d :
		TR_241 = TR_36 ;
	7'h4e :
		TR_241 = TR_36 ;
	7'h4f :
		TR_241 = TR_36 ;
	7'h50 :
		TR_241 = TR_36 ;
	7'h51 :
		TR_241 = TR_36 ;
	7'h52 :
		TR_241 = TR_36 ;
	7'h53 :
		TR_241 = TR_36 ;
	7'h54 :
		TR_241 = TR_36 ;
	7'h55 :
		TR_241 = TR_36 ;
	7'h56 :
		TR_241 = TR_36 ;
	7'h57 :
		TR_241 = TR_36 ;
	7'h58 :
		TR_241 = TR_36 ;
	7'h59 :
		TR_241 = TR_36 ;
	7'h5a :
		TR_241 = TR_36 ;
	7'h5b :
		TR_241 = TR_36 ;
	7'h5c :
		TR_241 = TR_36 ;
	7'h5d :
		TR_241 = TR_36 ;
	7'h5e :
		TR_241 = TR_36 ;
	7'h5f :
		TR_241 = TR_36 ;
	7'h60 :
		TR_241 = TR_36 ;
	7'h61 :
		TR_241 = TR_36 ;
	7'h62 :
		TR_241 = TR_36 ;
	7'h63 :
		TR_241 = TR_36 ;
	7'h64 :
		TR_241 = TR_36 ;
	7'h65 :
		TR_241 = TR_36 ;
	7'h66 :
		TR_241 = TR_36 ;
	7'h67 :
		TR_241 = TR_36 ;
	7'h68 :
		TR_241 = TR_36 ;
	7'h69 :
		TR_241 = TR_36 ;
	7'h6a :
		TR_241 = TR_36 ;
	7'h6b :
		TR_241 = TR_36 ;
	7'h6c :
		TR_241 = TR_36 ;
	7'h6d :
		TR_241 = TR_36 ;
	7'h6e :
		TR_241 = TR_36 ;
	7'h6f :
		TR_241 = TR_36 ;
	7'h70 :
		TR_241 = TR_36 ;
	7'h71 :
		TR_241 = TR_36 ;
	7'h72 :
		TR_241 = TR_36 ;
	7'h73 :
		TR_241 = TR_36 ;
	7'h74 :
		TR_241 = TR_36 ;
	7'h75 :
		TR_241 = TR_36 ;
	7'h76 :
		TR_241 = TR_36 ;
	7'h77 :
		TR_241 = TR_36 ;
	7'h78 :
		TR_241 = TR_36 ;
	7'h79 :
		TR_241 = TR_36 ;
	7'h7a :
		TR_241 = TR_36 ;
	7'h7b :
		TR_241 = TR_36 ;
	7'h7c :
		TR_241 = TR_36 ;
	7'h7d :
		TR_241 = TR_36 ;
	7'h7e :
		TR_241 = TR_36 ;
	7'h7f :
		TR_241 = TR_36 ;
	default :
		TR_241 = 9'hx ;
	endcase
always @ ( TR_241 or U_173 or sub8u_71ot or U_183 or RG_rl_141 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_24_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h18 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_24_t = ( ( { 9{ M_180 } } & RG_rl_141 )
		| ( { 9{ U_173 } } & TR_241 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_24_en = ( M_180 | RG_rl_24_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_24_en )
		RG_rl_24 <= RG_rl_24_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_37 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_240 = TR_37 ;
	7'h01 :
		TR_240 = TR_37 ;
	7'h02 :
		TR_240 = TR_37 ;
	7'h03 :
		TR_240 = TR_37 ;
	7'h04 :
		TR_240 = TR_37 ;
	7'h05 :
		TR_240 = TR_37 ;
	7'h06 :
		TR_240 = TR_37 ;
	7'h07 :
		TR_240 = TR_37 ;
	7'h08 :
		TR_240 = TR_37 ;
	7'h09 :
		TR_240 = TR_37 ;
	7'h0a :
		TR_240 = TR_37 ;
	7'h0b :
		TR_240 = TR_37 ;
	7'h0c :
		TR_240 = TR_37 ;
	7'h0d :
		TR_240 = TR_37 ;
	7'h0e :
		TR_240 = TR_37 ;
	7'h0f :
		TR_240 = TR_37 ;
	7'h10 :
		TR_240 = TR_37 ;
	7'h11 :
		TR_240 = TR_37 ;
	7'h12 :
		TR_240 = TR_37 ;
	7'h13 :
		TR_240 = TR_37 ;
	7'h14 :
		TR_240 = TR_37 ;
	7'h15 :
		TR_240 = TR_37 ;
	7'h16 :
		TR_240 = TR_37 ;
	7'h17 :
		TR_240 = TR_37 ;
	7'h18 :
		TR_240 = TR_37 ;
	7'h19 :
		TR_240 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1a :
		TR_240 = TR_37 ;
	7'h1b :
		TR_240 = TR_37 ;
	7'h1c :
		TR_240 = TR_37 ;
	7'h1d :
		TR_240 = TR_37 ;
	7'h1e :
		TR_240 = TR_37 ;
	7'h1f :
		TR_240 = TR_37 ;
	7'h20 :
		TR_240 = TR_37 ;
	7'h21 :
		TR_240 = TR_37 ;
	7'h22 :
		TR_240 = TR_37 ;
	7'h23 :
		TR_240 = TR_37 ;
	7'h24 :
		TR_240 = TR_37 ;
	7'h25 :
		TR_240 = TR_37 ;
	7'h26 :
		TR_240 = TR_37 ;
	7'h27 :
		TR_240 = TR_37 ;
	7'h28 :
		TR_240 = TR_37 ;
	7'h29 :
		TR_240 = TR_37 ;
	7'h2a :
		TR_240 = TR_37 ;
	7'h2b :
		TR_240 = TR_37 ;
	7'h2c :
		TR_240 = TR_37 ;
	7'h2d :
		TR_240 = TR_37 ;
	7'h2e :
		TR_240 = TR_37 ;
	7'h2f :
		TR_240 = TR_37 ;
	7'h30 :
		TR_240 = TR_37 ;
	7'h31 :
		TR_240 = TR_37 ;
	7'h32 :
		TR_240 = TR_37 ;
	7'h33 :
		TR_240 = TR_37 ;
	7'h34 :
		TR_240 = TR_37 ;
	7'h35 :
		TR_240 = TR_37 ;
	7'h36 :
		TR_240 = TR_37 ;
	7'h37 :
		TR_240 = TR_37 ;
	7'h38 :
		TR_240 = TR_37 ;
	7'h39 :
		TR_240 = TR_37 ;
	7'h3a :
		TR_240 = TR_37 ;
	7'h3b :
		TR_240 = TR_37 ;
	7'h3c :
		TR_240 = TR_37 ;
	7'h3d :
		TR_240 = TR_37 ;
	7'h3e :
		TR_240 = TR_37 ;
	7'h3f :
		TR_240 = TR_37 ;
	7'h40 :
		TR_240 = TR_37 ;
	7'h41 :
		TR_240 = TR_37 ;
	7'h42 :
		TR_240 = TR_37 ;
	7'h43 :
		TR_240 = TR_37 ;
	7'h44 :
		TR_240 = TR_37 ;
	7'h45 :
		TR_240 = TR_37 ;
	7'h46 :
		TR_240 = TR_37 ;
	7'h47 :
		TR_240 = TR_37 ;
	7'h48 :
		TR_240 = TR_37 ;
	7'h49 :
		TR_240 = TR_37 ;
	7'h4a :
		TR_240 = TR_37 ;
	7'h4b :
		TR_240 = TR_37 ;
	7'h4c :
		TR_240 = TR_37 ;
	7'h4d :
		TR_240 = TR_37 ;
	7'h4e :
		TR_240 = TR_37 ;
	7'h4f :
		TR_240 = TR_37 ;
	7'h50 :
		TR_240 = TR_37 ;
	7'h51 :
		TR_240 = TR_37 ;
	7'h52 :
		TR_240 = TR_37 ;
	7'h53 :
		TR_240 = TR_37 ;
	7'h54 :
		TR_240 = TR_37 ;
	7'h55 :
		TR_240 = TR_37 ;
	7'h56 :
		TR_240 = TR_37 ;
	7'h57 :
		TR_240 = TR_37 ;
	7'h58 :
		TR_240 = TR_37 ;
	7'h59 :
		TR_240 = TR_37 ;
	7'h5a :
		TR_240 = TR_37 ;
	7'h5b :
		TR_240 = TR_37 ;
	7'h5c :
		TR_240 = TR_37 ;
	7'h5d :
		TR_240 = TR_37 ;
	7'h5e :
		TR_240 = TR_37 ;
	7'h5f :
		TR_240 = TR_37 ;
	7'h60 :
		TR_240 = TR_37 ;
	7'h61 :
		TR_240 = TR_37 ;
	7'h62 :
		TR_240 = TR_37 ;
	7'h63 :
		TR_240 = TR_37 ;
	7'h64 :
		TR_240 = TR_37 ;
	7'h65 :
		TR_240 = TR_37 ;
	7'h66 :
		TR_240 = TR_37 ;
	7'h67 :
		TR_240 = TR_37 ;
	7'h68 :
		TR_240 = TR_37 ;
	7'h69 :
		TR_240 = TR_37 ;
	7'h6a :
		TR_240 = TR_37 ;
	7'h6b :
		TR_240 = TR_37 ;
	7'h6c :
		TR_240 = TR_37 ;
	7'h6d :
		TR_240 = TR_37 ;
	7'h6e :
		TR_240 = TR_37 ;
	7'h6f :
		TR_240 = TR_37 ;
	7'h70 :
		TR_240 = TR_37 ;
	7'h71 :
		TR_240 = TR_37 ;
	7'h72 :
		TR_240 = TR_37 ;
	7'h73 :
		TR_240 = TR_37 ;
	7'h74 :
		TR_240 = TR_37 ;
	7'h75 :
		TR_240 = TR_37 ;
	7'h76 :
		TR_240 = TR_37 ;
	7'h77 :
		TR_240 = TR_37 ;
	7'h78 :
		TR_240 = TR_37 ;
	7'h79 :
		TR_240 = TR_37 ;
	7'h7a :
		TR_240 = TR_37 ;
	7'h7b :
		TR_240 = TR_37 ;
	7'h7c :
		TR_240 = TR_37 ;
	7'h7d :
		TR_240 = TR_37 ;
	7'h7e :
		TR_240 = TR_37 ;
	7'h7f :
		TR_240 = TR_37 ;
	default :
		TR_240 = 9'hx ;
	endcase
always @ ( TR_240 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_10 or 
	U_174 or RG_rl_141 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_25_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h19 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_25_t = ( ( { 9{ ST1_03d } } & RG_rl_141 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_10 )
		| ( { 9{ U_173 } } & TR_240 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_25_en = ( ST1_03d | U_174 | RG_rl_25_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_25_en )
		RG_rl_25 <= RG_rl_25_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_38 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_239 = TR_38 ;
	7'h01 :
		TR_239 = TR_38 ;
	7'h02 :
		TR_239 = TR_38 ;
	7'h03 :
		TR_239 = TR_38 ;
	7'h04 :
		TR_239 = TR_38 ;
	7'h05 :
		TR_239 = TR_38 ;
	7'h06 :
		TR_239 = TR_38 ;
	7'h07 :
		TR_239 = TR_38 ;
	7'h08 :
		TR_239 = TR_38 ;
	7'h09 :
		TR_239 = TR_38 ;
	7'h0a :
		TR_239 = TR_38 ;
	7'h0b :
		TR_239 = TR_38 ;
	7'h0c :
		TR_239 = TR_38 ;
	7'h0d :
		TR_239 = TR_38 ;
	7'h0e :
		TR_239 = TR_38 ;
	7'h0f :
		TR_239 = TR_38 ;
	7'h10 :
		TR_239 = TR_38 ;
	7'h11 :
		TR_239 = TR_38 ;
	7'h12 :
		TR_239 = TR_38 ;
	7'h13 :
		TR_239 = TR_38 ;
	7'h14 :
		TR_239 = TR_38 ;
	7'h15 :
		TR_239 = TR_38 ;
	7'h16 :
		TR_239 = TR_38 ;
	7'h17 :
		TR_239 = TR_38 ;
	7'h18 :
		TR_239 = TR_38 ;
	7'h19 :
		TR_239 = TR_38 ;
	7'h1a :
		TR_239 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1b :
		TR_239 = TR_38 ;
	7'h1c :
		TR_239 = TR_38 ;
	7'h1d :
		TR_239 = TR_38 ;
	7'h1e :
		TR_239 = TR_38 ;
	7'h1f :
		TR_239 = TR_38 ;
	7'h20 :
		TR_239 = TR_38 ;
	7'h21 :
		TR_239 = TR_38 ;
	7'h22 :
		TR_239 = TR_38 ;
	7'h23 :
		TR_239 = TR_38 ;
	7'h24 :
		TR_239 = TR_38 ;
	7'h25 :
		TR_239 = TR_38 ;
	7'h26 :
		TR_239 = TR_38 ;
	7'h27 :
		TR_239 = TR_38 ;
	7'h28 :
		TR_239 = TR_38 ;
	7'h29 :
		TR_239 = TR_38 ;
	7'h2a :
		TR_239 = TR_38 ;
	7'h2b :
		TR_239 = TR_38 ;
	7'h2c :
		TR_239 = TR_38 ;
	7'h2d :
		TR_239 = TR_38 ;
	7'h2e :
		TR_239 = TR_38 ;
	7'h2f :
		TR_239 = TR_38 ;
	7'h30 :
		TR_239 = TR_38 ;
	7'h31 :
		TR_239 = TR_38 ;
	7'h32 :
		TR_239 = TR_38 ;
	7'h33 :
		TR_239 = TR_38 ;
	7'h34 :
		TR_239 = TR_38 ;
	7'h35 :
		TR_239 = TR_38 ;
	7'h36 :
		TR_239 = TR_38 ;
	7'h37 :
		TR_239 = TR_38 ;
	7'h38 :
		TR_239 = TR_38 ;
	7'h39 :
		TR_239 = TR_38 ;
	7'h3a :
		TR_239 = TR_38 ;
	7'h3b :
		TR_239 = TR_38 ;
	7'h3c :
		TR_239 = TR_38 ;
	7'h3d :
		TR_239 = TR_38 ;
	7'h3e :
		TR_239 = TR_38 ;
	7'h3f :
		TR_239 = TR_38 ;
	7'h40 :
		TR_239 = TR_38 ;
	7'h41 :
		TR_239 = TR_38 ;
	7'h42 :
		TR_239 = TR_38 ;
	7'h43 :
		TR_239 = TR_38 ;
	7'h44 :
		TR_239 = TR_38 ;
	7'h45 :
		TR_239 = TR_38 ;
	7'h46 :
		TR_239 = TR_38 ;
	7'h47 :
		TR_239 = TR_38 ;
	7'h48 :
		TR_239 = TR_38 ;
	7'h49 :
		TR_239 = TR_38 ;
	7'h4a :
		TR_239 = TR_38 ;
	7'h4b :
		TR_239 = TR_38 ;
	7'h4c :
		TR_239 = TR_38 ;
	7'h4d :
		TR_239 = TR_38 ;
	7'h4e :
		TR_239 = TR_38 ;
	7'h4f :
		TR_239 = TR_38 ;
	7'h50 :
		TR_239 = TR_38 ;
	7'h51 :
		TR_239 = TR_38 ;
	7'h52 :
		TR_239 = TR_38 ;
	7'h53 :
		TR_239 = TR_38 ;
	7'h54 :
		TR_239 = TR_38 ;
	7'h55 :
		TR_239 = TR_38 ;
	7'h56 :
		TR_239 = TR_38 ;
	7'h57 :
		TR_239 = TR_38 ;
	7'h58 :
		TR_239 = TR_38 ;
	7'h59 :
		TR_239 = TR_38 ;
	7'h5a :
		TR_239 = TR_38 ;
	7'h5b :
		TR_239 = TR_38 ;
	7'h5c :
		TR_239 = TR_38 ;
	7'h5d :
		TR_239 = TR_38 ;
	7'h5e :
		TR_239 = TR_38 ;
	7'h5f :
		TR_239 = TR_38 ;
	7'h60 :
		TR_239 = TR_38 ;
	7'h61 :
		TR_239 = TR_38 ;
	7'h62 :
		TR_239 = TR_38 ;
	7'h63 :
		TR_239 = TR_38 ;
	7'h64 :
		TR_239 = TR_38 ;
	7'h65 :
		TR_239 = TR_38 ;
	7'h66 :
		TR_239 = TR_38 ;
	7'h67 :
		TR_239 = TR_38 ;
	7'h68 :
		TR_239 = TR_38 ;
	7'h69 :
		TR_239 = TR_38 ;
	7'h6a :
		TR_239 = TR_38 ;
	7'h6b :
		TR_239 = TR_38 ;
	7'h6c :
		TR_239 = TR_38 ;
	7'h6d :
		TR_239 = TR_38 ;
	7'h6e :
		TR_239 = TR_38 ;
	7'h6f :
		TR_239 = TR_38 ;
	7'h70 :
		TR_239 = TR_38 ;
	7'h71 :
		TR_239 = TR_38 ;
	7'h72 :
		TR_239 = TR_38 ;
	7'h73 :
		TR_239 = TR_38 ;
	7'h74 :
		TR_239 = TR_38 ;
	7'h75 :
		TR_239 = TR_38 ;
	7'h76 :
		TR_239 = TR_38 ;
	7'h77 :
		TR_239 = TR_38 ;
	7'h78 :
		TR_239 = TR_38 ;
	7'h79 :
		TR_239 = TR_38 ;
	7'h7a :
		TR_239 = TR_38 ;
	7'h7b :
		TR_239 = TR_38 ;
	7'h7c :
		TR_239 = TR_38 ;
	7'h7d :
		TR_239 = TR_38 ;
	7'h7e :
		TR_239 = TR_38 ;
	7'h7f :
		TR_239 = TR_38 ;
	default :
		TR_239 = 9'hx ;
	endcase
always @ ( TR_239 or U_173 or sub8u_71ot or U_183 or RG_rl_142 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_26_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h1a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_26_t = ( ( { 9{ M_180 } } & RG_rl_142 )
		| ( { 9{ U_173 } } & TR_239 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_26_en = ( M_180 | RG_rl_26_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_26_en )
		RG_rl_26 <= RG_rl_26_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_39 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_238 = TR_39 ;
	7'h01 :
		TR_238 = TR_39 ;
	7'h02 :
		TR_238 = TR_39 ;
	7'h03 :
		TR_238 = TR_39 ;
	7'h04 :
		TR_238 = TR_39 ;
	7'h05 :
		TR_238 = TR_39 ;
	7'h06 :
		TR_238 = TR_39 ;
	7'h07 :
		TR_238 = TR_39 ;
	7'h08 :
		TR_238 = TR_39 ;
	7'h09 :
		TR_238 = TR_39 ;
	7'h0a :
		TR_238 = TR_39 ;
	7'h0b :
		TR_238 = TR_39 ;
	7'h0c :
		TR_238 = TR_39 ;
	7'h0d :
		TR_238 = TR_39 ;
	7'h0e :
		TR_238 = TR_39 ;
	7'h0f :
		TR_238 = TR_39 ;
	7'h10 :
		TR_238 = TR_39 ;
	7'h11 :
		TR_238 = TR_39 ;
	7'h12 :
		TR_238 = TR_39 ;
	7'h13 :
		TR_238 = TR_39 ;
	7'h14 :
		TR_238 = TR_39 ;
	7'h15 :
		TR_238 = TR_39 ;
	7'h16 :
		TR_238 = TR_39 ;
	7'h17 :
		TR_238 = TR_39 ;
	7'h18 :
		TR_238 = TR_39 ;
	7'h19 :
		TR_238 = TR_39 ;
	7'h1a :
		TR_238 = TR_39 ;
	7'h1b :
		TR_238 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1c :
		TR_238 = TR_39 ;
	7'h1d :
		TR_238 = TR_39 ;
	7'h1e :
		TR_238 = TR_39 ;
	7'h1f :
		TR_238 = TR_39 ;
	7'h20 :
		TR_238 = TR_39 ;
	7'h21 :
		TR_238 = TR_39 ;
	7'h22 :
		TR_238 = TR_39 ;
	7'h23 :
		TR_238 = TR_39 ;
	7'h24 :
		TR_238 = TR_39 ;
	7'h25 :
		TR_238 = TR_39 ;
	7'h26 :
		TR_238 = TR_39 ;
	7'h27 :
		TR_238 = TR_39 ;
	7'h28 :
		TR_238 = TR_39 ;
	7'h29 :
		TR_238 = TR_39 ;
	7'h2a :
		TR_238 = TR_39 ;
	7'h2b :
		TR_238 = TR_39 ;
	7'h2c :
		TR_238 = TR_39 ;
	7'h2d :
		TR_238 = TR_39 ;
	7'h2e :
		TR_238 = TR_39 ;
	7'h2f :
		TR_238 = TR_39 ;
	7'h30 :
		TR_238 = TR_39 ;
	7'h31 :
		TR_238 = TR_39 ;
	7'h32 :
		TR_238 = TR_39 ;
	7'h33 :
		TR_238 = TR_39 ;
	7'h34 :
		TR_238 = TR_39 ;
	7'h35 :
		TR_238 = TR_39 ;
	7'h36 :
		TR_238 = TR_39 ;
	7'h37 :
		TR_238 = TR_39 ;
	7'h38 :
		TR_238 = TR_39 ;
	7'h39 :
		TR_238 = TR_39 ;
	7'h3a :
		TR_238 = TR_39 ;
	7'h3b :
		TR_238 = TR_39 ;
	7'h3c :
		TR_238 = TR_39 ;
	7'h3d :
		TR_238 = TR_39 ;
	7'h3e :
		TR_238 = TR_39 ;
	7'h3f :
		TR_238 = TR_39 ;
	7'h40 :
		TR_238 = TR_39 ;
	7'h41 :
		TR_238 = TR_39 ;
	7'h42 :
		TR_238 = TR_39 ;
	7'h43 :
		TR_238 = TR_39 ;
	7'h44 :
		TR_238 = TR_39 ;
	7'h45 :
		TR_238 = TR_39 ;
	7'h46 :
		TR_238 = TR_39 ;
	7'h47 :
		TR_238 = TR_39 ;
	7'h48 :
		TR_238 = TR_39 ;
	7'h49 :
		TR_238 = TR_39 ;
	7'h4a :
		TR_238 = TR_39 ;
	7'h4b :
		TR_238 = TR_39 ;
	7'h4c :
		TR_238 = TR_39 ;
	7'h4d :
		TR_238 = TR_39 ;
	7'h4e :
		TR_238 = TR_39 ;
	7'h4f :
		TR_238 = TR_39 ;
	7'h50 :
		TR_238 = TR_39 ;
	7'h51 :
		TR_238 = TR_39 ;
	7'h52 :
		TR_238 = TR_39 ;
	7'h53 :
		TR_238 = TR_39 ;
	7'h54 :
		TR_238 = TR_39 ;
	7'h55 :
		TR_238 = TR_39 ;
	7'h56 :
		TR_238 = TR_39 ;
	7'h57 :
		TR_238 = TR_39 ;
	7'h58 :
		TR_238 = TR_39 ;
	7'h59 :
		TR_238 = TR_39 ;
	7'h5a :
		TR_238 = TR_39 ;
	7'h5b :
		TR_238 = TR_39 ;
	7'h5c :
		TR_238 = TR_39 ;
	7'h5d :
		TR_238 = TR_39 ;
	7'h5e :
		TR_238 = TR_39 ;
	7'h5f :
		TR_238 = TR_39 ;
	7'h60 :
		TR_238 = TR_39 ;
	7'h61 :
		TR_238 = TR_39 ;
	7'h62 :
		TR_238 = TR_39 ;
	7'h63 :
		TR_238 = TR_39 ;
	7'h64 :
		TR_238 = TR_39 ;
	7'h65 :
		TR_238 = TR_39 ;
	7'h66 :
		TR_238 = TR_39 ;
	7'h67 :
		TR_238 = TR_39 ;
	7'h68 :
		TR_238 = TR_39 ;
	7'h69 :
		TR_238 = TR_39 ;
	7'h6a :
		TR_238 = TR_39 ;
	7'h6b :
		TR_238 = TR_39 ;
	7'h6c :
		TR_238 = TR_39 ;
	7'h6d :
		TR_238 = TR_39 ;
	7'h6e :
		TR_238 = TR_39 ;
	7'h6f :
		TR_238 = TR_39 ;
	7'h70 :
		TR_238 = TR_39 ;
	7'h71 :
		TR_238 = TR_39 ;
	7'h72 :
		TR_238 = TR_39 ;
	7'h73 :
		TR_238 = TR_39 ;
	7'h74 :
		TR_238 = TR_39 ;
	7'h75 :
		TR_238 = TR_39 ;
	7'h76 :
		TR_238 = TR_39 ;
	7'h77 :
		TR_238 = TR_39 ;
	7'h78 :
		TR_238 = TR_39 ;
	7'h79 :
		TR_238 = TR_39 ;
	7'h7a :
		TR_238 = TR_39 ;
	7'h7b :
		TR_238 = TR_39 ;
	7'h7c :
		TR_238 = TR_39 ;
	7'h7d :
		TR_238 = TR_39 ;
	7'h7e :
		TR_238 = TR_39 ;
	7'h7f :
		TR_238 = TR_39 ;
	default :
		TR_238 = 9'hx ;
	endcase
always @ ( TR_238 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_11 or 
	U_174 or RG_rl_142 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_27_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h1b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_27_t = ( ( { 9{ ST1_03d } } & RG_rl_142 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_11 )
		| ( { 9{ U_173 } } & TR_238 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_27_en = ( ST1_03d | U_174 | RG_rl_27_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_27_en )
		RG_rl_27 <= RG_rl_27_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_40 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_237 = TR_40 ;
	7'h01 :
		TR_237 = TR_40 ;
	7'h02 :
		TR_237 = TR_40 ;
	7'h03 :
		TR_237 = TR_40 ;
	7'h04 :
		TR_237 = TR_40 ;
	7'h05 :
		TR_237 = TR_40 ;
	7'h06 :
		TR_237 = TR_40 ;
	7'h07 :
		TR_237 = TR_40 ;
	7'h08 :
		TR_237 = TR_40 ;
	7'h09 :
		TR_237 = TR_40 ;
	7'h0a :
		TR_237 = TR_40 ;
	7'h0b :
		TR_237 = TR_40 ;
	7'h0c :
		TR_237 = TR_40 ;
	7'h0d :
		TR_237 = TR_40 ;
	7'h0e :
		TR_237 = TR_40 ;
	7'h0f :
		TR_237 = TR_40 ;
	7'h10 :
		TR_237 = TR_40 ;
	7'h11 :
		TR_237 = TR_40 ;
	7'h12 :
		TR_237 = TR_40 ;
	7'h13 :
		TR_237 = TR_40 ;
	7'h14 :
		TR_237 = TR_40 ;
	7'h15 :
		TR_237 = TR_40 ;
	7'h16 :
		TR_237 = TR_40 ;
	7'h17 :
		TR_237 = TR_40 ;
	7'h18 :
		TR_237 = TR_40 ;
	7'h19 :
		TR_237 = TR_40 ;
	7'h1a :
		TR_237 = TR_40 ;
	7'h1b :
		TR_237 = TR_40 ;
	7'h1c :
		TR_237 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1d :
		TR_237 = TR_40 ;
	7'h1e :
		TR_237 = TR_40 ;
	7'h1f :
		TR_237 = TR_40 ;
	7'h20 :
		TR_237 = TR_40 ;
	7'h21 :
		TR_237 = TR_40 ;
	7'h22 :
		TR_237 = TR_40 ;
	7'h23 :
		TR_237 = TR_40 ;
	7'h24 :
		TR_237 = TR_40 ;
	7'h25 :
		TR_237 = TR_40 ;
	7'h26 :
		TR_237 = TR_40 ;
	7'h27 :
		TR_237 = TR_40 ;
	7'h28 :
		TR_237 = TR_40 ;
	7'h29 :
		TR_237 = TR_40 ;
	7'h2a :
		TR_237 = TR_40 ;
	7'h2b :
		TR_237 = TR_40 ;
	7'h2c :
		TR_237 = TR_40 ;
	7'h2d :
		TR_237 = TR_40 ;
	7'h2e :
		TR_237 = TR_40 ;
	7'h2f :
		TR_237 = TR_40 ;
	7'h30 :
		TR_237 = TR_40 ;
	7'h31 :
		TR_237 = TR_40 ;
	7'h32 :
		TR_237 = TR_40 ;
	7'h33 :
		TR_237 = TR_40 ;
	7'h34 :
		TR_237 = TR_40 ;
	7'h35 :
		TR_237 = TR_40 ;
	7'h36 :
		TR_237 = TR_40 ;
	7'h37 :
		TR_237 = TR_40 ;
	7'h38 :
		TR_237 = TR_40 ;
	7'h39 :
		TR_237 = TR_40 ;
	7'h3a :
		TR_237 = TR_40 ;
	7'h3b :
		TR_237 = TR_40 ;
	7'h3c :
		TR_237 = TR_40 ;
	7'h3d :
		TR_237 = TR_40 ;
	7'h3e :
		TR_237 = TR_40 ;
	7'h3f :
		TR_237 = TR_40 ;
	7'h40 :
		TR_237 = TR_40 ;
	7'h41 :
		TR_237 = TR_40 ;
	7'h42 :
		TR_237 = TR_40 ;
	7'h43 :
		TR_237 = TR_40 ;
	7'h44 :
		TR_237 = TR_40 ;
	7'h45 :
		TR_237 = TR_40 ;
	7'h46 :
		TR_237 = TR_40 ;
	7'h47 :
		TR_237 = TR_40 ;
	7'h48 :
		TR_237 = TR_40 ;
	7'h49 :
		TR_237 = TR_40 ;
	7'h4a :
		TR_237 = TR_40 ;
	7'h4b :
		TR_237 = TR_40 ;
	7'h4c :
		TR_237 = TR_40 ;
	7'h4d :
		TR_237 = TR_40 ;
	7'h4e :
		TR_237 = TR_40 ;
	7'h4f :
		TR_237 = TR_40 ;
	7'h50 :
		TR_237 = TR_40 ;
	7'h51 :
		TR_237 = TR_40 ;
	7'h52 :
		TR_237 = TR_40 ;
	7'h53 :
		TR_237 = TR_40 ;
	7'h54 :
		TR_237 = TR_40 ;
	7'h55 :
		TR_237 = TR_40 ;
	7'h56 :
		TR_237 = TR_40 ;
	7'h57 :
		TR_237 = TR_40 ;
	7'h58 :
		TR_237 = TR_40 ;
	7'h59 :
		TR_237 = TR_40 ;
	7'h5a :
		TR_237 = TR_40 ;
	7'h5b :
		TR_237 = TR_40 ;
	7'h5c :
		TR_237 = TR_40 ;
	7'h5d :
		TR_237 = TR_40 ;
	7'h5e :
		TR_237 = TR_40 ;
	7'h5f :
		TR_237 = TR_40 ;
	7'h60 :
		TR_237 = TR_40 ;
	7'h61 :
		TR_237 = TR_40 ;
	7'h62 :
		TR_237 = TR_40 ;
	7'h63 :
		TR_237 = TR_40 ;
	7'h64 :
		TR_237 = TR_40 ;
	7'h65 :
		TR_237 = TR_40 ;
	7'h66 :
		TR_237 = TR_40 ;
	7'h67 :
		TR_237 = TR_40 ;
	7'h68 :
		TR_237 = TR_40 ;
	7'h69 :
		TR_237 = TR_40 ;
	7'h6a :
		TR_237 = TR_40 ;
	7'h6b :
		TR_237 = TR_40 ;
	7'h6c :
		TR_237 = TR_40 ;
	7'h6d :
		TR_237 = TR_40 ;
	7'h6e :
		TR_237 = TR_40 ;
	7'h6f :
		TR_237 = TR_40 ;
	7'h70 :
		TR_237 = TR_40 ;
	7'h71 :
		TR_237 = TR_40 ;
	7'h72 :
		TR_237 = TR_40 ;
	7'h73 :
		TR_237 = TR_40 ;
	7'h74 :
		TR_237 = TR_40 ;
	7'h75 :
		TR_237 = TR_40 ;
	7'h76 :
		TR_237 = TR_40 ;
	7'h77 :
		TR_237 = TR_40 ;
	7'h78 :
		TR_237 = TR_40 ;
	7'h79 :
		TR_237 = TR_40 ;
	7'h7a :
		TR_237 = TR_40 ;
	7'h7b :
		TR_237 = TR_40 ;
	7'h7c :
		TR_237 = TR_40 ;
	7'h7d :
		TR_237 = TR_40 ;
	7'h7e :
		TR_237 = TR_40 ;
	7'h7f :
		TR_237 = TR_40 ;
	default :
		TR_237 = 9'hx ;
	endcase
always @ ( TR_237 or U_173 or sub8u_71ot or U_183 or RG_rl_143 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_28_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h1c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_28_t = ( ( { 9{ M_180 } } & RG_rl_143 )
		| ( { 9{ U_173 } } & TR_237 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_28_en = ( M_180 | RG_rl_28_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_28_en )
		RG_rl_28 <= RG_rl_28_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_41 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_236 = TR_41 ;
	7'h01 :
		TR_236 = TR_41 ;
	7'h02 :
		TR_236 = TR_41 ;
	7'h03 :
		TR_236 = TR_41 ;
	7'h04 :
		TR_236 = TR_41 ;
	7'h05 :
		TR_236 = TR_41 ;
	7'h06 :
		TR_236 = TR_41 ;
	7'h07 :
		TR_236 = TR_41 ;
	7'h08 :
		TR_236 = TR_41 ;
	7'h09 :
		TR_236 = TR_41 ;
	7'h0a :
		TR_236 = TR_41 ;
	7'h0b :
		TR_236 = TR_41 ;
	7'h0c :
		TR_236 = TR_41 ;
	7'h0d :
		TR_236 = TR_41 ;
	7'h0e :
		TR_236 = TR_41 ;
	7'h0f :
		TR_236 = TR_41 ;
	7'h10 :
		TR_236 = TR_41 ;
	7'h11 :
		TR_236 = TR_41 ;
	7'h12 :
		TR_236 = TR_41 ;
	7'h13 :
		TR_236 = TR_41 ;
	7'h14 :
		TR_236 = TR_41 ;
	7'h15 :
		TR_236 = TR_41 ;
	7'h16 :
		TR_236 = TR_41 ;
	7'h17 :
		TR_236 = TR_41 ;
	7'h18 :
		TR_236 = TR_41 ;
	7'h19 :
		TR_236 = TR_41 ;
	7'h1a :
		TR_236 = TR_41 ;
	7'h1b :
		TR_236 = TR_41 ;
	7'h1c :
		TR_236 = TR_41 ;
	7'h1d :
		TR_236 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1e :
		TR_236 = TR_41 ;
	7'h1f :
		TR_236 = TR_41 ;
	7'h20 :
		TR_236 = TR_41 ;
	7'h21 :
		TR_236 = TR_41 ;
	7'h22 :
		TR_236 = TR_41 ;
	7'h23 :
		TR_236 = TR_41 ;
	7'h24 :
		TR_236 = TR_41 ;
	7'h25 :
		TR_236 = TR_41 ;
	7'h26 :
		TR_236 = TR_41 ;
	7'h27 :
		TR_236 = TR_41 ;
	7'h28 :
		TR_236 = TR_41 ;
	7'h29 :
		TR_236 = TR_41 ;
	7'h2a :
		TR_236 = TR_41 ;
	7'h2b :
		TR_236 = TR_41 ;
	7'h2c :
		TR_236 = TR_41 ;
	7'h2d :
		TR_236 = TR_41 ;
	7'h2e :
		TR_236 = TR_41 ;
	7'h2f :
		TR_236 = TR_41 ;
	7'h30 :
		TR_236 = TR_41 ;
	7'h31 :
		TR_236 = TR_41 ;
	7'h32 :
		TR_236 = TR_41 ;
	7'h33 :
		TR_236 = TR_41 ;
	7'h34 :
		TR_236 = TR_41 ;
	7'h35 :
		TR_236 = TR_41 ;
	7'h36 :
		TR_236 = TR_41 ;
	7'h37 :
		TR_236 = TR_41 ;
	7'h38 :
		TR_236 = TR_41 ;
	7'h39 :
		TR_236 = TR_41 ;
	7'h3a :
		TR_236 = TR_41 ;
	7'h3b :
		TR_236 = TR_41 ;
	7'h3c :
		TR_236 = TR_41 ;
	7'h3d :
		TR_236 = TR_41 ;
	7'h3e :
		TR_236 = TR_41 ;
	7'h3f :
		TR_236 = TR_41 ;
	7'h40 :
		TR_236 = TR_41 ;
	7'h41 :
		TR_236 = TR_41 ;
	7'h42 :
		TR_236 = TR_41 ;
	7'h43 :
		TR_236 = TR_41 ;
	7'h44 :
		TR_236 = TR_41 ;
	7'h45 :
		TR_236 = TR_41 ;
	7'h46 :
		TR_236 = TR_41 ;
	7'h47 :
		TR_236 = TR_41 ;
	7'h48 :
		TR_236 = TR_41 ;
	7'h49 :
		TR_236 = TR_41 ;
	7'h4a :
		TR_236 = TR_41 ;
	7'h4b :
		TR_236 = TR_41 ;
	7'h4c :
		TR_236 = TR_41 ;
	7'h4d :
		TR_236 = TR_41 ;
	7'h4e :
		TR_236 = TR_41 ;
	7'h4f :
		TR_236 = TR_41 ;
	7'h50 :
		TR_236 = TR_41 ;
	7'h51 :
		TR_236 = TR_41 ;
	7'h52 :
		TR_236 = TR_41 ;
	7'h53 :
		TR_236 = TR_41 ;
	7'h54 :
		TR_236 = TR_41 ;
	7'h55 :
		TR_236 = TR_41 ;
	7'h56 :
		TR_236 = TR_41 ;
	7'h57 :
		TR_236 = TR_41 ;
	7'h58 :
		TR_236 = TR_41 ;
	7'h59 :
		TR_236 = TR_41 ;
	7'h5a :
		TR_236 = TR_41 ;
	7'h5b :
		TR_236 = TR_41 ;
	7'h5c :
		TR_236 = TR_41 ;
	7'h5d :
		TR_236 = TR_41 ;
	7'h5e :
		TR_236 = TR_41 ;
	7'h5f :
		TR_236 = TR_41 ;
	7'h60 :
		TR_236 = TR_41 ;
	7'h61 :
		TR_236 = TR_41 ;
	7'h62 :
		TR_236 = TR_41 ;
	7'h63 :
		TR_236 = TR_41 ;
	7'h64 :
		TR_236 = TR_41 ;
	7'h65 :
		TR_236 = TR_41 ;
	7'h66 :
		TR_236 = TR_41 ;
	7'h67 :
		TR_236 = TR_41 ;
	7'h68 :
		TR_236 = TR_41 ;
	7'h69 :
		TR_236 = TR_41 ;
	7'h6a :
		TR_236 = TR_41 ;
	7'h6b :
		TR_236 = TR_41 ;
	7'h6c :
		TR_236 = TR_41 ;
	7'h6d :
		TR_236 = TR_41 ;
	7'h6e :
		TR_236 = TR_41 ;
	7'h6f :
		TR_236 = TR_41 ;
	7'h70 :
		TR_236 = TR_41 ;
	7'h71 :
		TR_236 = TR_41 ;
	7'h72 :
		TR_236 = TR_41 ;
	7'h73 :
		TR_236 = TR_41 ;
	7'h74 :
		TR_236 = TR_41 ;
	7'h75 :
		TR_236 = TR_41 ;
	7'h76 :
		TR_236 = TR_41 ;
	7'h77 :
		TR_236 = TR_41 ;
	7'h78 :
		TR_236 = TR_41 ;
	7'h79 :
		TR_236 = TR_41 ;
	7'h7a :
		TR_236 = TR_41 ;
	7'h7b :
		TR_236 = TR_41 ;
	7'h7c :
		TR_236 = TR_41 ;
	7'h7d :
		TR_236 = TR_41 ;
	7'h7e :
		TR_236 = TR_41 ;
	7'h7f :
		TR_236 = TR_41 ;
	default :
		TR_236 = 9'hx ;
	endcase
always @ ( TR_236 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_12 or 
	U_174 or RG_rl_143 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_29_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h1d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_29_t = ( ( { 9{ ST1_03d } } & RG_rl_143 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_12 )
		| ( { 9{ U_173 } } & TR_236 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_29_en = ( ST1_03d | U_174 | RG_rl_29_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_29_en )
		RG_rl_29 <= RG_rl_29_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_42 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_235 = TR_42 ;
	7'h01 :
		TR_235 = TR_42 ;
	7'h02 :
		TR_235 = TR_42 ;
	7'h03 :
		TR_235 = TR_42 ;
	7'h04 :
		TR_235 = TR_42 ;
	7'h05 :
		TR_235 = TR_42 ;
	7'h06 :
		TR_235 = TR_42 ;
	7'h07 :
		TR_235 = TR_42 ;
	7'h08 :
		TR_235 = TR_42 ;
	7'h09 :
		TR_235 = TR_42 ;
	7'h0a :
		TR_235 = TR_42 ;
	7'h0b :
		TR_235 = TR_42 ;
	7'h0c :
		TR_235 = TR_42 ;
	7'h0d :
		TR_235 = TR_42 ;
	7'h0e :
		TR_235 = TR_42 ;
	7'h0f :
		TR_235 = TR_42 ;
	7'h10 :
		TR_235 = TR_42 ;
	7'h11 :
		TR_235 = TR_42 ;
	7'h12 :
		TR_235 = TR_42 ;
	7'h13 :
		TR_235 = TR_42 ;
	7'h14 :
		TR_235 = TR_42 ;
	7'h15 :
		TR_235 = TR_42 ;
	7'h16 :
		TR_235 = TR_42 ;
	7'h17 :
		TR_235 = TR_42 ;
	7'h18 :
		TR_235 = TR_42 ;
	7'h19 :
		TR_235 = TR_42 ;
	7'h1a :
		TR_235 = TR_42 ;
	7'h1b :
		TR_235 = TR_42 ;
	7'h1c :
		TR_235 = TR_42 ;
	7'h1d :
		TR_235 = TR_42 ;
	7'h1e :
		TR_235 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1f :
		TR_235 = TR_42 ;
	7'h20 :
		TR_235 = TR_42 ;
	7'h21 :
		TR_235 = TR_42 ;
	7'h22 :
		TR_235 = TR_42 ;
	7'h23 :
		TR_235 = TR_42 ;
	7'h24 :
		TR_235 = TR_42 ;
	7'h25 :
		TR_235 = TR_42 ;
	7'h26 :
		TR_235 = TR_42 ;
	7'h27 :
		TR_235 = TR_42 ;
	7'h28 :
		TR_235 = TR_42 ;
	7'h29 :
		TR_235 = TR_42 ;
	7'h2a :
		TR_235 = TR_42 ;
	7'h2b :
		TR_235 = TR_42 ;
	7'h2c :
		TR_235 = TR_42 ;
	7'h2d :
		TR_235 = TR_42 ;
	7'h2e :
		TR_235 = TR_42 ;
	7'h2f :
		TR_235 = TR_42 ;
	7'h30 :
		TR_235 = TR_42 ;
	7'h31 :
		TR_235 = TR_42 ;
	7'h32 :
		TR_235 = TR_42 ;
	7'h33 :
		TR_235 = TR_42 ;
	7'h34 :
		TR_235 = TR_42 ;
	7'h35 :
		TR_235 = TR_42 ;
	7'h36 :
		TR_235 = TR_42 ;
	7'h37 :
		TR_235 = TR_42 ;
	7'h38 :
		TR_235 = TR_42 ;
	7'h39 :
		TR_235 = TR_42 ;
	7'h3a :
		TR_235 = TR_42 ;
	7'h3b :
		TR_235 = TR_42 ;
	7'h3c :
		TR_235 = TR_42 ;
	7'h3d :
		TR_235 = TR_42 ;
	7'h3e :
		TR_235 = TR_42 ;
	7'h3f :
		TR_235 = TR_42 ;
	7'h40 :
		TR_235 = TR_42 ;
	7'h41 :
		TR_235 = TR_42 ;
	7'h42 :
		TR_235 = TR_42 ;
	7'h43 :
		TR_235 = TR_42 ;
	7'h44 :
		TR_235 = TR_42 ;
	7'h45 :
		TR_235 = TR_42 ;
	7'h46 :
		TR_235 = TR_42 ;
	7'h47 :
		TR_235 = TR_42 ;
	7'h48 :
		TR_235 = TR_42 ;
	7'h49 :
		TR_235 = TR_42 ;
	7'h4a :
		TR_235 = TR_42 ;
	7'h4b :
		TR_235 = TR_42 ;
	7'h4c :
		TR_235 = TR_42 ;
	7'h4d :
		TR_235 = TR_42 ;
	7'h4e :
		TR_235 = TR_42 ;
	7'h4f :
		TR_235 = TR_42 ;
	7'h50 :
		TR_235 = TR_42 ;
	7'h51 :
		TR_235 = TR_42 ;
	7'h52 :
		TR_235 = TR_42 ;
	7'h53 :
		TR_235 = TR_42 ;
	7'h54 :
		TR_235 = TR_42 ;
	7'h55 :
		TR_235 = TR_42 ;
	7'h56 :
		TR_235 = TR_42 ;
	7'h57 :
		TR_235 = TR_42 ;
	7'h58 :
		TR_235 = TR_42 ;
	7'h59 :
		TR_235 = TR_42 ;
	7'h5a :
		TR_235 = TR_42 ;
	7'h5b :
		TR_235 = TR_42 ;
	7'h5c :
		TR_235 = TR_42 ;
	7'h5d :
		TR_235 = TR_42 ;
	7'h5e :
		TR_235 = TR_42 ;
	7'h5f :
		TR_235 = TR_42 ;
	7'h60 :
		TR_235 = TR_42 ;
	7'h61 :
		TR_235 = TR_42 ;
	7'h62 :
		TR_235 = TR_42 ;
	7'h63 :
		TR_235 = TR_42 ;
	7'h64 :
		TR_235 = TR_42 ;
	7'h65 :
		TR_235 = TR_42 ;
	7'h66 :
		TR_235 = TR_42 ;
	7'h67 :
		TR_235 = TR_42 ;
	7'h68 :
		TR_235 = TR_42 ;
	7'h69 :
		TR_235 = TR_42 ;
	7'h6a :
		TR_235 = TR_42 ;
	7'h6b :
		TR_235 = TR_42 ;
	7'h6c :
		TR_235 = TR_42 ;
	7'h6d :
		TR_235 = TR_42 ;
	7'h6e :
		TR_235 = TR_42 ;
	7'h6f :
		TR_235 = TR_42 ;
	7'h70 :
		TR_235 = TR_42 ;
	7'h71 :
		TR_235 = TR_42 ;
	7'h72 :
		TR_235 = TR_42 ;
	7'h73 :
		TR_235 = TR_42 ;
	7'h74 :
		TR_235 = TR_42 ;
	7'h75 :
		TR_235 = TR_42 ;
	7'h76 :
		TR_235 = TR_42 ;
	7'h77 :
		TR_235 = TR_42 ;
	7'h78 :
		TR_235 = TR_42 ;
	7'h79 :
		TR_235 = TR_42 ;
	7'h7a :
		TR_235 = TR_42 ;
	7'h7b :
		TR_235 = TR_42 ;
	7'h7c :
		TR_235 = TR_42 ;
	7'h7d :
		TR_235 = TR_42 ;
	7'h7e :
		TR_235 = TR_42 ;
	7'h7f :
		TR_235 = TR_42 ;
	default :
		TR_235 = 9'hx ;
	endcase
always @ ( TR_235 or U_173 or sub8u_71ot or U_183 or RG_rl_144 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_30_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h1e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_30_t = ( ( { 9{ M_180 } } & RG_rl_144 )
		| ( { 9{ U_173 } } & TR_235 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_30_en = ( M_180 | RG_rl_30_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_30_en )
		RG_rl_30 <= RG_rl_30_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_43 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_234 = TR_43 ;
	7'h01 :
		TR_234 = TR_43 ;
	7'h02 :
		TR_234 = TR_43 ;
	7'h03 :
		TR_234 = TR_43 ;
	7'h04 :
		TR_234 = TR_43 ;
	7'h05 :
		TR_234 = TR_43 ;
	7'h06 :
		TR_234 = TR_43 ;
	7'h07 :
		TR_234 = TR_43 ;
	7'h08 :
		TR_234 = TR_43 ;
	7'h09 :
		TR_234 = TR_43 ;
	7'h0a :
		TR_234 = TR_43 ;
	7'h0b :
		TR_234 = TR_43 ;
	7'h0c :
		TR_234 = TR_43 ;
	7'h0d :
		TR_234 = TR_43 ;
	7'h0e :
		TR_234 = TR_43 ;
	7'h0f :
		TR_234 = TR_43 ;
	7'h10 :
		TR_234 = TR_43 ;
	7'h11 :
		TR_234 = TR_43 ;
	7'h12 :
		TR_234 = TR_43 ;
	7'h13 :
		TR_234 = TR_43 ;
	7'h14 :
		TR_234 = TR_43 ;
	7'h15 :
		TR_234 = TR_43 ;
	7'h16 :
		TR_234 = TR_43 ;
	7'h17 :
		TR_234 = TR_43 ;
	7'h18 :
		TR_234 = TR_43 ;
	7'h19 :
		TR_234 = TR_43 ;
	7'h1a :
		TR_234 = TR_43 ;
	7'h1b :
		TR_234 = TR_43 ;
	7'h1c :
		TR_234 = TR_43 ;
	7'h1d :
		TR_234 = TR_43 ;
	7'h1e :
		TR_234 = TR_43 ;
	7'h1f :
		TR_234 = 9'h000 ;	// line#=../rle.cpp:80
	7'h20 :
		TR_234 = TR_43 ;
	7'h21 :
		TR_234 = TR_43 ;
	7'h22 :
		TR_234 = TR_43 ;
	7'h23 :
		TR_234 = TR_43 ;
	7'h24 :
		TR_234 = TR_43 ;
	7'h25 :
		TR_234 = TR_43 ;
	7'h26 :
		TR_234 = TR_43 ;
	7'h27 :
		TR_234 = TR_43 ;
	7'h28 :
		TR_234 = TR_43 ;
	7'h29 :
		TR_234 = TR_43 ;
	7'h2a :
		TR_234 = TR_43 ;
	7'h2b :
		TR_234 = TR_43 ;
	7'h2c :
		TR_234 = TR_43 ;
	7'h2d :
		TR_234 = TR_43 ;
	7'h2e :
		TR_234 = TR_43 ;
	7'h2f :
		TR_234 = TR_43 ;
	7'h30 :
		TR_234 = TR_43 ;
	7'h31 :
		TR_234 = TR_43 ;
	7'h32 :
		TR_234 = TR_43 ;
	7'h33 :
		TR_234 = TR_43 ;
	7'h34 :
		TR_234 = TR_43 ;
	7'h35 :
		TR_234 = TR_43 ;
	7'h36 :
		TR_234 = TR_43 ;
	7'h37 :
		TR_234 = TR_43 ;
	7'h38 :
		TR_234 = TR_43 ;
	7'h39 :
		TR_234 = TR_43 ;
	7'h3a :
		TR_234 = TR_43 ;
	7'h3b :
		TR_234 = TR_43 ;
	7'h3c :
		TR_234 = TR_43 ;
	7'h3d :
		TR_234 = TR_43 ;
	7'h3e :
		TR_234 = TR_43 ;
	7'h3f :
		TR_234 = TR_43 ;
	7'h40 :
		TR_234 = TR_43 ;
	7'h41 :
		TR_234 = TR_43 ;
	7'h42 :
		TR_234 = TR_43 ;
	7'h43 :
		TR_234 = TR_43 ;
	7'h44 :
		TR_234 = TR_43 ;
	7'h45 :
		TR_234 = TR_43 ;
	7'h46 :
		TR_234 = TR_43 ;
	7'h47 :
		TR_234 = TR_43 ;
	7'h48 :
		TR_234 = TR_43 ;
	7'h49 :
		TR_234 = TR_43 ;
	7'h4a :
		TR_234 = TR_43 ;
	7'h4b :
		TR_234 = TR_43 ;
	7'h4c :
		TR_234 = TR_43 ;
	7'h4d :
		TR_234 = TR_43 ;
	7'h4e :
		TR_234 = TR_43 ;
	7'h4f :
		TR_234 = TR_43 ;
	7'h50 :
		TR_234 = TR_43 ;
	7'h51 :
		TR_234 = TR_43 ;
	7'h52 :
		TR_234 = TR_43 ;
	7'h53 :
		TR_234 = TR_43 ;
	7'h54 :
		TR_234 = TR_43 ;
	7'h55 :
		TR_234 = TR_43 ;
	7'h56 :
		TR_234 = TR_43 ;
	7'h57 :
		TR_234 = TR_43 ;
	7'h58 :
		TR_234 = TR_43 ;
	7'h59 :
		TR_234 = TR_43 ;
	7'h5a :
		TR_234 = TR_43 ;
	7'h5b :
		TR_234 = TR_43 ;
	7'h5c :
		TR_234 = TR_43 ;
	7'h5d :
		TR_234 = TR_43 ;
	7'h5e :
		TR_234 = TR_43 ;
	7'h5f :
		TR_234 = TR_43 ;
	7'h60 :
		TR_234 = TR_43 ;
	7'h61 :
		TR_234 = TR_43 ;
	7'h62 :
		TR_234 = TR_43 ;
	7'h63 :
		TR_234 = TR_43 ;
	7'h64 :
		TR_234 = TR_43 ;
	7'h65 :
		TR_234 = TR_43 ;
	7'h66 :
		TR_234 = TR_43 ;
	7'h67 :
		TR_234 = TR_43 ;
	7'h68 :
		TR_234 = TR_43 ;
	7'h69 :
		TR_234 = TR_43 ;
	7'h6a :
		TR_234 = TR_43 ;
	7'h6b :
		TR_234 = TR_43 ;
	7'h6c :
		TR_234 = TR_43 ;
	7'h6d :
		TR_234 = TR_43 ;
	7'h6e :
		TR_234 = TR_43 ;
	7'h6f :
		TR_234 = TR_43 ;
	7'h70 :
		TR_234 = TR_43 ;
	7'h71 :
		TR_234 = TR_43 ;
	7'h72 :
		TR_234 = TR_43 ;
	7'h73 :
		TR_234 = TR_43 ;
	7'h74 :
		TR_234 = TR_43 ;
	7'h75 :
		TR_234 = TR_43 ;
	7'h76 :
		TR_234 = TR_43 ;
	7'h77 :
		TR_234 = TR_43 ;
	7'h78 :
		TR_234 = TR_43 ;
	7'h79 :
		TR_234 = TR_43 ;
	7'h7a :
		TR_234 = TR_43 ;
	7'h7b :
		TR_234 = TR_43 ;
	7'h7c :
		TR_234 = TR_43 ;
	7'h7d :
		TR_234 = TR_43 ;
	7'h7e :
		TR_234 = TR_43 ;
	7'h7f :
		TR_234 = TR_43 ;
	default :
		TR_234 = 9'hx ;
	endcase
always @ ( TR_234 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_13 or 
	U_174 or RG_rl_144 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_31_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h1f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_31_t = ( ( { 9{ ST1_03d } } & RG_rl_144 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_13 )
		| ( { 9{ U_173 } } & TR_234 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_31_en = ( ST1_03d | U_174 | RG_rl_31_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_31_en )
		RG_rl_31 <= RG_rl_31_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_44 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_233 = TR_44 ;
	7'h01 :
		TR_233 = TR_44 ;
	7'h02 :
		TR_233 = TR_44 ;
	7'h03 :
		TR_233 = TR_44 ;
	7'h04 :
		TR_233 = TR_44 ;
	7'h05 :
		TR_233 = TR_44 ;
	7'h06 :
		TR_233 = TR_44 ;
	7'h07 :
		TR_233 = TR_44 ;
	7'h08 :
		TR_233 = TR_44 ;
	7'h09 :
		TR_233 = TR_44 ;
	7'h0a :
		TR_233 = TR_44 ;
	7'h0b :
		TR_233 = TR_44 ;
	7'h0c :
		TR_233 = TR_44 ;
	7'h0d :
		TR_233 = TR_44 ;
	7'h0e :
		TR_233 = TR_44 ;
	7'h0f :
		TR_233 = TR_44 ;
	7'h10 :
		TR_233 = TR_44 ;
	7'h11 :
		TR_233 = TR_44 ;
	7'h12 :
		TR_233 = TR_44 ;
	7'h13 :
		TR_233 = TR_44 ;
	7'h14 :
		TR_233 = TR_44 ;
	7'h15 :
		TR_233 = TR_44 ;
	7'h16 :
		TR_233 = TR_44 ;
	7'h17 :
		TR_233 = TR_44 ;
	7'h18 :
		TR_233 = TR_44 ;
	7'h19 :
		TR_233 = TR_44 ;
	7'h1a :
		TR_233 = TR_44 ;
	7'h1b :
		TR_233 = TR_44 ;
	7'h1c :
		TR_233 = TR_44 ;
	7'h1d :
		TR_233 = TR_44 ;
	7'h1e :
		TR_233 = TR_44 ;
	7'h1f :
		TR_233 = TR_44 ;
	7'h20 :
		TR_233 = 9'h000 ;	// line#=../rle.cpp:80
	7'h21 :
		TR_233 = TR_44 ;
	7'h22 :
		TR_233 = TR_44 ;
	7'h23 :
		TR_233 = TR_44 ;
	7'h24 :
		TR_233 = TR_44 ;
	7'h25 :
		TR_233 = TR_44 ;
	7'h26 :
		TR_233 = TR_44 ;
	7'h27 :
		TR_233 = TR_44 ;
	7'h28 :
		TR_233 = TR_44 ;
	7'h29 :
		TR_233 = TR_44 ;
	7'h2a :
		TR_233 = TR_44 ;
	7'h2b :
		TR_233 = TR_44 ;
	7'h2c :
		TR_233 = TR_44 ;
	7'h2d :
		TR_233 = TR_44 ;
	7'h2e :
		TR_233 = TR_44 ;
	7'h2f :
		TR_233 = TR_44 ;
	7'h30 :
		TR_233 = TR_44 ;
	7'h31 :
		TR_233 = TR_44 ;
	7'h32 :
		TR_233 = TR_44 ;
	7'h33 :
		TR_233 = TR_44 ;
	7'h34 :
		TR_233 = TR_44 ;
	7'h35 :
		TR_233 = TR_44 ;
	7'h36 :
		TR_233 = TR_44 ;
	7'h37 :
		TR_233 = TR_44 ;
	7'h38 :
		TR_233 = TR_44 ;
	7'h39 :
		TR_233 = TR_44 ;
	7'h3a :
		TR_233 = TR_44 ;
	7'h3b :
		TR_233 = TR_44 ;
	7'h3c :
		TR_233 = TR_44 ;
	7'h3d :
		TR_233 = TR_44 ;
	7'h3e :
		TR_233 = TR_44 ;
	7'h3f :
		TR_233 = TR_44 ;
	7'h40 :
		TR_233 = TR_44 ;
	7'h41 :
		TR_233 = TR_44 ;
	7'h42 :
		TR_233 = TR_44 ;
	7'h43 :
		TR_233 = TR_44 ;
	7'h44 :
		TR_233 = TR_44 ;
	7'h45 :
		TR_233 = TR_44 ;
	7'h46 :
		TR_233 = TR_44 ;
	7'h47 :
		TR_233 = TR_44 ;
	7'h48 :
		TR_233 = TR_44 ;
	7'h49 :
		TR_233 = TR_44 ;
	7'h4a :
		TR_233 = TR_44 ;
	7'h4b :
		TR_233 = TR_44 ;
	7'h4c :
		TR_233 = TR_44 ;
	7'h4d :
		TR_233 = TR_44 ;
	7'h4e :
		TR_233 = TR_44 ;
	7'h4f :
		TR_233 = TR_44 ;
	7'h50 :
		TR_233 = TR_44 ;
	7'h51 :
		TR_233 = TR_44 ;
	7'h52 :
		TR_233 = TR_44 ;
	7'h53 :
		TR_233 = TR_44 ;
	7'h54 :
		TR_233 = TR_44 ;
	7'h55 :
		TR_233 = TR_44 ;
	7'h56 :
		TR_233 = TR_44 ;
	7'h57 :
		TR_233 = TR_44 ;
	7'h58 :
		TR_233 = TR_44 ;
	7'h59 :
		TR_233 = TR_44 ;
	7'h5a :
		TR_233 = TR_44 ;
	7'h5b :
		TR_233 = TR_44 ;
	7'h5c :
		TR_233 = TR_44 ;
	7'h5d :
		TR_233 = TR_44 ;
	7'h5e :
		TR_233 = TR_44 ;
	7'h5f :
		TR_233 = TR_44 ;
	7'h60 :
		TR_233 = TR_44 ;
	7'h61 :
		TR_233 = TR_44 ;
	7'h62 :
		TR_233 = TR_44 ;
	7'h63 :
		TR_233 = TR_44 ;
	7'h64 :
		TR_233 = TR_44 ;
	7'h65 :
		TR_233 = TR_44 ;
	7'h66 :
		TR_233 = TR_44 ;
	7'h67 :
		TR_233 = TR_44 ;
	7'h68 :
		TR_233 = TR_44 ;
	7'h69 :
		TR_233 = TR_44 ;
	7'h6a :
		TR_233 = TR_44 ;
	7'h6b :
		TR_233 = TR_44 ;
	7'h6c :
		TR_233 = TR_44 ;
	7'h6d :
		TR_233 = TR_44 ;
	7'h6e :
		TR_233 = TR_44 ;
	7'h6f :
		TR_233 = TR_44 ;
	7'h70 :
		TR_233 = TR_44 ;
	7'h71 :
		TR_233 = TR_44 ;
	7'h72 :
		TR_233 = TR_44 ;
	7'h73 :
		TR_233 = TR_44 ;
	7'h74 :
		TR_233 = TR_44 ;
	7'h75 :
		TR_233 = TR_44 ;
	7'h76 :
		TR_233 = TR_44 ;
	7'h77 :
		TR_233 = TR_44 ;
	7'h78 :
		TR_233 = TR_44 ;
	7'h79 :
		TR_233 = TR_44 ;
	7'h7a :
		TR_233 = TR_44 ;
	7'h7b :
		TR_233 = TR_44 ;
	7'h7c :
		TR_233 = TR_44 ;
	7'h7d :
		TR_233 = TR_44 ;
	7'h7e :
		TR_233 = TR_44 ;
	7'h7f :
		TR_233 = TR_44 ;
	default :
		TR_233 = 9'hx ;
	endcase
always @ ( TR_233 or U_173 or sub8u_71ot or U_183 or RG_rl_145 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_32_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h20 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_32_t = ( ( { 9{ M_180 } } & RG_rl_145 )
		| ( { 9{ U_173 } } & TR_233 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_32_en = ( M_180 | RG_rl_32_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_32_en )
		RG_rl_32 <= RG_rl_32_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_45 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_232 = TR_45 ;
	7'h01 :
		TR_232 = TR_45 ;
	7'h02 :
		TR_232 = TR_45 ;
	7'h03 :
		TR_232 = TR_45 ;
	7'h04 :
		TR_232 = TR_45 ;
	7'h05 :
		TR_232 = TR_45 ;
	7'h06 :
		TR_232 = TR_45 ;
	7'h07 :
		TR_232 = TR_45 ;
	7'h08 :
		TR_232 = TR_45 ;
	7'h09 :
		TR_232 = TR_45 ;
	7'h0a :
		TR_232 = TR_45 ;
	7'h0b :
		TR_232 = TR_45 ;
	7'h0c :
		TR_232 = TR_45 ;
	7'h0d :
		TR_232 = TR_45 ;
	7'h0e :
		TR_232 = TR_45 ;
	7'h0f :
		TR_232 = TR_45 ;
	7'h10 :
		TR_232 = TR_45 ;
	7'h11 :
		TR_232 = TR_45 ;
	7'h12 :
		TR_232 = TR_45 ;
	7'h13 :
		TR_232 = TR_45 ;
	7'h14 :
		TR_232 = TR_45 ;
	7'h15 :
		TR_232 = TR_45 ;
	7'h16 :
		TR_232 = TR_45 ;
	7'h17 :
		TR_232 = TR_45 ;
	7'h18 :
		TR_232 = TR_45 ;
	7'h19 :
		TR_232 = TR_45 ;
	7'h1a :
		TR_232 = TR_45 ;
	7'h1b :
		TR_232 = TR_45 ;
	7'h1c :
		TR_232 = TR_45 ;
	7'h1d :
		TR_232 = TR_45 ;
	7'h1e :
		TR_232 = TR_45 ;
	7'h1f :
		TR_232 = TR_45 ;
	7'h20 :
		TR_232 = TR_45 ;
	7'h21 :
		TR_232 = 9'h000 ;	// line#=../rle.cpp:80
	7'h22 :
		TR_232 = TR_45 ;
	7'h23 :
		TR_232 = TR_45 ;
	7'h24 :
		TR_232 = TR_45 ;
	7'h25 :
		TR_232 = TR_45 ;
	7'h26 :
		TR_232 = TR_45 ;
	7'h27 :
		TR_232 = TR_45 ;
	7'h28 :
		TR_232 = TR_45 ;
	7'h29 :
		TR_232 = TR_45 ;
	7'h2a :
		TR_232 = TR_45 ;
	7'h2b :
		TR_232 = TR_45 ;
	7'h2c :
		TR_232 = TR_45 ;
	7'h2d :
		TR_232 = TR_45 ;
	7'h2e :
		TR_232 = TR_45 ;
	7'h2f :
		TR_232 = TR_45 ;
	7'h30 :
		TR_232 = TR_45 ;
	7'h31 :
		TR_232 = TR_45 ;
	7'h32 :
		TR_232 = TR_45 ;
	7'h33 :
		TR_232 = TR_45 ;
	7'h34 :
		TR_232 = TR_45 ;
	7'h35 :
		TR_232 = TR_45 ;
	7'h36 :
		TR_232 = TR_45 ;
	7'h37 :
		TR_232 = TR_45 ;
	7'h38 :
		TR_232 = TR_45 ;
	7'h39 :
		TR_232 = TR_45 ;
	7'h3a :
		TR_232 = TR_45 ;
	7'h3b :
		TR_232 = TR_45 ;
	7'h3c :
		TR_232 = TR_45 ;
	7'h3d :
		TR_232 = TR_45 ;
	7'h3e :
		TR_232 = TR_45 ;
	7'h3f :
		TR_232 = TR_45 ;
	7'h40 :
		TR_232 = TR_45 ;
	7'h41 :
		TR_232 = TR_45 ;
	7'h42 :
		TR_232 = TR_45 ;
	7'h43 :
		TR_232 = TR_45 ;
	7'h44 :
		TR_232 = TR_45 ;
	7'h45 :
		TR_232 = TR_45 ;
	7'h46 :
		TR_232 = TR_45 ;
	7'h47 :
		TR_232 = TR_45 ;
	7'h48 :
		TR_232 = TR_45 ;
	7'h49 :
		TR_232 = TR_45 ;
	7'h4a :
		TR_232 = TR_45 ;
	7'h4b :
		TR_232 = TR_45 ;
	7'h4c :
		TR_232 = TR_45 ;
	7'h4d :
		TR_232 = TR_45 ;
	7'h4e :
		TR_232 = TR_45 ;
	7'h4f :
		TR_232 = TR_45 ;
	7'h50 :
		TR_232 = TR_45 ;
	7'h51 :
		TR_232 = TR_45 ;
	7'h52 :
		TR_232 = TR_45 ;
	7'h53 :
		TR_232 = TR_45 ;
	7'h54 :
		TR_232 = TR_45 ;
	7'h55 :
		TR_232 = TR_45 ;
	7'h56 :
		TR_232 = TR_45 ;
	7'h57 :
		TR_232 = TR_45 ;
	7'h58 :
		TR_232 = TR_45 ;
	7'h59 :
		TR_232 = TR_45 ;
	7'h5a :
		TR_232 = TR_45 ;
	7'h5b :
		TR_232 = TR_45 ;
	7'h5c :
		TR_232 = TR_45 ;
	7'h5d :
		TR_232 = TR_45 ;
	7'h5e :
		TR_232 = TR_45 ;
	7'h5f :
		TR_232 = TR_45 ;
	7'h60 :
		TR_232 = TR_45 ;
	7'h61 :
		TR_232 = TR_45 ;
	7'h62 :
		TR_232 = TR_45 ;
	7'h63 :
		TR_232 = TR_45 ;
	7'h64 :
		TR_232 = TR_45 ;
	7'h65 :
		TR_232 = TR_45 ;
	7'h66 :
		TR_232 = TR_45 ;
	7'h67 :
		TR_232 = TR_45 ;
	7'h68 :
		TR_232 = TR_45 ;
	7'h69 :
		TR_232 = TR_45 ;
	7'h6a :
		TR_232 = TR_45 ;
	7'h6b :
		TR_232 = TR_45 ;
	7'h6c :
		TR_232 = TR_45 ;
	7'h6d :
		TR_232 = TR_45 ;
	7'h6e :
		TR_232 = TR_45 ;
	7'h6f :
		TR_232 = TR_45 ;
	7'h70 :
		TR_232 = TR_45 ;
	7'h71 :
		TR_232 = TR_45 ;
	7'h72 :
		TR_232 = TR_45 ;
	7'h73 :
		TR_232 = TR_45 ;
	7'h74 :
		TR_232 = TR_45 ;
	7'h75 :
		TR_232 = TR_45 ;
	7'h76 :
		TR_232 = TR_45 ;
	7'h77 :
		TR_232 = TR_45 ;
	7'h78 :
		TR_232 = TR_45 ;
	7'h79 :
		TR_232 = TR_45 ;
	7'h7a :
		TR_232 = TR_45 ;
	7'h7b :
		TR_232 = TR_45 ;
	7'h7c :
		TR_232 = TR_45 ;
	7'h7d :
		TR_232 = TR_45 ;
	7'h7e :
		TR_232 = TR_45 ;
	7'h7f :
		TR_232 = TR_45 ;
	default :
		TR_232 = 9'hx ;
	endcase
always @ ( TR_232 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_14 or 
	U_174 or RG_rl_145 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_33_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h21 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_33_t = ( ( { 9{ ST1_03d } } & RG_rl_145 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_14 )
		| ( { 9{ U_173 } } & TR_232 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_33_en = ( ST1_03d | U_174 | RG_rl_33_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_33_en )
		RG_rl_33 <= RG_rl_33_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_46 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_231 = TR_46 ;
	7'h01 :
		TR_231 = TR_46 ;
	7'h02 :
		TR_231 = TR_46 ;
	7'h03 :
		TR_231 = TR_46 ;
	7'h04 :
		TR_231 = TR_46 ;
	7'h05 :
		TR_231 = TR_46 ;
	7'h06 :
		TR_231 = TR_46 ;
	7'h07 :
		TR_231 = TR_46 ;
	7'h08 :
		TR_231 = TR_46 ;
	7'h09 :
		TR_231 = TR_46 ;
	7'h0a :
		TR_231 = TR_46 ;
	7'h0b :
		TR_231 = TR_46 ;
	7'h0c :
		TR_231 = TR_46 ;
	7'h0d :
		TR_231 = TR_46 ;
	7'h0e :
		TR_231 = TR_46 ;
	7'h0f :
		TR_231 = TR_46 ;
	7'h10 :
		TR_231 = TR_46 ;
	7'h11 :
		TR_231 = TR_46 ;
	7'h12 :
		TR_231 = TR_46 ;
	7'h13 :
		TR_231 = TR_46 ;
	7'h14 :
		TR_231 = TR_46 ;
	7'h15 :
		TR_231 = TR_46 ;
	7'h16 :
		TR_231 = TR_46 ;
	7'h17 :
		TR_231 = TR_46 ;
	7'h18 :
		TR_231 = TR_46 ;
	7'h19 :
		TR_231 = TR_46 ;
	7'h1a :
		TR_231 = TR_46 ;
	7'h1b :
		TR_231 = TR_46 ;
	7'h1c :
		TR_231 = TR_46 ;
	7'h1d :
		TR_231 = TR_46 ;
	7'h1e :
		TR_231 = TR_46 ;
	7'h1f :
		TR_231 = TR_46 ;
	7'h20 :
		TR_231 = TR_46 ;
	7'h21 :
		TR_231 = TR_46 ;
	7'h22 :
		TR_231 = 9'h000 ;	// line#=../rle.cpp:80
	7'h23 :
		TR_231 = TR_46 ;
	7'h24 :
		TR_231 = TR_46 ;
	7'h25 :
		TR_231 = TR_46 ;
	7'h26 :
		TR_231 = TR_46 ;
	7'h27 :
		TR_231 = TR_46 ;
	7'h28 :
		TR_231 = TR_46 ;
	7'h29 :
		TR_231 = TR_46 ;
	7'h2a :
		TR_231 = TR_46 ;
	7'h2b :
		TR_231 = TR_46 ;
	7'h2c :
		TR_231 = TR_46 ;
	7'h2d :
		TR_231 = TR_46 ;
	7'h2e :
		TR_231 = TR_46 ;
	7'h2f :
		TR_231 = TR_46 ;
	7'h30 :
		TR_231 = TR_46 ;
	7'h31 :
		TR_231 = TR_46 ;
	7'h32 :
		TR_231 = TR_46 ;
	7'h33 :
		TR_231 = TR_46 ;
	7'h34 :
		TR_231 = TR_46 ;
	7'h35 :
		TR_231 = TR_46 ;
	7'h36 :
		TR_231 = TR_46 ;
	7'h37 :
		TR_231 = TR_46 ;
	7'h38 :
		TR_231 = TR_46 ;
	7'h39 :
		TR_231 = TR_46 ;
	7'h3a :
		TR_231 = TR_46 ;
	7'h3b :
		TR_231 = TR_46 ;
	7'h3c :
		TR_231 = TR_46 ;
	7'h3d :
		TR_231 = TR_46 ;
	7'h3e :
		TR_231 = TR_46 ;
	7'h3f :
		TR_231 = TR_46 ;
	7'h40 :
		TR_231 = TR_46 ;
	7'h41 :
		TR_231 = TR_46 ;
	7'h42 :
		TR_231 = TR_46 ;
	7'h43 :
		TR_231 = TR_46 ;
	7'h44 :
		TR_231 = TR_46 ;
	7'h45 :
		TR_231 = TR_46 ;
	7'h46 :
		TR_231 = TR_46 ;
	7'h47 :
		TR_231 = TR_46 ;
	7'h48 :
		TR_231 = TR_46 ;
	7'h49 :
		TR_231 = TR_46 ;
	7'h4a :
		TR_231 = TR_46 ;
	7'h4b :
		TR_231 = TR_46 ;
	7'h4c :
		TR_231 = TR_46 ;
	7'h4d :
		TR_231 = TR_46 ;
	7'h4e :
		TR_231 = TR_46 ;
	7'h4f :
		TR_231 = TR_46 ;
	7'h50 :
		TR_231 = TR_46 ;
	7'h51 :
		TR_231 = TR_46 ;
	7'h52 :
		TR_231 = TR_46 ;
	7'h53 :
		TR_231 = TR_46 ;
	7'h54 :
		TR_231 = TR_46 ;
	7'h55 :
		TR_231 = TR_46 ;
	7'h56 :
		TR_231 = TR_46 ;
	7'h57 :
		TR_231 = TR_46 ;
	7'h58 :
		TR_231 = TR_46 ;
	7'h59 :
		TR_231 = TR_46 ;
	7'h5a :
		TR_231 = TR_46 ;
	7'h5b :
		TR_231 = TR_46 ;
	7'h5c :
		TR_231 = TR_46 ;
	7'h5d :
		TR_231 = TR_46 ;
	7'h5e :
		TR_231 = TR_46 ;
	7'h5f :
		TR_231 = TR_46 ;
	7'h60 :
		TR_231 = TR_46 ;
	7'h61 :
		TR_231 = TR_46 ;
	7'h62 :
		TR_231 = TR_46 ;
	7'h63 :
		TR_231 = TR_46 ;
	7'h64 :
		TR_231 = TR_46 ;
	7'h65 :
		TR_231 = TR_46 ;
	7'h66 :
		TR_231 = TR_46 ;
	7'h67 :
		TR_231 = TR_46 ;
	7'h68 :
		TR_231 = TR_46 ;
	7'h69 :
		TR_231 = TR_46 ;
	7'h6a :
		TR_231 = TR_46 ;
	7'h6b :
		TR_231 = TR_46 ;
	7'h6c :
		TR_231 = TR_46 ;
	7'h6d :
		TR_231 = TR_46 ;
	7'h6e :
		TR_231 = TR_46 ;
	7'h6f :
		TR_231 = TR_46 ;
	7'h70 :
		TR_231 = TR_46 ;
	7'h71 :
		TR_231 = TR_46 ;
	7'h72 :
		TR_231 = TR_46 ;
	7'h73 :
		TR_231 = TR_46 ;
	7'h74 :
		TR_231 = TR_46 ;
	7'h75 :
		TR_231 = TR_46 ;
	7'h76 :
		TR_231 = TR_46 ;
	7'h77 :
		TR_231 = TR_46 ;
	7'h78 :
		TR_231 = TR_46 ;
	7'h79 :
		TR_231 = TR_46 ;
	7'h7a :
		TR_231 = TR_46 ;
	7'h7b :
		TR_231 = TR_46 ;
	7'h7c :
		TR_231 = TR_46 ;
	7'h7d :
		TR_231 = TR_46 ;
	7'h7e :
		TR_231 = TR_46 ;
	7'h7f :
		TR_231 = TR_46 ;
	default :
		TR_231 = 9'hx ;
	endcase
always @ ( TR_231 or U_173 or sub8u_71ot or U_183 or RG_rl_146 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_34_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h22 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_34_t = ( ( { 9{ M_180 } } & RG_rl_146 )
		| ( { 9{ U_173 } } & TR_231 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_34_en = ( M_180 | RG_rl_34_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_34_en )
		RG_rl_34 <= RG_rl_34_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_47 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_230 = TR_47 ;
	7'h01 :
		TR_230 = TR_47 ;
	7'h02 :
		TR_230 = TR_47 ;
	7'h03 :
		TR_230 = TR_47 ;
	7'h04 :
		TR_230 = TR_47 ;
	7'h05 :
		TR_230 = TR_47 ;
	7'h06 :
		TR_230 = TR_47 ;
	7'h07 :
		TR_230 = TR_47 ;
	7'h08 :
		TR_230 = TR_47 ;
	7'h09 :
		TR_230 = TR_47 ;
	7'h0a :
		TR_230 = TR_47 ;
	7'h0b :
		TR_230 = TR_47 ;
	7'h0c :
		TR_230 = TR_47 ;
	7'h0d :
		TR_230 = TR_47 ;
	7'h0e :
		TR_230 = TR_47 ;
	7'h0f :
		TR_230 = TR_47 ;
	7'h10 :
		TR_230 = TR_47 ;
	7'h11 :
		TR_230 = TR_47 ;
	7'h12 :
		TR_230 = TR_47 ;
	7'h13 :
		TR_230 = TR_47 ;
	7'h14 :
		TR_230 = TR_47 ;
	7'h15 :
		TR_230 = TR_47 ;
	7'h16 :
		TR_230 = TR_47 ;
	7'h17 :
		TR_230 = TR_47 ;
	7'h18 :
		TR_230 = TR_47 ;
	7'h19 :
		TR_230 = TR_47 ;
	7'h1a :
		TR_230 = TR_47 ;
	7'h1b :
		TR_230 = TR_47 ;
	7'h1c :
		TR_230 = TR_47 ;
	7'h1d :
		TR_230 = TR_47 ;
	7'h1e :
		TR_230 = TR_47 ;
	7'h1f :
		TR_230 = TR_47 ;
	7'h20 :
		TR_230 = TR_47 ;
	7'h21 :
		TR_230 = TR_47 ;
	7'h22 :
		TR_230 = TR_47 ;
	7'h23 :
		TR_230 = 9'h000 ;	// line#=../rle.cpp:80
	7'h24 :
		TR_230 = TR_47 ;
	7'h25 :
		TR_230 = TR_47 ;
	7'h26 :
		TR_230 = TR_47 ;
	7'h27 :
		TR_230 = TR_47 ;
	7'h28 :
		TR_230 = TR_47 ;
	7'h29 :
		TR_230 = TR_47 ;
	7'h2a :
		TR_230 = TR_47 ;
	7'h2b :
		TR_230 = TR_47 ;
	7'h2c :
		TR_230 = TR_47 ;
	7'h2d :
		TR_230 = TR_47 ;
	7'h2e :
		TR_230 = TR_47 ;
	7'h2f :
		TR_230 = TR_47 ;
	7'h30 :
		TR_230 = TR_47 ;
	7'h31 :
		TR_230 = TR_47 ;
	7'h32 :
		TR_230 = TR_47 ;
	7'h33 :
		TR_230 = TR_47 ;
	7'h34 :
		TR_230 = TR_47 ;
	7'h35 :
		TR_230 = TR_47 ;
	7'h36 :
		TR_230 = TR_47 ;
	7'h37 :
		TR_230 = TR_47 ;
	7'h38 :
		TR_230 = TR_47 ;
	7'h39 :
		TR_230 = TR_47 ;
	7'h3a :
		TR_230 = TR_47 ;
	7'h3b :
		TR_230 = TR_47 ;
	7'h3c :
		TR_230 = TR_47 ;
	7'h3d :
		TR_230 = TR_47 ;
	7'h3e :
		TR_230 = TR_47 ;
	7'h3f :
		TR_230 = TR_47 ;
	7'h40 :
		TR_230 = TR_47 ;
	7'h41 :
		TR_230 = TR_47 ;
	7'h42 :
		TR_230 = TR_47 ;
	7'h43 :
		TR_230 = TR_47 ;
	7'h44 :
		TR_230 = TR_47 ;
	7'h45 :
		TR_230 = TR_47 ;
	7'h46 :
		TR_230 = TR_47 ;
	7'h47 :
		TR_230 = TR_47 ;
	7'h48 :
		TR_230 = TR_47 ;
	7'h49 :
		TR_230 = TR_47 ;
	7'h4a :
		TR_230 = TR_47 ;
	7'h4b :
		TR_230 = TR_47 ;
	7'h4c :
		TR_230 = TR_47 ;
	7'h4d :
		TR_230 = TR_47 ;
	7'h4e :
		TR_230 = TR_47 ;
	7'h4f :
		TR_230 = TR_47 ;
	7'h50 :
		TR_230 = TR_47 ;
	7'h51 :
		TR_230 = TR_47 ;
	7'h52 :
		TR_230 = TR_47 ;
	7'h53 :
		TR_230 = TR_47 ;
	7'h54 :
		TR_230 = TR_47 ;
	7'h55 :
		TR_230 = TR_47 ;
	7'h56 :
		TR_230 = TR_47 ;
	7'h57 :
		TR_230 = TR_47 ;
	7'h58 :
		TR_230 = TR_47 ;
	7'h59 :
		TR_230 = TR_47 ;
	7'h5a :
		TR_230 = TR_47 ;
	7'h5b :
		TR_230 = TR_47 ;
	7'h5c :
		TR_230 = TR_47 ;
	7'h5d :
		TR_230 = TR_47 ;
	7'h5e :
		TR_230 = TR_47 ;
	7'h5f :
		TR_230 = TR_47 ;
	7'h60 :
		TR_230 = TR_47 ;
	7'h61 :
		TR_230 = TR_47 ;
	7'h62 :
		TR_230 = TR_47 ;
	7'h63 :
		TR_230 = TR_47 ;
	7'h64 :
		TR_230 = TR_47 ;
	7'h65 :
		TR_230 = TR_47 ;
	7'h66 :
		TR_230 = TR_47 ;
	7'h67 :
		TR_230 = TR_47 ;
	7'h68 :
		TR_230 = TR_47 ;
	7'h69 :
		TR_230 = TR_47 ;
	7'h6a :
		TR_230 = TR_47 ;
	7'h6b :
		TR_230 = TR_47 ;
	7'h6c :
		TR_230 = TR_47 ;
	7'h6d :
		TR_230 = TR_47 ;
	7'h6e :
		TR_230 = TR_47 ;
	7'h6f :
		TR_230 = TR_47 ;
	7'h70 :
		TR_230 = TR_47 ;
	7'h71 :
		TR_230 = TR_47 ;
	7'h72 :
		TR_230 = TR_47 ;
	7'h73 :
		TR_230 = TR_47 ;
	7'h74 :
		TR_230 = TR_47 ;
	7'h75 :
		TR_230 = TR_47 ;
	7'h76 :
		TR_230 = TR_47 ;
	7'h77 :
		TR_230 = TR_47 ;
	7'h78 :
		TR_230 = TR_47 ;
	7'h79 :
		TR_230 = TR_47 ;
	7'h7a :
		TR_230 = TR_47 ;
	7'h7b :
		TR_230 = TR_47 ;
	7'h7c :
		TR_230 = TR_47 ;
	7'h7d :
		TR_230 = TR_47 ;
	7'h7e :
		TR_230 = TR_47 ;
	7'h7f :
		TR_230 = TR_47 ;
	default :
		TR_230 = 9'hx ;
	endcase
always @ ( TR_230 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_15 or 
	U_174 or RG_rl_146 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_35_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h23 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_35_t = ( ( { 9{ ST1_03d } } & RG_rl_146 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_15 )
		| ( { 9{ U_173 } } & TR_230 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_35_en = ( ST1_03d | U_174 | RG_rl_35_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_35_en )
		RG_rl_35 <= RG_rl_35_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_48 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_229 = TR_48 ;
	7'h01 :
		TR_229 = TR_48 ;
	7'h02 :
		TR_229 = TR_48 ;
	7'h03 :
		TR_229 = TR_48 ;
	7'h04 :
		TR_229 = TR_48 ;
	7'h05 :
		TR_229 = TR_48 ;
	7'h06 :
		TR_229 = TR_48 ;
	7'h07 :
		TR_229 = TR_48 ;
	7'h08 :
		TR_229 = TR_48 ;
	7'h09 :
		TR_229 = TR_48 ;
	7'h0a :
		TR_229 = TR_48 ;
	7'h0b :
		TR_229 = TR_48 ;
	7'h0c :
		TR_229 = TR_48 ;
	7'h0d :
		TR_229 = TR_48 ;
	7'h0e :
		TR_229 = TR_48 ;
	7'h0f :
		TR_229 = TR_48 ;
	7'h10 :
		TR_229 = TR_48 ;
	7'h11 :
		TR_229 = TR_48 ;
	7'h12 :
		TR_229 = TR_48 ;
	7'h13 :
		TR_229 = TR_48 ;
	7'h14 :
		TR_229 = TR_48 ;
	7'h15 :
		TR_229 = TR_48 ;
	7'h16 :
		TR_229 = TR_48 ;
	7'h17 :
		TR_229 = TR_48 ;
	7'h18 :
		TR_229 = TR_48 ;
	7'h19 :
		TR_229 = TR_48 ;
	7'h1a :
		TR_229 = TR_48 ;
	7'h1b :
		TR_229 = TR_48 ;
	7'h1c :
		TR_229 = TR_48 ;
	7'h1d :
		TR_229 = TR_48 ;
	7'h1e :
		TR_229 = TR_48 ;
	7'h1f :
		TR_229 = TR_48 ;
	7'h20 :
		TR_229 = TR_48 ;
	7'h21 :
		TR_229 = TR_48 ;
	7'h22 :
		TR_229 = TR_48 ;
	7'h23 :
		TR_229 = TR_48 ;
	7'h24 :
		TR_229 = 9'h000 ;	// line#=../rle.cpp:80
	7'h25 :
		TR_229 = TR_48 ;
	7'h26 :
		TR_229 = TR_48 ;
	7'h27 :
		TR_229 = TR_48 ;
	7'h28 :
		TR_229 = TR_48 ;
	7'h29 :
		TR_229 = TR_48 ;
	7'h2a :
		TR_229 = TR_48 ;
	7'h2b :
		TR_229 = TR_48 ;
	7'h2c :
		TR_229 = TR_48 ;
	7'h2d :
		TR_229 = TR_48 ;
	7'h2e :
		TR_229 = TR_48 ;
	7'h2f :
		TR_229 = TR_48 ;
	7'h30 :
		TR_229 = TR_48 ;
	7'h31 :
		TR_229 = TR_48 ;
	7'h32 :
		TR_229 = TR_48 ;
	7'h33 :
		TR_229 = TR_48 ;
	7'h34 :
		TR_229 = TR_48 ;
	7'h35 :
		TR_229 = TR_48 ;
	7'h36 :
		TR_229 = TR_48 ;
	7'h37 :
		TR_229 = TR_48 ;
	7'h38 :
		TR_229 = TR_48 ;
	7'h39 :
		TR_229 = TR_48 ;
	7'h3a :
		TR_229 = TR_48 ;
	7'h3b :
		TR_229 = TR_48 ;
	7'h3c :
		TR_229 = TR_48 ;
	7'h3d :
		TR_229 = TR_48 ;
	7'h3e :
		TR_229 = TR_48 ;
	7'h3f :
		TR_229 = TR_48 ;
	7'h40 :
		TR_229 = TR_48 ;
	7'h41 :
		TR_229 = TR_48 ;
	7'h42 :
		TR_229 = TR_48 ;
	7'h43 :
		TR_229 = TR_48 ;
	7'h44 :
		TR_229 = TR_48 ;
	7'h45 :
		TR_229 = TR_48 ;
	7'h46 :
		TR_229 = TR_48 ;
	7'h47 :
		TR_229 = TR_48 ;
	7'h48 :
		TR_229 = TR_48 ;
	7'h49 :
		TR_229 = TR_48 ;
	7'h4a :
		TR_229 = TR_48 ;
	7'h4b :
		TR_229 = TR_48 ;
	7'h4c :
		TR_229 = TR_48 ;
	7'h4d :
		TR_229 = TR_48 ;
	7'h4e :
		TR_229 = TR_48 ;
	7'h4f :
		TR_229 = TR_48 ;
	7'h50 :
		TR_229 = TR_48 ;
	7'h51 :
		TR_229 = TR_48 ;
	7'h52 :
		TR_229 = TR_48 ;
	7'h53 :
		TR_229 = TR_48 ;
	7'h54 :
		TR_229 = TR_48 ;
	7'h55 :
		TR_229 = TR_48 ;
	7'h56 :
		TR_229 = TR_48 ;
	7'h57 :
		TR_229 = TR_48 ;
	7'h58 :
		TR_229 = TR_48 ;
	7'h59 :
		TR_229 = TR_48 ;
	7'h5a :
		TR_229 = TR_48 ;
	7'h5b :
		TR_229 = TR_48 ;
	7'h5c :
		TR_229 = TR_48 ;
	7'h5d :
		TR_229 = TR_48 ;
	7'h5e :
		TR_229 = TR_48 ;
	7'h5f :
		TR_229 = TR_48 ;
	7'h60 :
		TR_229 = TR_48 ;
	7'h61 :
		TR_229 = TR_48 ;
	7'h62 :
		TR_229 = TR_48 ;
	7'h63 :
		TR_229 = TR_48 ;
	7'h64 :
		TR_229 = TR_48 ;
	7'h65 :
		TR_229 = TR_48 ;
	7'h66 :
		TR_229 = TR_48 ;
	7'h67 :
		TR_229 = TR_48 ;
	7'h68 :
		TR_229 = TR_48 ;
	7'h69 :
		TR_229 = TR_48 ;
	7'h6a :
		TR_229 = TR_48 ;
	7'h6b :
		TR_229 = TR_48 ;
	7'h6c :
		TR_229 = TR_48 ;
	7'h6d :
		TR_229 = TR_48 ;
	7'h6e :
		TR_229 = TR_48 ;
	7'h6f :
		TR_229 = TR_48 ;
	7'h70 :
		TR_229 = TR_48 ;
	7'h71 :
		TR_229 = TR_48 ;
	7'h72 :
		TR_229 = TR_48 ;
	7'h73 :
		TR_229 = TR_48 ;
	7'h74 :
		TR_229 = TR_48 ;
	7'h75 :
		TR_229 = TR_48 ;
	7'h76 :
		TR_229 = TR_48 ;
	7'h77 :
		TR_229 = TR_48 ;
	7'h78 :
		TR_229 = TR_48 ;
	7'h79 :
		TR_229 = TR_48 ;
	7'h7a :
		TR_229 = TR_48 ;
	7'h7b :
		TR_229 = TR_48 ;
	7'h7c :
		TR_229 = TR_48 ;
	7'h7d :
		TR_229 = TR_48 ;
	7'h7e :
		TR_229 = TR_48 ;
	7'h7f :
		TR_229 = TR_48 ;
	default :
		TR_229 = 9'hx ;
	endcase
always @ ( TR_229 or U_173 or sub8u_71ot or U_183 or RG_rl_147 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_36_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h24 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_36_t = ( ( { 9{ M_180 } } & RG_rl_147 )
		| ( { 9{ U_173 } } & TR_229 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_36_en = ( M_180 | RG_rl_36_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_36_en )
		RG_rl_36 <= RG_rl_36_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_49 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_228 = TR_49 ;
	7'h01 :
		TR_228 = TR_49 ;
	7'h02 :
		TR_228 = TR_49 ;
	7'h03 :
		TR_228 = TR_49 ;
	7'h04 :
		TR_228 = TR_49 ;
	7'h05 :
		TR_228 = TR_49 ;
	7'h06 :
		TR_228 = TR_49 ;
	7'h07 :
		TR_228 = TR_49 ;
	7'h08 :
		TR_228 = TR_49 ;
	7'h09 :
		TR_228 = TR_49 ;
	7'h0a :
		TR_228 = TR_49 ;
	7'h0b :
		TR_228 = TR_49 ;
	7'h0c :
		TR_228 = TR_49 ;
	7'h0d :
		TR_228 = TR_49 ;
	7'h0e :
		TR_228 = TR_49 ;
	7'h0f :
		TR_228 = TR_49 ;
	7'h10 :
		TR_228 = TR_49 ;
	7'h11 :
		TR_228 = TR_49 ;
	7'h12 :
		TR_228 = TR_49 ;
	7'h13 :
		TR_228 = TR_49 ;
	7'h14 :
		TR_228 = TR_49 ;
	7'h15 :
		TR_228 = TR_49 ;
	7'h16 :
		TR_228 = TR_49 ;
	7'h17 :
		TR_228 = TR_49 ;
	7'h18 :
		TR_228 = TR_49 ;
	7'h19 :
		TR_228 = TR_49 ;
	7'h1a :
		TR_228 = TR_49 ;
	7'h1b :
		TR_228 = TR_49 ;
	7'h1c :
		TR_228 = TR_49 ;
	7'h1d :
		TR_228 = TR_49 ;
	7'h1e :
		TR_228 = TR_49 ;
	7'h1f :
		TR_228 = TR_49 ;
	7'h20 :
		TR_228 = TR_49 ;
	7'h21 :
		TR_228 = TR_49 ;
	7'h22 :
		TR_228 = TR_49 ;
	7'h23 :
		TR_228 = TR_49 ;
	7'h24 :
		TR_228 = TR_49 ;
	7'h25 :
		TR_228 = 9'h000 ;	// line#=../rle.cpp:80
	7'h26 :
		TR_228 = TR_49 ;
	7'h27 :
		TR_228 = TR_49 ;
	7'h28 :
		TR_228 = TR_49 ;
	7'h29 :
		TR_228 = TR_49 ;
	7'h2a :
		TR_228 = TR_49 ;
	7'h2b :
		TR_228 = TR_49 ;
	7'h2c :
		TR_228 = TR_49 ;
	7'h2d :
		TR_228 = TR_49 ;
	7'h2e :
		TR_228 = TR_49 ;
	7'h2f :
		TR_228 = TR_49 ;
	7'h30 :
		TR_228 = TR_49 ;
	7'h31 :
		TR_228 = TR_49 ;
	7'h32 :
		TR_228 = TR_49 ;
	7'h33 :
		TR_228 = TR_49 ;
	7'h34 :
		TR_228 = TR_49 ;
	7'h35 :
		TR_228 = TR_49 ;
	7'h36 :
		TR_228 = TR_49 ;
	7'h37 :
		TR_228 = TR_49 ;
	7'h38 :
		TR_228 = TR_49 ;
	7'h39 :
		TR_228 = TR_49 ;
	7'h3a :
		TR_228 = TR_49 ;
	7'h3b :
		TR_228 = TR_49 ;
	7'h3c :
		TR_228 = TR_49 ;
	7'h3d :
		TR_228 = TR_49 ;
	7'h3e :
		TR_228 = TR_49 ;
	7'h3f :
		TR_228 = TR_49 ;
	7'h40 :
		TR_228 = TR_49 ;
	7'h41 :
		TR_228 = TR_49 ;
	7'h42 :
		TR_228 = TR_49 ;
	7'h43 :
		TR_228 = TR_49 ;
	7'h44 :
		TR_228 = TR_49 ;
	7'h45 :
		TR_228 = TR_49 ;
	7'h46 :
		TR_228 = TR_49 ;
	7'h47 :
		TR_228 = TR_49 ;
	7'h48 :
		TR_228 = TR_49 ;
	7'h49 :
		TR_228 = TR_49 ;
	7'h4a :
		TR_228 = TR_49 ;
	7'h4b :
		TR_228 = TR_49 ;
	7'h4c :
		TR_228 = TR_49 ;
	7'h4d :
		TR_228 = TR_49 ;
	7'h4e :
		TR_228 = TR_49 ;
	7'h4f :
		TR_228 = TR_49 ;
	7'h50 :
		TR_228 = TR_49 ;
	7'h51 :
		TR_228 = TR_49 ;
	7'h52 :
		TR_228 = TR_49 ;
	7'h53 :
		TR_228 = TR_49 ;
	7'h54 :
		TR_228 = TR_49 ;
	7'h55 :
		TR_228 = TR_49 ;
	7'h56 :
		TR_228 = TR_49 ;
	7'h57 :
		TR_228 = TR_49 ;
	7'h58 :
		TR_228 = TR_49 ;
	7'h59 :
		TR_228 = TR_49 ;
	7'h5a :
		TR_228 = TR_49 ;
	7'h5b :
		TR_228 = TR_49 ;
	7'h5c :
		TR_228 = TR_49 ;
	7'h5d :
		TR_228 = TR_49 ;
	7'h5e :
		TR_228 = TR_49 ;
	7'h5f :
		TR_228 = TR_49 ;
	7'h60 :
		TR_228 = TR_49 ;
	7'h61 :
		TR_228 = TR_49 ;
	7'h62 :
		TR_228 = TR_49 ;
	7'h63 :
		TR_228 = TR_49 ;
	7'h64 :
		TR_228 = TR_49 ;
	7'h65 :
		TR_228 = TR_49 ;
	7'h66 :
		TR_228 = TR_49 ;
	7'h67 :
		TR_228 = TR_49 ;
	7'h68 :
		TR_228 = TR_49 ;
	7'h69 :
		TR_228 = TR_49 ;
	7'h6a :
		TR_228 = TR_49 ;
	7'h6b :
		TR_228 = TR_49 ;
	7'h6c :
		TR_228 = TR_49 ;
	7'h6d :
		TR_228 = TR_49 ;
	7'h6e :
		TR_228 = TR_49 ;
	7'h6f :
		TR_228 = TR_49 ;
	7'h70 :
		TR_228 = TR_49 ;
	7'h71 :
		TR_228 = TR_49 ;
	7'h72 :
		TR_228 = TR_49 ;
	7'h73 :
		TR_228 = TR_49 ;
	7'h74 :
		TR_228 = TR_49 ;
	7'h75 :
		TR_228 = TR_49 ;
	7'h76 :
		TR_228 = TR_49 ;
	7'h77 :
		TR_228 = TR_49 ;
	7'h78 :
		TR_228 = TR_49 ;
	7'h79 :
		TR_228 = TR_49 ;
	7'h7a :
		TR_228 = TR_49 ;
	7'h7b :
		TR_228 = TR_49 ;
	7'h7c :
		TR_228 = TR_49 ;
	7'h7d :
		TR_228 = TR_49 ;
	7'h7e :
		TR_228 = TR_49 ;
	7'h7f :
		TR_228 = TR_49 ;
	default :
		TR_228 = 9'hx ;
	endcase
always @ ( TR_228 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_16 or 
	U_174 or RG_rl_147 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_37_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h25 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_37_t = ( ( { 9{ ST1_03d } } & RG_rl_147 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_16 )
		| ( { 9{ U_173 } } & TR_228 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_37_en = ( ST1_03d | U_174 | RG_rl_37_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_37_en )
		RG_rl_37 <= RG_rl_37_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_50 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_227 = TR_50 ;
	7'h01 :
		TR_227 = TR_50 ;
	7'h02 :
		TR_227 = TR_50 ;
	7'h03 :
		TR_227 = TR_50 ;
	7'h04 :
		TR_227 = TR_50 ;
	7'h05 :
		TR_227 = TR_50 ;
	7'h06 :
		TR_227 = TR_50 ;
	7'h07 :
		TR_227 = TR_50 ;
	7'h08 :
		TR_227 = TR_50 ;
	7'h09 :
		TR_227 = TR_50 ;
	7'h0a :
		TR_227 = TR_50 ;
	7'h0b :
		TR_227 = TR_50 ;
	7'h0c :
		TR_227 = TR_50 ;
	7'h0d :
		TR_227 = TR_50 ;
	7'h0e :
		TR_227 = TR_50 ;
	7'h0f :
		TR_227 = TR_50 ;
	7'h10 :
		TR_227 = TR_50 ;
	7'h11 :
		TR_227 = TR_50 ;
	7'h12 :
		TR_227 = TR_50 ;
	7'h13 :
		TR_227 = TR_50 ;
	7'h14 :
		TR_227 = TR_50 ;
	7'h15 :
		TR_227 = TR_50 ;
	7'h16 :
		TR_227 = TR_50 ;
	7'h17 :
		TR_227 = TR_50 ;
	7'h18 :
		TR_227 = TR_50 ;
	7'h19 :
		TR_227 = TR_50 ;
	7'h1a :
		TR_227 = TR_50 ;
	7'h1b :
		TR_227 = TR_50 ;
	7'h1c :
		TR_227 = TR_50 ;
	7'h1d :
		TR_227 = TR_50 ;
	7'h1e :
		TR_227 = TR_50 ;
	7'h1f :
		TR_227 = TR_50 ;
	7'h20 :
		TR_227 = TR_50 ;
	7'h21 :
		TR_227 = TR_50 ;
	7'h22 :
		TR_227 = TR_50 ;
	7'h23 :
		TR_227 = TR_50 ;
	7'h24 :
		TR_227 = TR_50 ;
	7'h25 :
		TR_227 = TR_50 ;
	7'h26 :
		TR_227 = 9'h000 ;	// line#=../rle.cpp:80
	7'h27 :
		TR_227 = TR_50 ;
	7'h28 :
		TR_227 = TR_50 ;
	7'h29 :
		TR_227 = TR_50 ;
	7'h2a :
		TR_227 = TR_50 ;
	7'h2b :
		TR_227 = TR_50 ;
	7'h2c :
		TR_227 = TR_50 ;
	7'h2d :
		TR_227 = TR_50 ;
	7'h2e :
		TR_227 = TR_50 ;
	7'h2f :
		TR_227 = TR_50 ;
	7'h30 :
		TR_227 = TR_50 ;
	7'h31 :
		TR_227 = TR_50 ;
	7'h32 :
		TR_227 = TR_50 ;
	7'h33 :
		TR_227 = TR_50 ;
	7'h34 :
		TR_227 = TR_50 ;
	7'h35 :
		TR_227 = TR_50 ;
	7'h36 :
		TR_227 = TR_50 ;
	7'h37 :
		TR_227 = TR_50 ;
	7'h38 :
		TR_227 = TR_50 ;
	7'h39 :
		TR_227 = TR_50 ;
	7'h3a :
		TR_227 = TR_50 ;
	7'h3b :
		TR_227 = TR_50 ;
	7'h3c :
		TR_227 = TR_50 ;
	7'h3d :
		TR_227 = TR_50 ;
	7'h3e :
		TR_227 = TR_50 ;
	7'h3f :
		TR_227 = TR_50 ;
	7'h40 :
		TR_227 = TR_50 ;
	7'h41 :
		TR_227 = TR_50 ;
	7'h42 :
		TR_227 = TR_50 ;
	7'h43 :
		TR_227 = TR_50 ;
	7'h44 :
		TR_227 = TR_50 ;
	7'h45 :
		TR_227 = TR_50 ;
	7'h46 :
		TR_227 = TR_50 ;
	7'h47 :
		TR_227 = TR_50 ;
	7'h48 :
		TR_227 = TR_50 ;
	7'h49 :
		TR_227 = TR_50 ;
	7'h4a :
		TR_227 = TR_50 ;
	7'h4b :
		TR_227 = TR_50 ;
	7'h4c :
		TR_227 = TR_50 ;
	7'h4d :
		TR_227 = TR_50 ;
	7'h4e :
		TR_227 = TR_50 ;
	7'h4f :
		TR_227 = TR_50 ;
	7'h50 :
		TR_227 = TR_50 ;
	7'h51 :
		TR_227 = TR_50 ;
	7'h52 :
		TR_227 = TR_50 ;
	7'h53 :
		TR_227 = TR_50 ;
	7'h54 :
		TR_227 = TR_50 ;
	7'h55 :
		TR_227 = TR_50 ;
	7'h56 :
		TR_227 = TR_50 ;
	7'h57 :
		TR_227 = TR_50 ;
	7'h58 :
		TR_227 = TR_50 ;
	7'h59 :
		TR_227 = TR_50 ;
	7'h5a :
		TR_227 = TR_50 ;
	7'h5b :
		TR_227 = TR_50 ;
	7'h5c :
		TR_227 = TR_50 ;
	7'h5d :
		TR_227 = TR_50 ;
	7'h5e :
		TR_227 = TR_50 ;
	7'h5f :
		TR_227 = TR_50 ;
	7'h60 :
		TR_227 = TR_50 ;
	7'h61 :
		TR_227 = TR_50 ;
	7'h62 :
		TR_227 = TR_50 ;
	7'h63 :
		TR_227 = TR_50 ;
	7'h64 :
		TR_227 = TR_50 ;
	7'h65 :
		TR_227 = TR_50 ;
	7'h66 :
		TR_227 = TR_50 ;
	7'h67 :
		TR_227 = TR_50 ;
	7'h68 :
		TR_227 = TR_50 ;
	7'h69 :
		TR_227 = TR_50 ;
	7'h6a :
		TR_227 = TR_50 ;
	7'h6b :
		TR_227 = TR_50 ;
	7'h6c :
		TR_227 = TR_50 ;
	7'h6d :
		TR_227 = TR_50 ;
	7'h6e :
		TR_227 = TR_50 ;
	7'h6f :
		TR_227 = TR_50 ;
	7'h70 :
		TR_227 = TR_50 ;
	7'h71 :
		TR_227 = TR_50 ;
	7'h72 :
		TR_227 = TR_50 ;
	7'h73 :
		TR_227 = TR_50 ;
	7'h74 :
		TR_227 = TR_50 ;
	7'h75 :
		TR_227 = TR_50 ;
	7'h76 :
		TR_227 = TR_50 ;
	7'h77 :
		TR_227 = TR_50 ;
	7'h78 :
		TR_227 = TR_50 ;
	7'h79 :
		TR_227 = TR_50 ;
	7'h7a :
		TR_227 = TR_50 ;
	7'h7b :
		TR_227 = TR_50 ;
	7'h7c :
		TR_227 = TR_50 ;
	7'h7d :
		TR_227 = TR_50 ;
	7'h7e :
		TR_227 = TR_50 ;
	7'h7f :
		TR_227 = TR_50 ;
	default :
		TR_227 = 9'hx ;
	endcase
always @ ( TR_227 or U_173 or sub8u_71ot or U_183 or RG_rl_148 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_38_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h26 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_38_t = ( ( { 9{ M_180 } } & RG_rl_148 )
		| ( { 9{ U_173 } } & TR_227 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_38_en = ( M_180 | RG_rl_38_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_38_en )
		RG_rl_38 <= RG_rl_38_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_51 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_226 = TR_51 ;
	7'h01 :
		TR_226 = TR_51 ;
	7'h02 :
		TR_226 = TR_51 ;
	7'h03 :
		TR_226 = TR_51 ;
	7'h04 :
		TR_226 = TR_51 ;
	7'h05 :
		TR_226 = TR_51 ;
	7'h06 :
		TR_226 = TR_51 ;
	7'h07 :
		TR_226 = TR_51 ;
	7'h08 :
		TR_226 = TR_51 ;
	7'h09 :
		TR_226 = TR_51 ;
	7'h0a :
		TR_226 = TR_51 ;
	7'h0b :
		TR_226 = TR_51 ;
	7'h0c :
		TR_226 = TR_51 ;
	7'h0d :
		TR_226 = TR_51 ;
	7'h0e :
		TR_226 = TR_51 ;
	7'h0f :
		TR_226 = TR_51 ;
	7'h10 :
		TR_226 = TR_51 ;
	7'h11 :
		TR_226 = TR_51 ;
	7'h12 :
		TR_226 = TR_51 ;
	7'h13 :
		TR_226 = TR_51 ;
	7'h14 :
		TR_226 = TR_51 ;
	7'h15 :
		TR_226 = TR_51 ;
	7'h16 :
		TR_226 = TR_51 ;
	7'h17 :
		TR_226 = TR_51 ;
	7'h18 :
		TR_226 = TR_51 ;
	7'h19 :
		TR_226 = TR_51 ;
	7'h1a :
		TR_226 = TR_51 ;
	7'h1b :
		TR_226 = TR_51 ;
	7'h1c :
		TR_226 = TR_51 ;
	7'h1d :
		TR_226 = TR_51 ;
	7'h1e :
		TR_226 = TR_51 ;
	7'h1f :
		TR_226 = TR_51 ;
	7'h20 :
		TR_226 = TR_51 ;
	7'h21 :
		TR_226 = TR_51 ;
	7'h22 :
		TR_226 = TR_51 ;
	7'h23 :
		TR_226 = TR_51 ;
	7'h24 :
		TR_226 = TR_51 ;
	7'h25 :
		TR_226 = TR_51 ;
	7'h26 :
		TR_226 = TR_51 ;
	7'h27 :
		TR_226 = 9'h000 ;	// line#=../rle.cpp:80
	7'h28 :
		TR_226 = TR_51 ;
	7'h29 :
		TR_226 = TR_51 ;
	7'h2a :
		TR_226 = TR_51 ;
	7'h2b :
		TR_226 = TR_51 ;
	7'h2c :
		TR_226 = TR_51 ;
	7'h2d :
		TR_226 = TR_51 ;
	7'h2e :
		TR_226 = TR_51 ;
	7'h2f :
		TR_226 = TR_51 ;
	7'h30 :
		TR_226 = TR_51 ;
	7'h31 :
		TR_226 = TR_51 ;
	7'h32 :
		TR_226 = TR_51 ;
	7'h33 :
		TR_226 = TR_51 ;
	7'h34 :
		TR_226 = TR_51 ;
	7'h35 :
		TR_226 = TR_51 ;
	7'h36 :
		TR_226 = TR_51 ;
	7'h37 :
		TR_226 = TR_51 ;
	7'h38 :
		TR_226 = TR_51 ;
	7'h39 :
		TR_226 = TR_51 ;
	7'h3a :
		TR_226 = TR_51 ;
	7'h3b :
		TR_226 = TR_51 ;
	7'h3c :
		TR_226 = TR_51 ;
	7'h3d :
		TR_226 = TR_51 ;
	7'h3e :
		TR_226 = TR_51 ;
	7'h3f :
		TR_226 = TR_51 ;
	7'h40 :
		TR_226 = TR_51 ;
	7'h41 :
		TR_226 = TR_51 ;
	7'h42 :
		TR_226 = TR_51 ;
	7'h43 :
		TR_226 = TR_51 ;
	7'h44 :
		TR_226 = TR_51 ;
	7'h45 :
		TR_226 = TR_51 ;
	7'h46 :
		TR_226 = TR_51 ;
	7'h47 :
		TR_226 = TR_51 ;
	7'h48 :
		TR_226 = TR_51 ;
	7'h49 :
		TR_226 = TR_51 ;
	7'h4a :
		TR_226 = TR_51 ;
	7'h4b :
		TR_226 = TR_51 ;
	7'h4c :
		TR_226 = TR_51 ;
	7'h4d :
		TR_226 = TR_51 ;
	7'h4e :
		TR_226 = TR_51 ;
	7'h4f :
		TR_226 = TR_51 ;
	7'h50 :
		TR_226 = TR_51 ;
	7'h51 :
		TR_226 = TR_51 ;
	7'h52 :
		TR_226 = TR_51 ;
	7'h53 :
		TR_226 = TR_51 ;
	7'h54 :
		TR_226 = TR_51 ;
	7'h55 :
		TR_226 = TR_51 ;
	7'h56 :
		TR_226 = TR_51 ;
	7'h57 :
		TR_226 = TR_51 ;
	7'h58 :
		TR_226 = TR_51 ;
	7'h59 :
		TR_226 = TR_51 ;
	7'h5a :
		TR_226 = TR_51 ;
	7'h5b :
		TR_226 = TR_51 ;
	7'h5c :
		TR_226 = TR_51 ;
	7'h5d :
		TR_226 = TR_51 ;
	7'h5e :
		TR_226 = TR_51 ;
	7'h5f :
		TR_226 = TR_51 ;
	7'h60 :
		TR_226 = TR_51 ;
	7'h61 :
		TR_226 = TR_51 ;
	7'h62 :
		TR_226 = TR_51 ;
	7'h63 :
		TR_226 = TR_51 ;
	7'h64 :
		TR_226 = TR_51 ;
	7'h65 :
		TR_226 = TR_51 ;
	7'h66 :
		TR_226 = TR_51 ;
	7'h67 :
		TR_226 = TR_51 ;
	7'h68 :
		TR_226 = TR_51 ;
	7'h69 :
		TR_226 = TR_51 ;
	7'h6a :
		TR_226 = TR_51 ;
	7'h6b :
		TR_226 = TR_51 ;
	7'h6c :
		TR_226 = TR_51 ;
	7'h6d :
		TR_226 = TR_51 ;
	7'h6e :
		TR_226 = TR_51 ;
	7'h6f :
		TR_226 = TR_51 ;
	7'h70 :
		TR_226 = TR_51 ;
	7'h71 :
		TR_226 = TR_51 ;
	7'h72 :
		TR_226 = TR_51 ;
	7'h73 :
		TR_226 = TR_51 ;
	7'h74 :
		TR_226 = TR_51 ;
	7'h75 :
		TR_226 = TR_51 ;
	7'h76 :
		TR_226 = TR_51 ;
	7'h77 :
		TR_226 = TR_51 ;
	7'h78 :
		TR_226 = TR_51 ;
	7'h79 :
		TR_226 = TR_51 ;
	7'h7a :
		TR_226 = TR_51 ;
	7'h7b :
		TR_226 = TR_51 ;
	7'h7c :
		TR_226 = TR_51 ;
	7'h7d :
		TR_226 = TR_51 ;
	7'h7e :
		TR_226 = TR_51 ;
	7'h7f :
		TR_226 = TR_51 ;
	default :
		TR_226 = 9'hx ;
	endcase
always @ ( TR_226 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_17 or 
	U_174 or RG_rl_148 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_39_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h27 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_39_t = ( ( { 9{ ST1_03d } } & RG_rl_148 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_17 )
		| ( { 9{ U_173 } } & TR_226 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_39_en = ( ST1_03d | U_174 | RG_rl_39_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_39_en )
		RG_rl_39 <= RG_rl_39_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_52 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_225 = TR_52 ;
	7'h01 :
		TR_225 = TR_52 ;
	7'h02 :
		TR_225 = TR_52 ;
	7'h03 :
		TR_225 = TR_52 ;
	7'h04 :
		TR_225 = TR_52 ;
	7'h05 :
		TR_225 = TR_52 ;
	7'h06 :
		TR_225 = TR_52 ;
	7'h07 :
		TR_225 = TR_52 ;
	7'h08 :
		TR_225 = TR_52 ;
	7'h09 :
		TR_225 = TR_52 ;
	7'h0a :
		TR_225 = TR_52 ;
	7'h0b :
		TR_225 = TR_52 ;
	7'h0c :
		TR_225 = TR_52 ;
	7'h0d :
		TR_225 = TR_52 ;
	7'h0e :
		TR_225 = TR_52 ;
	7'h0f :
		TR_225 = TR_52 ;
	7'h10 :
		TR_225 = TR_52 ;
	7'h11 :
		TR_225 = TR_52 ;
	7'h12 :
		TR_225 = TR_52 ;
	7'h13 :
		TR_225 = TR_52 ;
	7'h14 :
		TR_225 = TR_52 ;
	7'h15 :
		TR_225 = TR_52 ;
	7'h16 :
		TR_225 = TR_52 ;
	7'h17 :
		TR_225 = TR_52 ;
	7'h18 :
		TR_225 = TR_52 ;
	7'h19 :
		TR_225 = TR_52 ;
	7'h1a :
		TR_225 = TR_52 ;
	7'h1b :
		TR_225 = TR_52 ;
	7'h1c :
		TR_225 = TR_52 ;
	7'h1d :
		TR_225 = TR_52 ;
	7'h1e :
		TR_225 = TR_52 ;
	7'h1f :
		TR_225 = TR_52 ;
	7'h20 :
		TR_225 = TR_52 ;
	7'h21 :
		TR_225 = TR_52 ;
	7'h22 :
		TR_225 = TR_52 ;
	7'h23 :
		TR_225 = TR_52 ;
	7'h24 :
		TR_225 = TR_52 ;
	7'h25 :
		TR_225 = TR_52 ;
	7'h26 :
		TR_225 = TR_52 ;
	7'h27 :
		TR_225 = TR_52 ;
	7'h28 :
		TR_225 = 9'h000 ;	// line#=../rle.cpp:80
	7'h29 :
		TR_225 = TR_52 ;
	7'h2a :
		TR_225 = TR_52 ;
	7'h2b :
		TR_225 = TR_52 ;
	7'h2c :
		TR_225 = TR_52 ;
	7'h2d :
		TR_225 = TR_52 ;
	7'h2e :
		TR_225 = TR_52 ;
	7'h2f :
		TR_225 = TR_52 ;
	7'h30 :
		TR_225 = TR_52 ;
	7'h31 :
		TR_225 = TR_52 ;
	7'h32 :
		TR_225 = TR_52 ;
	7'h33 :
		TR_225 = TR_52 ;
	7'h34 :
		TR_225 = TR_52 ;
	7'h35 :
		TR_225 = TR_52 ;
	7'h36 :
		TR_225 = TR_52 ;
	7'h37 :
		TR_225 = TR_52 ;
	7'h38 :
		TR_225 = TR_52 ;
	7'h39 :
		TR_225 = TR_52 ;
	7'h3a :
		TR_225 = TR_52 ;
	7'h3b :
		TR_225 = TR_52 ;
	7'h3c :
		TR_225 = TR_52 ;
	7'h3d :
		TR_225 = TR_52 ;
	7'h3e :
		TR_225 = TR_52 ;
	7'h3f :
		TR_225 = TR_52 ;
	7'h40 :
		TR_225 = TR_52 ;
	7'h41 :
		TR_225 = TR_52 ;
	7'h42 :
		TR_225 = TR_52 ;
	7'h43 :
		TR_225 = TR_52 ;
	7'h44 :
		TR_225 = TR_52 ;
	7'h45 :
		TR_225 = TR_52 ;
	7'h46 :
		TR_225 = TR_52 ;
	7'h47 :
		TR_225 = TR_52 ;
	7'h48 :
		TR_225 = TR_52 ;
	7'h49 :
		TR_225 = TR_52 ;
	7'h4a :
		TR_225 = TR_52 ;
	7'h4b :
		TR_225 = TR_52 ;
	7'h4c :
		TR_225 = TR_52 ;
	7'h4d :
		TR_225 = TR_52 ;
	7'h4e :
		TR_225 = TR_52 ;
	7'h4f :
		TR_225 = TR_52 ;
	7'h50 :
		TR_225 = TR_52 ;
	7'h51 :
		TR_225 = TR_52 ;
	7'h52 :
		TR_225 = TR_52 ;
	7'h53 :
		TR_225 = TR_52 ;
	7'h54 :
		TR_225 = TR_52 ;
	7'h55 :
		TR_225 = TR_52 ;
	7'h56 :
		TR_225 = TR_52 ;
	7'h57 :
		TR_225 = TR_52 ;
	7'h58 :
		TR_225 = TR_52 ;
	7'h59 :
		TR_225 = TR_52 ;
	7'h5a :
		TR_225 = TR_52 ;
	7'h5b :
		TR_225 = TR_52 ;
	7'h5c :
		TR_225 = TR_52 ;
	7'h5d :
		TR_225 = TR_52 ;
	7'h5e :
		TR_225 = TR_52 ;
	7'h5f :
		TR_225 = TR_52 ;
	7'h60 :
		TR_225 = TR_52 ;
	7'h61 :
		TR_225 = TR_52 ;
	7'h62 :
		TR_225 = TR_52 ;
	7'h63 :
		TR_225 = TR_52 ;
	7'h64 :
		TR_225 = TR_52 ;
	7'h65 :
		TR_225 = TR_52 ;
	7'h66 :
		TR_225 = TR_52 ;
	7'h67 :
		TR_225 = TR_52 ;
	7'h68 :
		TR_225 = TR_52 ;
	7'h69 :
		TR_225 = TR_52 ;
	7'h6a :
		TR_225 = TR_52 ;
	7'h6b :
		TR_225 = TR_52 ;
	7'h6c :
		TR_225 = TR_52 ;
	7'h6d :
		TR_225 = TR_52 ;
	7'h6e :
		TR_225 = TR_52 ;
	7'h6f :
		TR_225 = TR_52 ;
	7'h70 :
		TR_225 = TR_52 ;
	7'h71 :
		TR_225 = TR_52 ;
	7'h72 :
		TR_225 = TR_52 ;
	7'h73 :
		TR_225 = TR_52 ;
	7'h74 :
		TR_225 = TR_52 ;
	7'h75 :
		TR_225 = TR_52 ;
	7'h76 :
		TR_225 = TR_52 ;
	7'h77 :
		TR_225 = TR_52 ;
	7'h78 :
		TR_225 = TR_52 ;
	7'h79 :
		TR_225 = TR_52 ;
	7'h7a :
		TR_225 = TR_52 ;
	7'h7b :
		TR_225 = TR_52 ;
	7'h7c :
		TR_225 = TR_52 ;
	7'h7d :
		TR_225 = TR_52 ;
	7'h7e :
		TR_225 = TR_52 ;
	7'h7f :
		TR_225 = TR_52 ;
	default :
		TR_225 = 9'hx ;
	endcase
always @ ( TR_225 or U_173 or sub8u_71ot or U_183 or RG_rl_149 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_40_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h28 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_40_t = ( ( { 9{ M_180 } } & RG_rl_149 )
		| ( { 9{ U_173 } } & TR_225 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_40_en = ( M_180 | RG_rl_40_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_40_en )
		RG_rl_40 <= RG_rl_40_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_53 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_224 = TR_53 ;
	7'h01 :
		TR_224 = TR_53 ;
	7'h02 :
		TR_224 = TR_53 ;
	7'h03 :
		TR_224 = TR_53 ;
	7'h04 :
		TR_224 = TR_53 ;
	7'h05 :
		TR_224 = TR_53 ;
	7'h06 :
		TR_224 = TR_53 ;
	7'h07 :
		TR_224 = TR_53 ;
	7'h08 :
		TR_224 = TR_53 ;
	7'h09 :
		TR_224 = TR_53 ;
	7'h0a :
		TR_224 = TR_53 ;
	7'h0b :
		TR_224 = TR_53 ;
	7'h0c :
		TR_224 = TR_53 ;
	7'h0d :
		TR_224 = TR_53 ;
	7'h0e :
		TR_224 = TR_53 ;
	7'h0f :
		TR_224 = TR_53 ;
	7'h10 :
		TR_224 = TR_53 ;
	7'h11 :
		TR_224 = TR_53 ;
	7'h12 :
		TR_224 = TR_53 ;
	7'h13 :
		TR_224 = TR_53 ;
	7'h14 :
		TR_224 = TR_53 ;
	7'h15 :
		TR_224 = TR_53 ;
	7'h16 :
		TR_224 = TR_53 ;
	7'h17 :
		TR_224 = TR_53 ;
	7'h18 :
		TR_224 = TR_53 ;
	7'h19 :
		TR_224 = TR_53 ;
	7'h1a :
		TR_224 = TR_53 ;
	7'h1b :
		TR_224 = TR_53 ;
	7'h1c :
		TR_224 = TR_53 ;
	7'h1d :
		TR_224 = TR_53 ;
	7'h1e :
		TR_224 = TR_53 ;
	7'h1f :
		TR_224 = TR_53 ;
	7'h20 :
		TR_224 = TR_53 ;
	7'h21 :
		TR_224 = TR_53 ;
	7'h22 :
		TR_224 = TR_53 ;
	7'h23 :
		TR_224 = TR_53 ;
	7'h24 :
		TR_224 = TR_53 ;
	7'h25 :
		TR_224 = TR_53 ;
	7'h26 :
		TR_224 = TR_53 ;
	7'h27 :
		TR_224 = TR_53 ;
	7'h28 :
		TR_224 = TR_53 ;
	7'h29 :
		TR_224 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2a :
		TR_224 = TR_53 ;
	7'h2b :
		TR_224 = TR_53 ;
	7'h2c :
		TR_224 = TR_53 ;
	7'h2d :
		TR_224 = TR_53 ;
	7'h2e :
		TR_224 = TR_53 ;
	7'h2f :
		TR_224 = TR_53 ;
	7'h30 :
		TR_224 = TR_53 ;
	7'h31 :
		TR_224 = TR_53 ;
	7'h32 :
		TR_224 = TR_53 ;
	7'h33 :
		TR_224 = TR_53 ;
	7'h34 :
		TR_224 = TR_53 ;
	7'h35 :
		TR_224 = TR_53 ;
	7'h36 :
		TR_224 = TR_53 ;
	7'h37 :
		TR_224 = TR_53 ;
	7'h38 :
		TR_224 = TR_53 ;
	7'h39 :
		TR_224 = TR_53 ;
	7'h3a :
		TR_224 = TR_53 ;
	7'h3b :
		TR_224 = TR_53 ;
	7'h3c :
		TR_224 = TR_53 ;
	7'h3d :
		TR_224 = TR_53 ;
	7'h3e :
		TR_224 = TR_53 ;
	7'h3f :
		TR_224 = TR_53 ;
	7'h40 :
		TR_224 = TR_53 ;
	7'h41 :
		TR_224 = TR_53 ;
	7'h42 :
		TR_224 = TR_53 ;
	7'h43 :
		TR_224 = TR_53 ;
	7'h44 :
		TR_224 = TR_53 ;
	7'h45 :
		TR_224 = TR_53 ;
	7'h46 :
		TR_224 = TR_53 ;
	7'h47 :
		TR_224 = TR_53 ;
	7'h48 :
		TR_224 = TR_53 ;
	7'h49 :
		TR_224 = TR_53 ;
	7'h4a :
		TR_224 = TR_53 ;
	7'h4b :
		TR_224 = TR_53 ;
	7'h4c :
		TR_224 = TR_53 ;
	7'h4d :
		TR_224 = TR_53 ;
	7'h4e :
		TR_224 = TR_53 ;
	7'h4f :
		TR_224 = TR_53 ;
	7'h50 :
		TR_224 = TR_53 ;
	7'h51 :
		TR_224 = TR_53 ;
	7'h52 :
		TR_224 = TR_53 ;
	7'h53 :
		TR_224 = TR_53 ;
	7'h54 :
		TR_224 = TR_53 ;
	7'h55 :
		TR_224 = TR_53 ;
	7'h56 :
		TR_224 = TR_53 ;
	7'h57 :
		TR_224 = TR_53 ;
	7'h58 :
		TR_224 = TR_53 ;
	7'h59 :
		TR_224 = TR_53 ;
	7'h5a :
		TR_224 = TR_53 ;
	7'h5b :
		TR_224 = TR_53 ;
	7'h5c :
		TR_224 = TR_53 ;
	7'h5d :
		TR_224 = TR_53 ;
	7'h5e :
		TR_224 = TR_53 ;
	7'h5f :
		TR_224 = TR_53 ;
	7'h60 :
		TR_224 = TR_53 ;
	7'h61 :
		TR_224 = TR_53 ;
	7'h62 :
		TR_224 = TR_53 ;
	7'h63 :
		TR_224 = TR_53 ;
	7'h64 :
		TR_224 = TR_53 ;
	7'h65 :
		TR_224 = TR_53 ;
	7'h66 :
		TR_224 = TR_53 ;
	7'h67 :
		TR_224 = TR_53 ;
	7'h68 :
		TR_224 = TR_53 ;
	7'h69 :
		TR_224 = TR_53 ;
	7'h6a :
		TR_224 = TR_53 ;
	7'h6b :
		TR_224 = TR_53 ;
	7'h6c :
		TR_224 = TR_53 ;
	7'h6d :
		TR_224 = TR_53 ;
	7'h6e :
		TR_224 = TR_53 ;
	7'h6f :
		TR_224 = TR_53 ;
	7'h70 :
		TR_224 = TR_53 ;
	7'h71 :
		TR_224 = TR_53 ;
	7'h72 :
		TR_224 = TR_53 ;
	7'h73 :
		TR_224 = TR_53 ;
	7'h74 :
		TR_224 = TR_53 ;
	7'h75 :
		TR_224 = TR_53 ;
	7'h76 :
		TR_224 = TR_53 ;
	7'h77 :
		TR_224 = TR_53 ;
	7'h78 :
		TR_224 = TR_53 ;
	7'h79 :
		TR_224 = TR_53 ;
	7'h7a :
		TR_224 = TR_53 ;
	7'h7b :
		TR_224 = TR_53 ;
	7'h7c :
		TR_224 = TR_53 ;
	7'h7d :
		TR_224 = TR_53 ;
	7'h7e :
		TR_224 = TR_53 ;
	7'h7f :
		TR_224 = TR_53 ;
	default :
		TR_224 = 9'hx ;
	endcase
always @ ( TR_224 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_18 or 
	U_174 or RG_rl_149 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_41_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h29 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_41_t = ( ( { 9{ ST1_03d } } & RG_rl_149 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_18 )
		| ( { 9{ U_173 } } & TR_224 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_41_en = ( ST1_03d | U_174 | RG_rl_41_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_41_en )
		RG_rl_41 <= RG_rl_41_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_54 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_223 = TR_54 ;
	7'h01 :
		TR_223 = TR_54 ;
	7'h02 :
		TR_223 = TR_54 ;
	7'h03 :
		TR_223 = TR_54 ;
	7'h04 :
		TR_223 = TR_54 ;
	7'h05 :
		TR_223 = TR_54 ;
	7'h06 :
		TR_223 = TR_54 ;
	7'h07 :
		TR_223 = TR_54 ;
	7'h08 :
		TR_223 = TR_54 ;
	7'h09 :
		TR_223 = TR_54 ;
	7'h0a :
		TR_223 = TR_54 ;
	7'h0b :
		TR_223 = TR_54 ;
	7'h0c :
		TR_223 = TR_54 ;
	7'h0d :
		TR_223 = TR_54 ;
	7'h0e :
		TR_223 = TR_54 ;
	7'h0f :
		TR_223 = TR_54 ;
	7'h10 :
		TR_223 = TR_54 ;
	7'h11 :
		TR_223 = TR_54 ;
	7'h12 :
		TR_223 = TR_54 ;
	7'h13 :
		TR_223 = TR_54 ;
	7'h14 :
		TR_223 = TR_54 ;
	7'h15 :
		TR_223 = TR_54 ;
	7'h16 :
		TR_223 = TR_54 ;
	7'h17 :
		TR_223 = TR_54 ;
	7'h18 :
		TR_223 = TR_54 ;
	7'h19 :
		TR_223 = TR_54 ;
	7'h1a :
		TR_223 = TR_54 ;
	7'h1b :
		TR_223 = TR_54 ;
	7'h1c :
		TR_223 = TR_54 ;
	7'h1d :
		TR_223 = TR_54 ;
	7'h1e :
		TR_223 = TR_54 ;
	7'h1f :
		TR_223 = TR_54 ;
	7'h20 :
		TR_223 = TR_54 ;
	7'h21 :
		TR_223 = TR_54 ;
	7'h22 :
		TR_223 = TR_54 ;
	7'h23 :
		TR_223 = TR_54 ;
	7'h24 :
		TR_223 = TR_54 ;
	7'h25 :
		TR_223 = TR_54 ;
	7'h26 :
		TR_223 = TR_54 ;
	7'h27 :
		TR_223 = TR_54 ;
	7'h28 :
		TR_223 = TR_54 ;
	7'h29 :
		TR_223 = TR_54 ;
	7'h2a :
		TR_223 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2b :
		TR_223 = TR_54 ;
	7'h2c :
		TR_223 = TR_54 ;
	7'h2d :
		TR_223 = TR_54 ;
	7'h2e :
		TR_223 = TR_54 ;
	7'h2f :
		TR_223 = TR_54 ;
	7'h30 :
		TR_223 = TR_54 ;
	7'h31 :
		TR_223 = TR_54 ;
	7'h32 :
		TR_223 = TR_54 ;
	7'h33 :
		TR_223 = TR_54 ;
	7'h34 :
		TR_223 = TR_54 ;
	7'h35 :
		TR_223 = TR_54 ;
	7'h36 :
		TR_223 = TR_54 ;
	7'h37 :
		TR_223 = TR_54 ;
	7'h38 :
		TR_223 = TR_54 ;
	7'h39 :
		TR_223 = TR_54 ;
	7'h3a :
		TR_223 = TR_54 ;
	7'h3b :
		TR_223 = TR_54 ;
	7'h3c :
		TR_223 = TR_54 ;
	7'h3d :
		TR_223 = TR_54 ;
	7'h3e :
		TR_223 = TR_54 ;
	7'h3f :
		TR_223 = TR_54 ;
	7'h40 :
		TR_223 = TR_54 ;
	7'h41 :
		TR_223 = TR_54 ;
	7'h42 :
		TR_223 = TR_54 ;
	7'h43 :
		TR_223 = TR_54 ;
	7'h44 :
		TR_223 = TR_54 ;
	7'h45 :
		TR_223 = TR_54 ;
	7'h46 :
		TR_223 = TR_54 ;
	7'h47 :
		TR_223 = TR_54 ;
	7'h48 :
		TR_223 = TR_54 ;
	7'h49 :
		TR_223 = TR_54 ;
	7'h4a :
		TR_223 = TR_54 ;
	7'h4b :
		TR_223 = TR_54 ;
	7'h4c :
		TR_223 = TR_54 ;
	7'h4d :
		TR_223 = TR_54 ;
	7'h4e :
		TR_223 = TR_54 ;
	7'h4f :
		TR_223 = TR_54 ;
	7'h50 :
		TR_223 = TR_54 ;
	7'h51 :
		TR_223 = TR_54 ;
	7'h52 :
		TR_223 = TR_54 ;
	7'h53 :
		TR_223 = TR_54 ;
	7'h54 :
		TR_223 = TR_54 ;
	7'h55 :
		TR_223 = TR_54 ;
	7'h56 :
		TR_223 = TR_54 ;
	7'h57 :
		TR_223 = TR_54 ;
	7'h58 :
		TR_223 = TR_54 ;
	7'h59 :
		TR_223 = TR_54 ;
	7'h5a :
		TR_223 = TR_54 ;
	7'h5b :
		TR_223 = TR_54 ;
	7'h5c :
		TR_223 = TR_54 ;
	7'h5d :
		TR_223 = TR_54 ;
	7'h5e :
		TR_223 = TR_54 ;
	7'h5f :
		TR_223 = TR_54 ;
	7'h60 :
		TR_223 = TR_54 ;
	7'h61 :
		TR_223 = TR_54 ;
	7'h62 :
		TR_223 = TR_54 ;
	7'h63 :
		TR_223 = TR_54 ;
	7'h64 :
		TR_223 = TR_54 ;
	7'h65 :
		TR_223 = TR_54 ;
	7'h66 :
		TR_223 = TR_54 ;
	7'h67 :
		TR_223 = TR_54 ;
	7'h68 :
		TR_223 = TR_54 ;
	7'h69 :
		TR_223 = TR_54 ;
	7'h6a :
		TR_223 = TR_54 ;
	7'h6b :
		TR_223 = TR_54 ;
	7'h6c :
		TR_223 = TR_54 ;
	7'h6d :
		TR_223 = TR_54 ;
	7'h6e :
		TR_223 = TR_54 ;
	7'h6f :
		TR_223 = TR_54 ;
	7'h70 :
		TR_223 = TR_54 ;
	7'h71 :
		TR_223 = TR_54 ;
	7'h72 :
		TR_223 = TR_54 ;
	7'h73 :
		TR_223 = TR_54 ;
	7'h74 :
		TR_223 = TR_54 ;
	7'h75 :
		TR_223 = TR_54 ;
	7'h76 :
		TR_223 = TR_54 ;
	7'h77 :
		TR_223 = TR_54 ;
	7'h78 :
		TR_223 = TR_54 ;
	7'h79 :
		TR_223 = TR_54 ;
	7'h7a :
		TR_223 = TR_54 ;
	7'h7b :
		TR_223 = TR_54 ;
	7'h7c :
		TR_223 = TR_54 ;
	7'h7d :
		TR_223 = TR_54 ;
	7'h7e :
		TR_223 = TR_54 ;
	7'h7f :
		TR_223 = TR_54 ;
	default :
		TR_223 = 9'hx ;
	endcase
always @ ( TR_223 or U_173 or sub8u_71ot or U_183 or RG_rl_150 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_42_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h2a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_42_t = ( ( { 9{ M_180 } } & RG_rl_150 )
		| ( { 9{ U_173 } } & TR_223 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_42_en = ( M_180 | RG_rl_42_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_42_en )
		RG_rl_42 <= RG_rl_42_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_55 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_222 = TR_55 ;
	7'h01 :
		TR_222 = TR_55 ;
	7'h02 :
		TR_222 = TR_55 ;
	7'h03 :
		TR_222 = TR_55 ;
	7'h04 :
		TR_222 = TR_55 ;
	7'h05 :
		TR_222 = TR_55 ;
	7'h06 :
		TR_222 = TR_55 ;
	7'h07 :
		TR_222 = TR_55 ;
	7'h08 :
		TR_222 = TR_55 ;
	7'h09 :
		TR_222 = TR_55 ;
	7'h0a :
		TR_222 = TR_55 ;
	7'h0b :
		TR_222 = TR_55 ;
	7'h0c :
		TR_222 = TR_55 ;
	7'h0d :
		TR_222 = TR_55 ;
	7'h0e :
		TR_222 = TR_55 ;
	7'h0f :
		TR_222 = TR_55 ;
	7'h10 :
		TR_222 = TR_55 ;
	7'h11 :
		TR_222 = TR_55 ;
	7'h12 :
		TR_222 = TR_55 ;
	7'h13 :
		TR_222 = TR_55 ;
	7'h14 :
		TR_222 = TR_55 ;
	7'h15 :
		TR_222 = TR_55 ;
	7'h16 :
		TR_222 = TR_55 ;
	7'h17 :
		TR_222 = TR_55 ;
	7'h18 :
		TR_222 = TR_55 ;
	7'h19 :
		TR_222 = TR_55 ;
	7'h1a :
		TR_222 = TR_55 ;
	7'h1b :
		TR_222 = TR_55 ;
	7'h1c :
		TR_222 = TR_55 ;
	7'h1d :
		TR_222 = TR_55 ;
	7'h1e :
		TR_222 = TR_55 ;
	7'h1f :
		TR_222 = TR_55 ;
	7'h20 :
		TR_222 = TR_55 ;
	7'h21 :
		TR_222 = TR_55 ;
	7'h22 :
		TR_222 = TR_55 ;
	7'h23 :
		TR_222 = TR_55 ;
	7'h24 :
		TR_222 = TR_55 ;
	7'h25 :
		TR_222 = TR_55 ;
	7'h26 :
		TR_222 = TR_55 ;
	7'h27 :
		TR_222 = TR_55 ;
	7'h28 :
		TR_222 = TR_55 ;
	7'h29 :
		TR_222 = TR_55 ;
	7'h2a :
		TR_222 = TR_55 ;
	7'h2b :
		TR_222 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2c :
		TR_222 = TR_55 ;
	7'h2d :
		TR_222 = TR_55 ;
	7'h2e :
		TR_222 = TR_55 ;
	7'h2f :
		TR_222 = TR_55 ;
	7'h30 :
		TR_222 = TR_55 ;
	7'h31 :
		TR_222 = TR_55 ;
	7'h32 :
		TR_222 = TR_55 ;
	7'h33 :
		TR_222 = TR_55 ;
	7'h34 :
		TR_222 = TR_55 ;
	7'h35 :
		TR_222 = TR_55 ;
	7'h36 :
		TR_222 = TR_55 ;
	7'h37 :
		TR_222 = TR_55 ;
	7'h38 :
		TR_222 = TR_55 ;
	7'h39 :
		TR_222 = TR_55 ;
	7'h3a :
		TR_222 = TR_55 ;
	7'h3b :
		TR_222 = TR_55 ;
	7'h3c :
		TR_222 = TR_55 ;
	7'h3d :
		TR_222 = TR_55 ;
	7'h3e :
		TR_222 = TR_55 ;
	7'h3f :
		TR_222 = TR_55 ;
	7'h40 :
		TR_222 = TR_55 ;
	7'h41 :
		TR_222 = TR_55 ;
	7'h42 :
		TR_222 = TR_55 ;
	7'h43 :
		TR_222 = TR_55 ;
	7'h44 :
		TR_222 = TR_55 ;
	7'h45 :
		TR_222 = TR_55 ;
	7'h46 :
		TR_222 = TR_55 ;
	7'h47 :
		TR_222 = TR_55 ;
	7'h48 :
		TR_222 = TR_55 ;
	7'h49 :
		TR_222 = TR_55 ;
	7'h4a :
		TR_222 = TR_55 ;
	7'h4b :
		TR_222 = TR_55 ;
	7'h4c :
		TR_222 = TR_55 ;
	7'h4d :
		TR_222 = TR_55 ;
	7'h4e :
		TR_222 = TR_55 ;
	7'h4f :
		TR_222 = TR_55 ;
	7'h50 :
		TR_222 = TR_55 ;
	7'h51 :
		TR_222 = TR_55 ;
	7'h52 :
		TR_222 = TR_55 ;
	7'h53 :
		TR_222 = TR_55 ;
	7'h54 :
		TR_222 = TR_55 ;
	7'h55 :
		TR_222 = TR_55 ;
	7'h56 :
		TR_222 = TR_55 ;
	7'h57 :
		TR_222 = TR_55 ;
	7'h58 :
		TR_222 = TR_55 ;
	7'h59 :
		TR_222 = TR_55 ;
	7'h5a :
		TR_222 = TR_55 ;
	7'h5b :
		TR_222 = TR_55 ;
	7'h5c :
		TR_222 = TR_55 ;
	7'h5d :
		TR_222 = TR_55 ;
	7'h5e :
		TR_222 = TR_55 ;
	7'h5f :
		TR_222 = TR_55 ;
	7'h60 :
		TR_222 = TR_55 ;
	7'h61 :
		TR_222 = TR_55 ;
	7'h62 :
		TR_222 = TR_55 ;
	7'h63 :
		TR_222 = TR_55 ;
	7'h64 :
		TR_222 = TR_55 ;
	7'h65 :
		TR_222 = TR_55 ;
	7'h66 :
		TR_222 = TR_55 ;
	7'h67 :
		TR_222 = TR_55 ;
	7'h68 :
		TR_222 = TR_55 ;
	7'h69 :
		TR_222 = TR_55 ;
	7'h6a :
		TR_222 = TR_55 ;
	7'h6b :
		TR_222 = TR_55 ;
	7'h6c :
		TR_222 = TR_55 ;
	7'h6d :
		TR_222 = TR_55 ;
	7'h6e :
		TR_222 = TR_55 ;
	7'h6f :
		TR_222 = TR_55 ;
	7'h70 :
		TR_222 = TR_55 ;
	7'h71 :
		TR_222 = TR_55 ;
	7'h72 :
		TR_222 = TR_55 ;
	7'h73 :
		TR_222 = TR_55 ;
	7'h74 :
		TR_222 = TR_55 ;
	7'h75 :
		TR_222 = TR_55 ;
	7'h76 :
		TR_222 = TR_55 ;
	7'h77 :
		TR_222 = TR_55 ;
	7'h78 :
		TR_222 = TR_55 ;
	7'h79 :
		TR_222 = TR_55 ;
	7'h7a :
		TR_222 = TR_55 ;
	7'h7b :
		TR_222 = TR_55 ;
	7'h7c :
		TR_222 = TR_55 ;
	7'h7d :
		TR_222 = TR_55 ;
	7'h7e :
		TR_222 = TR_55 ;
	7'h7f :
		TR_222 = TR_55 ;
	default :
		TR_222 = 9'hx ;
	endcase
always @ ( TR_222 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_19 or 
	U_174 or RG_rl_150 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_43_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h2b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_43_t = ( ( { 9{ ST1_03d } } & RG_rl_150 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_19 )
		| ( { 9{ U_173 } } & TR_222 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_43_en = ( ST1_03d | U_174 | RG_rl_43_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_43_en )
		RG_rl_43 <= RG_rl_43_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_56 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_221 = TR_56 ;
	7'h01 :
		TR_221 = TR_56 ;
	7'h02 :
		TR_221 = TR_56 ;
	7'h03 :
		TR_221 = TR_56 ;
	7'h04 :
		TR_221 = TR_56 ;
	7'h05 :
		TR_221 = TR_56 ;
	7'h06 :
		TR_221 = TR_56 ;
	7'h07 :
		TR_221 = TR_56 ;
	7'h08 :
		TR_221 = TR_56 ;
	7'h09 :
		TR_221 = TR_56 ;
	7'h0a :
		TR_221 = TR_56 ;
	7'h0b :
		TR_221 = TR_56 ;
	7'h0c :
		TR_221 = TR_56 ;
	7'h0d :
		TR_221 = TR_56 ;
	7'h0e :
		TR_221 = TR_56 ;
	7'h0f :
		TR_221 = TR_56 ;
	7'h10 :
		TR_221 = TR_56 ;
	7'h11 :
		TR_221 = TR_56 ;
	7'h12 :
		TR_221 = TR_56 ;
	7'h13 :
		TR_221 = TR_56 ;
	7'h14 :
		TR_221 = TR_56 ;
	7'h15 :
		TR_221 = TR_56 ;
	7'h16 :
		TR_221 = TR_56 ;
	7'h17 :
		TR_221 = TR_56 ;
	7'h18 :
		TR_221 = TR_56 ;
	7'h19 :
		TR_221 = TR_56 ;
	7'h1a :
		TR_221 = TR_56 ;
	7'h1b :
		TR_221 = TR_56 ;
	7'h1c :
		TR_221 = TR_56 ;
	7'h1d :
		TR_221 = TR_56 ;
	7'h1e :
		TR_221 = TR_56 ;
	7'h1f :
		TR_221 = TR_56 ;
	7'h20 :
		TR_221 = TR_56 ;
	7'h21 :
		TR_221 = TR_56 ;
	7'h22 :
		TR_221 = TR_56 ;
	7'h23 :
		TR_221 = TR_56 ;
	7'h24 :
		TR_221 = TR_56 ;
	7'h25 :
		TR_221 = TR_56 ;
	7'h26 :
		TR_221 = TR_56 ;
	7'h27 :
		TR_221 = TR_56 ;
	7'h28 :
		TR_221 = TR_56 ;
	7'h29 :
		TR_221 = TR_56 ;
	7'h2a :
		TR_221 = TR_56 ;
	7'h2b :
		TR_221 = TR_56 ;
	7'h2c :
		TR_221 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2d :
		TR_221 = TR_56 ;
	7'h2e :
		TR_221 = TR_56 ;
	7'h2f :
		TR_221 = TR_56 ;
	7'h30 :
		TR_221 = TR_56 ;
	7'h31 :
		TR_221 = TR_56 ;
	7'h32 :
		TR_221 = TR_56 ;
	7'h33 :
		TR_221 = TR_56 ;
	7'h34 :
		TR_221 = TR_56 ;
	7'h35 :
		TR_221 = TR_56 ;
	7'h36 :
		TR_221 = TR_56 ;
	7'h37 :
		TR_221 = TR_56 ;
	7'h38 :
		TR_221 = TR_56 ;
	7'h39 :
		TR_221 = TR_56 ;
	7'h3a :
		TR_221 = TR_56 ;
	7'h3b :
		TR_221 = TR_56 ;
	7'h3c :
		TR_221 = TR_56 ;
	7'h3d :
		TR_221 = TR_56 ;
	7'h3e :
		TR_221 = TR_56 ;
	7'h3f :
		TR_221 = TR_56 ;
	7'h40 :
		TR_221 = TR_56 ;
	7'h41 :
		TR_221 = TR_56 ;
	7'h42 :
		TR_221 = TR_56 ;
	7'h43 :
		TR_221 = TR_56 ;
	7'h44 :
		TR_221 = TR_56 ;
	7'h45 :
		TR_221 = TR_56 ;
	7'h46 :
		TR_221 = TR_56 ;
	7'h47 :
		TR_221 = TR_56 ;
	7'h48 :
		TR_221 = TR_56 ;
	7'h49 :
		TR_221 = TR_56 ;
	7'h4a :
		TR_221 = TR_56 ;
	7'h4b :
		TR_221 = TR_56 ;
	7'h4c :
		TR_221 = TR_56 ;
	7'h4d :
		TR_221 = TR_56 ;
	7'h4e :
		TR_221 = TR_56 ;
	7'h4f :
		TR_221 = TR_56 ;
	7'h50 :
		TR_221 = TR_56 ;
	7'h51 :
		TR_221 = TR_56 ;
	7'h52 :
		TR_221 = TR_56 ;
	7'h53 :
		TR_221 = TR_56 ;
	7'h54 :
		TR_221 = TR_56 ;
	7'h55 :
		TR_221 = TR_56 ;
	7'h56 :
		TR_221 = TR_56 ;
	7'h57 :
		TR_221 = TR_56 ;
	7'h58 :
		TR_221 = TR_56 ;
	7'h59 :
		TR_221 = TR_56 ;
	7'h5a :
		TR_221 = TR_56 ;
	7'h5b :
		TR_221 = TR_56 ;
	7'h5c :
		TR_221 = TR_56 ;
	7'h5d :
		TR_221 = TR_56 ;
	7'h5e :
		TR_221 = TR_56 ;
	7'h5f :
		TR_221 = TR_56 ;
	7'h60 :
		TR_221 = TR_56 ;
	7'h61 :
		TR_221 = TR_56 ;
	7'h62 :
		TR_221 = TR_56 ;
	7'h63 :
		TR_221 = TR_56 ;
	7'h64 :
		TR_221 = TR_56 ;
	7'h65 :
		TR_221 = TR_56 ;
	7'h66 :
		TR_221 = TR_56 ;
	7'h67 :
		TR_221 = TR_56 ;
	7'h68 :
		TR_221 = TR_56 ;
	7'h69 :
		TR_221 = TR_56 ;
	7'h6a :
		TR_221 = TR_56 ;
	7'h6b :
		TR_221 = TR_56 ;
	7'h6c :
		TR_221 = TR_56 ;
	7'h6d :
		TR_221 = TR_56 ;
	7'h6e :
		TR_221 = TR_56 ;
	7'h6f :
		TR_221 = TR_56 ;
	7'h70 :
		TR_221 = TR_56 ;
	7'h71 :
		TR_221 = TR_56 ;
	7'h72 :
		TR_221 = TR_56 ;
	7'h73 :
		TR_221 = TR_56 ;
	7'h74 :
		TR_221 = TR_56 ;
	7'h75 :
		TR_221 = TR_56 ;
	7'h76 :
		TR_221 = TR_56 ;
	7'h77 :
		TR_221 = TR_56 ;
	7'h78 :
		TR_221 = TR_56 ;
	7'h79 :
		TR_221 = TR_56 ;
	7'h7a :
		TR_221 = TR_56 ;
	7'h7b :
		TR_221 = TR_56 ;
	7'h7c :
		TR_221 = TR_56 ;
	7'h7d :
		TR_221 = TR_56 ;
	7'h7e :
		TR_221 = TR_56 ;
	7'h7f :
		TR_221 = TR_56 ;
	default :
		TR_221 = 9'hx ;
	endcase
always @ ( TR_221 or U_173 or sub8u_71ot or U_183 or RG_rl_151 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_44_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h2c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_44_t = ( ( { 9{ M_180 } } & RG_rl_151 )
		| ( { 9{ U_173 } } & TR_221 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_44_en = ( M_180 | RG_rl_44_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_44_en )
		RG_rl_44 <= RG_rl_44_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_57 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_220 = TR_57 ;
	7'h01 :
		TR_220 = TR_57 ;
	7'h02 :
		TR_220 = TR_57 ;
	7'h03 :
		TR_220 = TR_57 ;
	7'h04 :
		TR_220 = TR_57 ;
	7'h05 :
		TR_220 = TR_57 ;
	7'h06 :
		TR_220 = TR_57 ;
	7'h07 :
		TR_220 = TR_57 ;
	7'h08 :
		TR_220 = TR_57 ;
	7'h09 :
		TR_220 = TR_57 ;
	7'h0a :
		TR_220 = TR_57 ;
	7'h0b :
		TR_220 = TR_57 ;
	7'h0c :
		TR_220 = TR_57 ;
	7'h0d :
		TR_220 = TR_57 ;
	7'h0e :
		TR_220 = TR_57 ;
	7'h0f :
		TR_220 = TR_57 ;
	7'h10 :
		TR_220 = TR_57 ;
	7'h11 :
		TR_220 = TR_57 ;
	7'h12 :
		TR_220 = TR_57 ;
	7'h13 :
		TR_220 = TR_57 ;
	7'h14 :
		TR_220 = TR_57 ;
	7'h15 :
		TR_220 = TR_57 ;
	7'h16 :
		TR_220 = TR_57 ;
	7'h17 :
		TR_220 = TR_57 ;
	7'h18 :
		TR_220 = TR_57 ;
	7'h19 :
		TR_220 = TR_57 ;
	7'h1a :
		TR_220 = TR_57 ;
	7'h1b :
		TR_220 = TR_57 ;
	7'h1c :
		TR_220 = TR_57 ;
	7'h1d :
		TR_220 = TR_57 ;
	7'h1e :
		TR_220 = TR_57 ;
	7'h1f :
		TR_220 = TR_57 ;
	7'h20 :
		TR_220 = TR_57 ;
	7'h21 :
		TR_220 = TR_57 ;
	7'h22 :
		TR_220 = TR_57 ;
	7'h23 :
		TR_220 = TR_57 ;
	7'h24 :
		TR_220 = TR_57 ;
	7'h25 :
		TR_220 = TR_57 ;
	7'h26 :
		TR_220 = TR_57 ;
	7'h27 :
		TR_220 = TR_57 ;
	7'h28 :
		TR_220 = TR_57 ;
	7'h29 :
		TR_220 = TR_57 ;
	7'h2a :
		TR_220 = TR_57 ;
	7'h2b :
		TR_220 = TR_57 ;
	7'h2c :
		TR_220 = TR_57 ;
	7'h2d :
		TR_220 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2e :
		TR_220 = TR_57 ;
	7'h2f :
		TR_220 = TR_57 ;
	7'h30 :
		TR_220 = TR_57 ;
	7'h31 :
		TR_220 = TR_57 ;
	7'h32 :
		TR_220 = TR_57 ;
	7'h33 :
		TR_220 = TR_57 ;
	7'h34 :
		TR_220 = TR_57 ;
	7'h35 :
		TR_220 = TR_57 ;
	7'h36 :
		TR_220 = TR_57 ;
	7'h37 :
		TR_220 = TR_57 ;
	7'h38 :
		TR_220 = TR_57 ;
	7'h39 :
		TR_220 = TR_57 ;
	7'h3a :
		TR_220 = TR_57 ;
	7'h3b :
		TR_220 = TR_57 ;
	7'h3c :
		TR_220 = TR_57 ;
	7'h3d :
		TR_220 = TR_57 ;
	7'h3e :
		TR_220 = TR_57 ;
	7'h3f :
		TR_220 = TR_57 ;
	7'h40 :
		TR_220 = TR_57 ;
	7'h41 :
		TR_220 = TR_57 ;
	7'h42 :
		TR_220 = TR_57 ;
	7'h43 :
		TR_220 = TR_57 ;
	7'h44 :
		TR_220 = TR_57 ;
	7'h45 :
		TR_220 = TR_57 ;
	7'h46 :
		TR_220 = TR_57 ;
	7'h47 :
		TR_220 = TR_57 ;
	7'h48 :
		TR_220 = TR_57 ;
	7'h49 :
		TR_220 = TR_57 ;
	7'h4a :
		TR_220 = TR_57 ;
	7'h4b :
		TR_220 = TR_57 ;
	7'h4c :
		TR_220 = TR_57 ;
	7'h4d :
		TR_220 = TR_57 ;
	7'h4e :
		TR_220 = TR_57 ;
	7'h4f :
		TR_220 = TR_57 ;
	7'h50 :
		TR_220 = TR_57 ;
	7'h51 :
		TR_220 = TR_57 ;
	7'h52 :
		TR_220 = TR_57 ;
	7'h53 :
		TR_220 = TR_57 ;
	7'h54 :
		TR_220 = TR_57 ;
	7'h55 :
		TR_220 = TR_57 ;
	7'h56 :
		TR_220 = TR_57 ;
	7'h57 :
		TR_220 = TR_57 ;
	7'h58 :
		TR_220 = TR_57 ;
	7'h59 :
		TR_220 = TR_57 ;
	7'h5a :
		TR_220 = TR_57 ;
	7'h5b :
		TR_220 = TR_57 ;
	7'h5c :
		TR_220 = TR_57 ;
	7'h5d :
		TR_220 = TR_57 ;
	7'h5e :
		TR_220 = TR_57 ;
	7'h5f :
		TR_220 = TR_57 ;
	7'h60 :
		TR_220 = TR_57 ;
	7'h61 :
		TR_220 = TR_57 ;
	7'h62 :
		TR_220 = TR_57 ;
	7'h63 :
		TR_220 = TR_57 ;
	7'h64 :
		TR_220 = TR_57 ;
	7'h65 :
		TR_220 = TR_57 ;
	7'h66 :
		TR_220 = TR_57 ;
	7'h67 :
		TR_220 = TR_57 ;
	7'h68 :
		TR_220 = TR_57 ;
	7'h69 :
		TR_220 = TR_57 ;
	7'h6a :
		TR_220 = TR_57 ;
	7'h6b :
		TR_220 = TR_57 ;
	7'h6c :
		TR_220 = TR_57 ;
	7'h6d :
		TR_220 = TR_57 ;
	7'h6e :
		TR_220 = TR_57 ;
	7'h6f :
		TR_220 = TR_57 ;
	7'h70 :
		TR_220 = TR_57 ;
	7'h71 :
		TR_220 = TR_57 ;
	7'h72 :
		TR_220 = TR_57 ;
	7'h73 :
		TR_220 = TR_57 ;
	7'h74 :
		TR_220 = TR_57 ;
	7'h75 :
		TR_220 = TR_57 ;
	7'h76 :
		TR_220 = TR_57 ;
	7'h77 :
		TR_220 = TR_57 ;
	7'h78 :
		TR_220 = TR_57 ;
	7'h79 :
		TR_220 = TR_57 ;
	7'h7a :
		TR_220 = TR_57 ;
	7'h7b :
		TR_220 = TR_57 ;
	7'h7c :
		TR_220 = TR_57 ;
	7'h7d :
		TR_220 = TR_57 ;
	7'h7e :
		TR_220 = TR_57 ;
	7'h7f :
		TR_220 = TR_57 ;
	default :
		TR_220 = 9'hx ;
	endcase
always @ ( TR_220 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_20 or 
	U_174 or RG_rl_151 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_45_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h2d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_45_t = ( ( { 9{ ST1_03d } } & RG_rl_151 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_20 )
		| ( { 9{ U_173 } } & TR_220 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_45_en = ( ST1_03d | U_174 | RG_rl_45_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_45_en )
		RG_rl_45 <= RG_rl_45_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_58 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_219 = TR_58 ;
	7'h01 :
		TR_219 = TR_58 ;
	7'h02 :
		TR_219 = TR_58 ;
	7'h03 :
		TR_219 = TR_58 ;
	7'h04 :
		TR_219 = TR_58 ;
	7'h05 :
		TR_219 = TR_58 ;
	7'h06 :
		TR_219 = TR_58 ;
	7'h07 :
		TR_219 = TR_58 ;
	7'h08 :
		TR_219 = TR_58 ;
	7'h09 :
		TR_219 = TR_58 ;
	7'h0a :
		TR_219 = TR_58 ;
	7'h0b :
		TR_219 = TR_58 ;
	7'h0c :
		TR_219 = TR_58 ;
	7'h0d :
		TR_219 = TR_58 ;
	7'h0e :
		TR_219 = TR_58 ;
	7'h0f :
		TR_219 = TR_58 ;
	7'h10 :
		TR_219 = TR_58 ;
	7'h11 :
		TR_219 = TR_58 ;
	7'h12 :
		TR_219 = TR_58 ;
	7'h13 :
		TR_219 = TR_58 ;
	7'h14 :
		TR_219 = TR_58 ;
	7'h15 :
		TR_219 = TR_58 ;
	7'h16 :
		TR_219 = TR_58 ;
	7'h17 :
		TR_219 = TR_58 ;
	7'h18 :
		TR_219 = TR_58 ;
	7'h19 :
		TR_219 = TR_58 ;
	7'h1a :
		TR_219 = TR_58 ;
	7'h1b :
		TR_219 = TR_58 ;
	7'h1c :
		TR_219 = TR_58 ;
	7'h1d :
		TR_219 = TR_58 ;
	7'h1e :
		TR_219 = TR_58 ;
	7'h1f :
		TR_219 = TR_58 ;
	7'h20 :
		TR_219 = TR_58 ;
	7'h21 :
		TR_219 = TR_58 ;
	7'h22 :
		TR_219 = TR_58 ;
	7'h23 :
		TR_219 = TR_58 ;
	7'h24 :
		TR_219 = TR_58 ;
	7'h25 :
		TR_219 = TR_58 ;
	7'h26 :
		TR_219 = TR_58 ;
	7'h27 :
		TR_219 = TR_58 ;
	7'h28 :
		TR_219 = TR_58 ;
	7'h29 :
		TR_219 = TR_58 ;
	7'h2a :
		TR_219 = TR_58 ;
	7'h2b :
		TR_219 = TR_58 ;
	7'h2c :
		TR_219 = TR_58 ;
	7'h2d :
		TR_219 = TR_58 ;
	7'h2e :
		TR_219 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2f :
		TR_219 = TR_58 ;
	7'h30 :
		TR_219 = TR_58 ;
	7'h31 :
		TR_219 = TR_58 ;
	7'h32 :
		TR_219 = TR_58 ;
	7'h33 :
		TR_219 = TR_58 ;
	7'h34 :
		TR_219 = TR_58 ;
	7'h35 :
		TR_219 = TR_58 ;
	7'h36 :
		TR_219 = TR_58 ;
	7'h37 :
		TR_219 = TR_58 ;
	7'h38 :
		TR_219 = TR_58 ;
	7'h39 :
		TR_219 = TR_58 ;
	7'h3a :
		TR_219 = TR_58 ;
	7'h3b :
		TR_219 = TR_58 ;
	7'h3c :
		TR_219 = TR_58 ;
	7'h3d :
		TR_219 = TR_58 ;
	7'h3e :
		TR_219 = TR_58 ;
	7'h3f :
		TR_219 = TR_58 ;
	7'h40 :
		TR_219 = TR_58 ;
	7'h41 :
		TR_219 = TR_58 ;
	7'h42 :
		TR_219 = TR_58 ;
	7'h43 :
		TR_219 = TR_58 ;
	7'h44 :
		TR_219 = TR_58 ;
	7'h45 :
		TR_219 = TR_58 ;
	7'h46 :
		TR_219 = TR_58 ;
	7'h47 :
		TR_219 = TR_58 ;
	7'h48 :
		TR_219 = TR_58 ;
	7'h49 :
		TR_219 = TR_58 ;
	7'h4a :
		TR_219 = TR_58 ;
	7'h4b :
		TR_219 = TR_58 ;
	7'h4c :
		TR_219 = TR_58 ;
	7'h4d :
		TR_219 = TR_58 ;
	7'h4e :
		TR_219 = TR_58 ;
	7'h4f :
		TR_219 = TR_58 ;
	7'h50 :
		TR_219 = TR_58 ;
	7'h51 :
		TR_219 = TR_58 ;
	7'h52 :
		TR_219 = TR_58 ;
	7'h53 :
		TR_219 = TR_58 ;
	7'h54 :
		TR_219 = TR_58 ;
	7'h55 :
		TR_219 = TR_58 ;
	7'h56 :
		TR_219 = TR_58 ;
	7'h57 :
		TR_219 = TR_58 ;
	7'h58 :
		TR_219 = TR_58 ;
	7'h59 :
		TR_219 = TR_58 ;
	7'h5a :
		TR_219 = TR_58 ;
	7'h5b :
		TR_219 = TR_58 ;
	7'h5c :
		TR_219 = TR_58 ;
	7'h5d :
		TR_219 = TR_58 ;
	7'h5e :
		TR_219 = TR_58 ;
	7'h5f :
		TR_219 = TR_58 ;
	7'h60 :
		TR_219 = TR_58 ;
	7'h61 :
		TR_219 = TR_58 ;
	7'h62 :
		TR_219 = TR_58 ;
	7'h63 :
		TR_219 = TR_58 ;
	7'h64 :
		TR_219 = TR_58 ;
	7'h65 :
		TR_219 = TR_58 ;
	7'h66 :
		TR_219 = TR_58 ;
	7'h67 :
		TR_219 = TR_58 ;
	7'h68 :
		TR_219 = TR_58 ;
	7'h69 :
		TR_219 = TR_58 ;
	7'h6a :
		TR_219 = TR_58 ;
	7'h6b :
		TR_219 = TR_58 ;
	7'h6c :
		TR_219 = TR_58 ;
	7'h6d :
		TR_219 = TR_58 ;
	7'h6e :
		TR_219 = TR_58 ;
	7'h6f :
		TR_219 = TR_58 ;
	7'h70 :
		TR_219 = TR_58 ;
	7'h71 :
		TR_219 = TR_58 ;
	7'h72 :
		TR_219 = TR_58 ;
	7'h73 :
		TR_219 = TR_58 ;
	7'h74 :
		TR_219 = TR_58 ;
	7'h75 :
		TR_219 = TR_58 ;
	7'h76 :
		TR_219 = TR_58 ;
	7'h77 :
		TR_219 = TR_58 ;
	7'h78 :
		TR_219 = TR_58 ;
	7'h79 :
		TR_219 = TR_58 ;
	7'h7a :
		TR_219 = TR_58 ;
	7'h7b :
		TR_219 = TR_58 ;
	7'h7c :
		TR_219 = TR_58 ;
	7'h7d :
		TR_219 = TR_58 ;
	7'h7e :
		TR_219 = TR_58 ;
	7'h7f :
		TR_219 = TR_58 ;
	default :
		TR_219 = 9'hx ;
	endcase
always @ ( TR_219 or U_173 or sub8u_71ot or U_183 or RG_rl_152 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_46_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h2e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_46_t = ( ( { 9{ M_180 } } & RG_rl_152 )
		| ( { 9{ U_173 } } & TR_219 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_46_en = ( M_180 | RG_rl_46_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_46_en )
		RG_rl_46 <= RG_rl_46_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_59 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_218 = TR_59 ;
	7'h01 :
		TR_218 = TR_59 ;
	7'h02 :
		TR_218 = TR_59 ;
	7'h03 :
		TR_218 = TR_59 ;
	7'h04 :
		TR_218 = TR_59 ;
	7'h05 :
		TR_218 = TR_59 ;
	7'h06 :
		TR_218 = TR_59 ;
	7'h07 :
		TR_218 = TR_59 ;
	7'h08 :
		TR_218 = TR_59 ;
	7'h09 :
		TR_218 = TR_59 ;
	7'h0a :
		TR_218 = TR_59 ;
	7'h0b :
		TR_218 = TR_59 ;
	7'h0c :
		TR_218 = TR_59 ;
	7'h0d :
		TR_218 = TR_59 ;
	7'h0e :
		TR_218 = TR_59 ;
	7'h0f :
		TR_218 = TR_59 ;
	7'h10 :
		TR_218 = TR_59 ;
	7'h11 :
		TR_218 = TR_59 ;
	7'h12 :
		TR_218 = TR_59 ;
	7'h13 :
		TR_218 = TR_59 ;
	7'h14 :
		TR_218 = TR_59 ;
	7'h15 :
		TR_218 = TR_59 ;
	7'h16 :
		TR_218 = TR_59 ;
	7'h17 :
		TR_218 = TR_59 ;
	7'h18 :
		TR_218 = TR_59 ;
	7'h19 :
		TR_218 = TR_59 ;
	7'h1a :
		TR_218 = TR_59 ;
	7'h1b :
		TR_218 = TR_59 ;
	7'h1c :
		TR_218 = TR_59 ;
	7'h1d :
		TR_218 = TR_59 ;
	7'h1e :
		TR_218 = TR_59 ;
	7'h1f :
		TR_218 = TR_59 ;
	7'h20 :
		TR_218 = TR_59 ;
	7'h21 :
		TR_218 = TR_59 ;
	7'h22 :
		TR_218 = TR_59 ;
	7'h23 :
		TR_218 = TR_59 ;
	7'h24 :
		TR_218 = TR_59 ;
	7'h25 :
		TR_218 = TR_59 ;
	7'h26 :
		TR_218 = TR_59 ;
	7'h27 :
		TR_218 = TR_59 ;
	7'h28 :
		TR_218 = TR_59 ;
	7'h29 :
		TR_218 = TR_59 ;
	7'h2a :
		TR_218 = TR_59 ;
	7'h2b :
		TR_218 = TR_59 ;
	7'h2c :
		TR_218 = TR_59 ;
	7'h2d :
		TR_218 = TR_59 ;
	7'h2e :
		TR_218 = TR_59 ;
	7'h2f :
		TR_218 = 9'h000 ;	// line#=../rle.cpp:80
	7'h30 :
		TR_218 = TR_59 ;
	7'h31 :
		TR_218 = TR_59 ;
	7'h32 :
		TR_218 = TR_59 ;
	7'h33 :
		TR_218 = TR_59 ;
	7'h34 :
		TR_218 = TR_59 ;
	7'h35 :
		TR_218 = TR_59 ;
	7'h36 :
		TR_218 = TR_59 ;
	7'h37 :
		TR_218 = TR_59 ;
	7'h38 :
		TR_218 = TR_59 ;
	7'h39 :
		TR_218 = TR_59 ;
	7'h3a :
		TR_218 = TR_59 ;
	7'h3b :
		TR_218 = TR_59 ;
	7'h3c :
		TR_218 = TR_59 ;
	7'h3d :
		TR_218 = TR_59 ;
	7'h3e :
		TR_218 = TR_59 ;
	7'h3f :
		TR_218 = TR_59 ;
	7'h40 :
		TR_218 = TR_59 ;
	7'h41 :
		TR_218 = TR_59 ;
	7'h42 :
		TR_218 = TR_59 ;
	7'h43 :
		TR_218 = TR_59 ;
	7'h44 :
		TR_218 = TR_59 ;
	7'h45 :
		TR_218 = TR_59 ;
	7'h46 :
		TR_218 = TR_59 ;
	7'h47 :
		TR_218 = TR_59 ;
	7'h48 :
		TR_218 = TR_59 ;
	7'h49 :
		TR_218 = TR_59 ;
	7'h4a :
		TR_218 = TR_59 ;
	7'h4b :
		TR_218 = TR_59 ;
	7'h4c :
		TR_218 = TR_59 ;
	7'h4d :
		TR_218 = TR_59 ;
	7'h4e :
		TR_218 = TR_59 ;
	7'h4f :
		TR_218 = TR_59 ;
	7'h50 :
		TR_218 = TR_59 ;
	7'h51 :
		TR_218 = TR_59 ;
	7'h52 :
		TR_218 = TR_59 ;
	7'h53 :
		TR_218 = TR_59 ;
	7'h54 :
		TR_218 = TR_59 ;
	7'h55 :
		TR_218 = TR_59 ;
	7'h56 :
		TR_218 = TR_59 ;
	7'h57 :
		TR_218 = TR_59 ;
	7'h58 :
		TR_218 = TR_59 ;
	7'h59 :
		TR_218 = TR_59 ;
	7'h5a :
		TR_218 = TR_59 ;
	7'h5b :
		TR_218 = TR_59 ;
	7'h5c :
		TR_218 = TR_59 ;
	7'h5d :
		TR_218 = TR_59 ;
	7'h5e :
		TR_218 = TR_59 ;
	7'h5f :
		TR_218 = TR_59 ;
	7'h60 :
		TR_218 = TR_59 ;
	7'h61 :
		TR_218 = TR_59 ;
	7'h62 :
		TR_218 = TR_59 ;
	7'h63 :
		TR_218 = TR_59 ;
	7'h64 :
		TR_218 = TR_59 ;
	7'h65 :
		TR_218 = TR_59 ;
	7'h66 :
		TR_218 = TR_59 ;
	7'h67 :
		TR_218 = TR_59 ;
	7'h68 :
		TR_218 = TR_59 ;
	7'h69 :
		TR_218 = TR_59 ;
	7'h6a :
		TR_218 = TR_59 ;
	7'h6b :
		TR_218 = TR_59 ;
	7'h6c :
		TR_218 = TR_59 ;
	7'h6d :
		TR_218 = TR_59 ;
	7'h6e :
		TR_218 = TR_59 ;
	7'h6f :
		TR_218 = TR_59 ;
	7'h70 :
		TR_218 = TR_59 ;
	7'h71 :
		TR_218 = TR_59 ;
	7'h72 :
		TR_218 = TR_59 ;
	7'h73 :
		TR_218 = TR_59 ;
	7'h74 :
		TR_218 = TR_59 ;
	7'h75 :
		TR_218 = TR_59 ;
	7'h76 :
		TR_218 = TR_59 ;
	7'h77 :
		TR_218 = TR_59 ;
	7'h78 :
		TR_218 = TR_59 ;
	7'h79 :
		TR_218 = TR_59 ;
	7'h7a :
		TR_218 = TR_59 ;
	7'h7b :
		TR_218 = TR_59 ;
	7'h7c :
		TR_218 = TR_59 ;
	7'h7d :
		TR_218 = TR_59 ;
	7'h7e :
		TR_218 = TR_59 ;
	7'h7f :
		TR_218 = TR_59 ;
	default :
		TR_218 = 9'hx ;
	endcase
always @ ( TR_218 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_21 or 
	U_174 or RG_rl_152 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_47_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h2f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_47_t = ( ( { 9{ ST1_03d } } & RG_rl_152 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_21 )
		| ( { 9{ U_173 } } & TR_218 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_47_en = ( ST1_03d | U_174 | RG_rl_47_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_47_en )
		RG_rl_47 <= RG_rl_47_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_60 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_217 = TR_60 ;
	7'h01 :
		TR_217 = TR_60 ;
	7'h02 :
		TR_217 = TR_60 ;
	7'h03 :
		TR_217 = TR_60 ;
	7'h04 :
		TR_217 = TR_60 ;
	7'h05 :
		TR_217 = TR_60 ;
	7'h06 :
		TR_217 = TR_60 ;
	7'h07 :
		TR_217 = TR_60 ;
	7'h08 :
		TR_217 = TR_60 ;
	7'h09 :
		TR_217 = TR_60 ;
	7'h0a :
		TR_217 = TR_60 ;
	7'h0b :
		TR_217 = TR_60 ;
	7'h0c :
		TR_217 = TR_60 ;
	7'h0d :
		TR_217 = TR_60 ;
	7'h0e :
		TR_217 = TR_60 ;
	7'h0f :
		TR_217 = TR_60 ;
	7'h10 :
		TR_217 = TR_60 ;
	7'h11 :
		TR_217 = TR_60 ;
	7'h12 :
		TR_217 = TR_60 ;
	7'h13 :
		TR_217 = TR_60 ;
	7'h14 :
		TR_217 = TR_60 ;
	7'h15 :
		TR_217 = TR_60 ;
	7'h16 :
		TR_217 = TR_60 ;
	7'h17 :
		TR_217 = TR_60 ;
	7'h18 :
		TR_217 = TR_60 ;
	7'h19 :
		TR_217 = TR_60 ;
	7'h1a :
		TR_217 = TR_60 ;
	7'h1b :
		TR_217 = TR_60 ;
	7'h1c :
		TR_217 = TR_60 ;
	7'h1d :
		TR_217 = TR_60 ;
	7'h1e :
		TR_217 = TR_60 ;
	7'h1f :
		TR_217 = TR_60 ;
	7'h20 :
		TR_217 = TR_60 ;
	7'h21 :
		TR_217 = TR_60 ;
	7'h22 :
		TR_217 = TR_60 ;
	7'h23 :
		TR_217 = TR_60 ;
	7'h24 :
		TR_217 = TR_60 ;
	7'h25 :
		TR_217 = TR_60 ;
	7'h26 :
		TR_217 = TR_60 ;
	7'h27 :
		TR_217 = TR_60 ;
	7'h28 :
		TR_217 = TR_60 ;
	7'h29 :
		TR_217 = TR_60 ;
	7'h2a :
		TR_217 = TR_60 ;
	7'h2b :
		TR_217 = TR_60 ;
	7'h2c :
		TR_217 = TR_60 ;
	7'h2d :
		TR_217 = TR_60 ;
	7'h2e :
		TR_217 = TR_60 ;
	7'h2f :
		TR_217 = TR_60 ;
	7'h30 :
		TR_217 = 9'h000 ;	// line#=../rle.cpp:80
	7'h31 :
		TR_217 = TR_60 ;
	7'h32 :
		TR_217 = TR_60 ;
	7'h33 :
		TR_217 = TR_60 ;
	7'h34 :
		TR_217 = TR_60 ;
	7'h35 :
		TR_217 = TR_60 ;
	7'h36 :
		TR_217 = TR_60 ;
	7'h37 :
		TR_217 = TR_60 ;
	7'h38 :
		TR_217 = TR_60 ;
	7'h39 :
		TR_217 = TR_60 ;
	7'h3a :
		TR_217 = TR_60 ;
	7'h3b :
		TR_217 = TR_60 ;
	7'h3c :
		TR_217 = TR_60 ;
	7'h3d :
		TR_217 = TR_60 ;
	7'h3e :
		TR_217 = TR_60 ;
	7'h3f :
		TR_217 = TR_60 ;
	7'h40 :
		TR_217 = TR_60 ;
	7'h41 :
		TR_217 = TR_60 ;
	7'h42 :
		TR_217 = TR_60 ;
	7'h43 :
		TR_217 = TR_60 ;
	7'h44 :
		TR_217 = TR_60 ;
	7'h45 :
		TR_217 = TR_60 ;
	7'h46 :
		TR_217 = TR_60 ;
	7'h47 :
		TR_217 = TR_60 ;
	7'h48 :
		TR_217 = TR_60 ;
	7'h49 :
		TR_217 = TR_60 ;
	7'h4a :
		TR_217 = TR_60 ;
	7'h4b :
		TR_217 = TR_60 ;
	7'h4c :
		TR_217 = TR_60 ;
	7'h4d :
		TR_217 = TR_60 ;
	7'h4e :
		TR_217 = TR_60 ;
	7'h4f :
		TR_217 = TR_60 ;
	7'h50 :
		TR_217 = TR_60 ;
	7'h51 :
		TR_217 = TR_60 ;
	7'h52 :
		TR_217 = TR_60 ;
	7'h53 :
		TR_217 = TR_60 ;
	7'h54 :
		TR_217 = TR_60 ;
	7'h55 :
		TR_217 = TR_60 ;
	7'h56 :
		TR_217 = TR_60 ;
	7'h57 :
		TR_217 = TR_60 ;
	7'h58 :
		TR_217 = TR_60 ;
	7'h59 :
		TR_217 = TR_60 ;
	7'h5a :
		TR_217 = TR_60 ;
	7'h5b :
		TR_217 = TR_60 ;
	7'h5c :
		TR_217 = TR_60 ;
	7'h5d :
		TR_217 = TR_60 ;
	7'h5e :
		TR_217 = TR_60 ;
	7'h5f :
		TR_217 = TR_60 ;
	7'h60 :
		TR_217 = TR_60 ;
	7'h61 :
		TR_217 = TR_60 ;
	7'h62 :
		TR_217 = TR_60 ;
	7'h63 :
		TR_217 = TR_60 ;
	7'h64 :
		TR_217 = TR_60 ;
	7'h65 :
		TR_217 = TR_60 ;
	7'h66 :
		TR_217 = TR_60 ;
	7'h67 :
		TR_217 = TR_60 ;
	7'h68 :
		TR_217 = TR_60 ;
	7'h69 :
		TR_217 = TR_60 ;
	7'h6a :
		TR_217 = TR_60 ;
	7'h6b :
		TR_217 = TR_60 ;
	7'h6c :
		TR_217 = TR_60 ;
	7'h6d :
		TR_217 = TR_60 ;
	7'h6e :
		TR_217 = TR_60 ;
	7'h6f :
		TR_217 = TR_60 ;
	7'h70 :
		TR_217 = TR_60 ;
	7'h71 :
		TR_217 = TR_60 ;
	7'h72 :
		TR_217 = TR_60 ;
	7'h73 :
		TR_217 = TR_60 ;
	7'h74 :
		TR_217 = TR_60 ;
	7'h75 :
		TR_217 = TR_60 ;
	7'h76 :
		TR_217 = TR_60 ;
	7'h77 :
		TR_217 = TR_60 ;
	7'h78 :
		TR_217 = TR_60 ;
	7'h79 :
		TR_217 = TR_60 ;
	7'h7a :
		TR_217 = TR_60 ;
	7'h7b :
		TR_217 = TR_60 ;
	7'h7c :
		TR_217 = TR_60 ;
	7'h7d :
		TR_217 = TR_60 ;
	7'h7e :
		TR_217 = TR_60 ;
	7'h7f :
		TR_217 = TR_60 ;
	default :
		TR_217 = 9'hx ;
	endcase
always @ ( TR_217 or U_173 or sub8u_71ot or U_183 or RG_rl_153 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_48_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h30 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_48_t = ( ( { 9{ M_180 } } & RG_rl_153 )
		| ( { 9{ U_173 } } & TR_217 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_48_en = ( M_180 | RG_rl_48_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_48_en )
		RG_rl_48 <= RG_rl_48_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_61 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_216 = TR_61 ;
	7'h01 :
		TR_216 = TR_61 ;
	7'h02 :
		TR_216 = TR_61 ;
	7'h03 :
		TR_216 = TR_61 ;
	7'h04 :
		TR_216 = TR_61 ;
	7'h05 :
		TR_216 = TR_61 ;
	7'h06 :
		TR_216 = TR_61 ;
	7'h07 :
		TR_216 = TR_61 ;
	7'h08 :
		TR_216 = TR_61 ;
	7'h09 :
		TR_216 = TR_61 ;
	7'h0a :
		TR_216 = TR_61 ;
	7'h0b :
		TR_216 = TR_61 ;
	7'h0c :
		TR_216 = TR_61 ;
	7'h0d :
		TR_216 = TR_61 ;
	7'h0e :
		TR_216 = TR_61 ;
	7'h0f :
		TR_216 = TR_61 ;
	7'h10 :
		TR_216 = TR_61 ;
	7'h11 :
		TR_216 = TR_61 ;
	7'h12 :
		TR_216 = TR_61 ;
	7'h13 :
		TR_216 = TR_61 ;
	7'h14 :
		TR_216 = TR_61 ;
	7'h15 :
		TR_216 = TR_61 ;
	7'h16 :
		TR_216 = TR_61 ;
	7'h17 :
		TR_216 = TR_61 ;
	7'h18 :
		TR_216 = TR_61 ;
	7'h19 :
		TR_216 = TR_61 ;
	7'h1a :
		TR_216 = TR_61 ;
	7'h1b :
		TR_216 = TR_61 ;
	7'h1c :
		TR_216 = TR_61 ;
	7'h1d :
		TR_216 = TR_61 ;
	7'h1e :
		TR_216 = TR_61 ;
	7'h1f :
		TR_216 = TR_61 ;
	7'h20 :
		TR_216 = TR_61 ;
	7'h21 :
		TR_216 = TR_61 ;
	7'h22 :
		TR_216 = TR_61 ;
	7'h23 :
		TR_216 = TR_61 ;
	7'h24 :
		TR_216 = TR_61 ;
	7'h25 :
		TR_216 = TR_61 ;
	7'h26 :
		TR_216 = TR_61 ;
	7'h27 :
		TR_216 = TR_61 ;
	7'h28 :
		TR_216 = TR_61 ;
	7'h29 :
		TR_216 = TR_61 ;
	7'h2a :
		TR_216 = TR_61 ;
	7'h2b :
		TR_216 = TR_61 ;
	7'h2c :
		TR_216 = TR_61 ;
	7'h2d :
		TR_216 = TR_61 ;
	7'h2e :
		TR_216 = TR_61 ;
	7'h2f :
		TR_216 = TR_61 ;
	7'h30 :
		TR_216 = TR_61 ;
	7'h31 :
		TR_216 = 9'h000 ;	// line#=../rle.cpp:80
	7'h32 :
		TR_216 = TR_61 ;
	7'h33 :
		TR_216 = TR_61 ;
	7'h34 :
		TR_216 = TR_61 ;
	7'h35 :
		TR_216 = TR_61 ;
	7'h36 :
		TR_216 = TR_61 ;
	7'h37 :
		TR_216 = TR_61 ;
	7'h38 :
		TR_216 = TR_61 ;
	7'h39 :
		TR_216 = TR_61 ;
	7'h3a :
		TR_216 = TR_61 ;
	7'h3b :
		TR_216 = TR_61 ;
	7'h3c :
		TR_216 = TR_61 ;
	7'h3d :
		TR_216 = TR_61 ;
	7'h3e :
		TR_216 = TR_61 ;
	7'h3f :
		TR_216 = TR_61 ;
	7'h40 :
		TR_216 = TR_61 ;
	7'h41 :
		TR_216 = TR_61 ;
	7'h42 :
		TR_216 = TR_61 ;
	7'h43 :
		TR_216 = TR_61 ;
	7'h44 :
		TR_216 = TR_61 ;
	7'h45 :
		TR_216 = TR_61 ;
	7'h46 :
		TR_216 = TR_61 ;
	7'h47 :
		TR_216 = TR_61 ;
	7'h48 :
		TR_216 = TR_61 ;
	7'h49 :
		TR_216 = TR_61 ;
	7'h4a :
		TR_216 = TR_61 ;
	7'h4b :
		TR_216 = TR_61 ;
	7'h4c :
		TR_216 = TR_61 ;
	7'h4d :
		TR_216 = TR_61 ;
	7'h4e :
		TR_216 = TR_61 ;
	7'h4f :
		TR_216 = TR_61 ;
	7'h50 :
		TR_216 = TR_61 ;
	7'h51 :
		TR_216 = TR_61 ;
	7'h52 :
		TR_216 = TR_61 ;
	7'h53 :
		TR_216 = TR_61 ;
	7'h54 :
		TR_216 = TR_61 ;
	7'h55 :
		TR_216 = TR_61 ;
	7'h56 :
		TR_216 = TR_61 ;
	7'h57 :
		TR_216 = TR_61 ;
	7'h58 :
		TR_216 = TR_61 ;
	7'h59 :
		TR_216 = TR_61 ;
	7'h5a :
		TR_216 = TR_61 ;
	7'h5b :
		TR_216 = TR_61 ;
	7'h5c :
		TR_216 = TR_61 ;
	7'h5d :
		TR_216 = TR_61 ;
	7'h5e :
		TR_216 = TR_61 ;
	7'h5f :
		TR_216 = TR_61 ;
	7'h60 :
		TR_216 = TR_61 ;
	7'h61 :
		TR_216 = TR_61 ;
	7'h62 :
		TR_216 = TR_61 ;
	7'h63 :
		TR_216 = TR_61 ;
	7'h64 :
		TR_216 = TR_61 ;
	7'h65 :
		TR_216 = TR_61 ;
	7'h66 :
		TR_216 = TR_61 ;
	7'h67 :
		TR_216 = TR_61 ;
	7'h68 :
		TR_216 = TR_61 ;
	7'h69 :
		TR_216 = TR_61 ;
	7'h6a :
		TR_216 = TR_61 ;
	7'h6b :
		TR_216 = TR_61 ;
	7'h6c :
		TR_216 = TR_61 ;
	7'h6d :
		TR_216 = TR_61 ;
	7'h6e :
		TR_216 = TR_61 ;
	7'h6f :
		TR_216 = TR_61 ;
	7'h70 :
		TR_216 = TR_61 ;
	7'h71 :
		TR_216 = TR_61 ;
	7'h72 :
		TR_216 = TR_61 ;
	7'h73 :
		TR_216 = TR_61 ;
	7'h74 :
		TR_216 = TR_61 ;
	7'h75 :
		TR_216 = TR_61 ;
	7'h76 :
		TR_216 = TR_61 ;
	7'h77 :
		TR_216 = TR_61 ;
	7'h78 :
		TR_216 = TR_61 ;
	7'h79 :
		TR_216 = TR_61 ;
	7'h7a :
		TR_216 = TR_61 ;
	7'h7b :
		TR_216 = TR_61 ;
	7'h7c :
		TR_216 = TR_61 ;
	7'h7d :
		TR_216 = TR_61 ;
	7'h7e :
		TR_216 = TR_61 ;
	7'h7f :
		TR_216 = TR_61 ;
	default :
		TR_216 = 9'hx ;
	endcase
always @ ( TR_216 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_22 or 
	U_174 or RG_rl_153 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_49_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h31 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_49_t = ( ( { 9{ ST1_03d } } & RG_rl_153 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_22 )
		| ( { 9{ U_173 } } & TR_216 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_49_en = ( ST1_03d | U_174 | RG_rl_49_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_49_en )
		RG_rl_49 <= RG_rl_49_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_62 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_215 = TR_62 ;
	7'h01 :
		TR_215 = TR_62 ;
	7'h02 :
		TR_215 = TR_62 ;
	7'h03 :
		TR_215 = TR_62 ;
	7'h04 :
		TR_215 = TR_62 ;
	7'h05 :
		TR_215 = TR_62 ;
	7'h06 :
		TR_215 = TR_62 ;
	7'h07 :
		TR_215 = TR_62 ;
	7'h08 :
		TR_215 = TR_62 ;
	7'h09 :
		TR_215 = TR_62 ;
	7'h0a :
		TR_215 = TR_62 ;
	7'h0b :
		TR_215 = TR_62 ;
	7'h0c :
		TR_215 = TR_62 ;
	7'h0d :
		TR_215 = TR_62 ;
	7'h0e :
		TR_215 = TR_62 ;
	7'h0f :
		TR_215 = TR_62 ;
	7'h10 :
		TR_215 = TR_62 ;
	7'h11 :
		TR_215 = TR_62 ;
	7'h12 :
		TR_215 = TR_62 ;
	7'h13 :
		TR_215 = TR_62 ;
	7'h14 :
		TR_215 = TR_62 ;
	7'h15 :
		TR_215 = TR_62 ;
	7'h16 :
		TR_215 = TR_62 ;
	7'h17 :
		TR_215 = TR_62 ;
	7'h18 :
		TR_215 = TR_62 ;
	7'h19 :
		TR_215 = TR_62 ;
	7'h1a :
		TR_215 = TR_62 ;
	7'h1b :
		TR_215 = TR_62 ;
	7'h1c :
		TR_215 = TR_62 ;
	7'h1d :
		TR_215 = TR_62 ;
	7'h1e :
		TR_215 = TR_62 ;
	7'h1f :
		TR_215 = TR_62 ;
	7'h20 :
		TR_215 = TR_62 ;
	7'h21 :
		TR_215 = TR_62 ;
	7'h22 :
		TR_215 = TR_62 ;
	7'h23 :
		TR_215 = TR_62 ;
	7'h24 :
		TR_215 = TR_62 ;
	7'h25 :
		TR_215 = TR_62 ;
	7'h26 :
		TR_215 = TR_62 ;
	7'h27 :
		TR_215 = TR_62 ;
	7'h28 :
		TR_215 = TR_62 ;
	7'h29 :
		TR_215 = TR_62 ;
	7'h2a :
		TR_215 = TR_62 ;
	7'h2b :
		TR_215 = TR_62 ;
	7'h2c :
		TR_215 = TR_62 ;
	7'h2d :
		TR_215 = TR_62 ;
	7'h2e :
		TR_215 = TR_62 ;
	7'h2f :
		TR_215 = TR_62 ;
	7'h30 :
		TR_215 = TR_62 ;
	7'h31 :
		TR_215 = TR_62 ;
	7'h32 :
		TR_215 = 9'h000 ;	// line#=../rle.cpp:80
	7'h33 :
		TR_215 = TR_62 ;
	7'h34 :
		TR_215 = TR_62 ;
	7'h35 :
		TR_215 = TR_62 ;
	7'h36 :
		TR_215 = TR_62 ;
	7'h37 :
		TR_215 = TR_62 ;
	7'h38 :
		TR_215 = TR_62 ;
	7'h39 :
		TR_215 = TR_62 ;
	7'h3a :
		TR_215 = TR_62 ;
	7'h3b :
		TR_215 = TR_62 ;
	7'h3c :
		TR_215 = TR_62 ;
	7'h3d :
		TR_215 = TR_62 ;
	7'h3e :
		TR_215 = TR_62 ;
	7'h3f :
		TR_215 = TR_62 ;
	7'h40 :
		TR_215 = TR_62 ;
	7'h41 :
		TR_215 = TR_62 ;
	7'h42 :
		TR_215 = TR_62 ;
	7'h43 :
		TR_215 = TR_62 ;
	7'h44 :
		TR_215 = TR_62 ;
	7'h45 :
		TR_215 = TR_62 ;
	7'h46 :
		TR_215 = TR_62 ;
	7'h47 :
		TR_215 = TR_62 ;
	7'h48 :
		TR_215 = TR_62 ;
	7'h49 :
		TR_215 = TR_62 ;
	7'h4a :
		TR_215 = TR_62 ;
	7'h4b :
		TR_215 = TR_62 ;
	7'h4c :
		TR_215 = TR_62 ;
	7'h4d :
		TR_215 = TR_62 ;
	7'h4e :
		TR_215 = TR_62 ;
	7'h4f :
		TR_215 = TR_62 ;
	7'h50 :
		TR_215 = TR_62 ;
	7'h51 :
		TR_215 = TR_62 ;
	7'h52 :
		TR_215 = TR_62 ;
	7'h53 :
		TR_215 = TR_62 ;
	7'h54 :
		TR_215 = TR_62 ;
	7'h55 :
		TR_215 = TR_62 ;
	7'h56 :
		TR_215 = TR_62 ;
	7'h57 :
		TR_215 = TR_62 ;
	7'h58 :
		TR_215 = TR_62 ;
	7'h59 :
		TR_215 = TR_62 ;
	7'h5a :
		TR_215 = TR_62 ;
	7'h5b :
		TR_215 = TR_62 ;
	7'h5c :
		TR_215 = TR_62 ;
	7'h5d :
		TR_215 = TR_62 ;
	7'h5e :
		TR_215 = TR_62 ;
	7'h5f :
		TR_215 = TR_62 ;
	7'h60 :
		TR_215 = TR_62 ;
	7'h61 :
		TR_215 = TR_62 ;
	7'h62 :
		TR_215 = TR_62 ;
	7'h63 :
		TR_215 = TR_62 ;
	7'h64 :
		TR_215 = TR_62 ;
	7'h65 :
		TR_215 = TR_62 ;
	7'h66 :
		TR_215 = TR_62 ;
	7'h67 :
		TR_215 = TR_62 ;
	7'h68 :
		TR_215 = TR_62 ;
	7'h69 :
		TR_215 = TR_62 ;
	7'h6a :
		TR_215 = TR_62 ;
	7'h6b :
		TR_215 = TR_62 ;
	7'h6c :
		TR_215 = TR_62 ;
	7'h6d :
		TR_215 = TR_62 ;
	7'h6e :
		TR_215 = TR_62 ;
	7'h6f :
		TR_215 = TR_62 ;
	7'h70 :
		TR_215 = TR_62 ;
	7'h71 :
		TR_215 = TR_62 ;
	7'h72 :
		TR_215 = TR_62 ;
	7'h73 :
		TR_215 = TR_62 ;
	7'h74 :
		TR_215 = TR_62 ;
	7'h75 :
		TR_215 = TR_62 ;
	7'h76 :
		TR_215 = TR_62 ;
	7'h77 :
		TR_215 = TR_62 ;
	7'h78 :
		TR_215 = TR_62 ;
	7'h79 :
		TR_215 = TR_62 ;
	7'h7a :
		TR_215 = TR_62 ;
	7'h7b :
		TR_215 = TR_62 ;
	7'h7c :
		TR_215 = TR_62 ;
	7'h7d :
		TR_215 = TR_62 ;
	7'h7e :
		TR_215 = TR_62 ;
	7'h7f :
		TR_215 = TR_62 ;
	default :
		TR_215 = 9'hx ;
	endcase
always @ ( TR_215 or U_173 or sub8u_71ot or U_183 or RG_rl_154 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_50_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h32 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_50_t = ( ( { 9{ M_180 } } & RG_rl_154 )
		| ( { 9{ U_173 } } & TR_215 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_50_en = ( M_180 | RG_rl_50_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_50_en )
		RG_rl_50 <= RG_rl_50_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_63 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_214 = TR_63 ;
	7'h01 :
		TR_214 = TR_63 ;
	7'h02 :
		TR_214 = TR_63 ;
	7'h03 :
		TR_214 = TR_63 ;
	7'h04 :
		TR_214 = TR_63 ;
	7'h05 :
		TR_214 = TR_63 ;
	7'h06 :
		TR_214 = TR_63 ;
	7'h07 :
		TR_214 = TR_63 ;
	7'h08 :
		TR_214 = TR_63 ;
	7'h09 :
		TR_214 = TR_63 ;
	7'h0a :
		TR_214 = TR_63 ;
	7'h0b :
		TR_214 = TR_63 ;
	7'h0c :
		TR_214 = TR_63 ;
	7'h0d :
		TR_214 = TR_63 ;
	7'h0e :
		TR_214 = TR_63 ;
	7'h0f :
		TR_214 = TR_63 ;
	7'h10 :
		TR_214 = TR_63 ;
	7'h11 :
		TR_214 = TR_63 ;
	7'h12 :
		TR_214 = TR_63 ;
	7'h13 :
		TR_214 = TR_63 ;
	7'h14 :
		TR_214 = TR_63 ;
	7'h15 :
		TR_214 = TR_63 ;
	7'h16 :
		TR_214 = TR_63 ;
	7'h17 :
		TR_214 = TR_63 ;
	7'h18 :
		TR_214 = TR_63 ;
	7'h19 :
		TR_214 = TR_63 ;
	7'h1a :
		TR_214 = TR_63 ;
	7'h1b :
		TR_214 = TR_63 ;
	7'h1c :
		TR_214 = TR_63 ;
	7'h1d :
		TR_214 = TR_63 ;
	7'h1e :
		TR_214 = TR_63 ;
	7'h1f :
		TR_214 = TR_63 ;
	7'h20 :
		TR_214 = TR_63 ;
	7'h21 :
		TR_214 = TR_63 ;
	7'h22 :
		TR_214 = TR_63 ;
	7'h23 :
		TR_214 = TR_63 ;
	7'h24 :
		TR_214 = TR_63 ;
	7'h25 :
		TR_214 = TR_63 ;
	7'h26 :
		TR_214 = TR_63 ;
	7'h27 :
		TR_214 = TR_63 ;
	7'h28 :
		TR_214 = TR_63 ;
	7'h29 :
		TR_214 = TR_63 ;
	7'h2a :
		TR_214 = TR_63 ;
	7'h2b :
		TR_214 = TR_63 ;
	7'h2c :
		TR_214 = TR_63 ;
	7'h2d :
		TR_214 = TR_63 ;
	7'h2e :
		TR_214 = TR_63 ;
	7'h2f :
		TR_214 = TR_63 ;
	7'h30 :
		TR_214 = TR_63 ;
	7'h31 :
		TR_214 = TR_63 ;
	7'h32 :
		TR_214 = TR_63 ;
	7'h33 :
		TR_214 = 9'h000 ;	// line#=../rle.cpp:80
	7'h34 :
		TR_214 = TR_63 ;
	7'h35 :
		TR_214 = TR_63 ;
	7'h36 :
		TR_214 = TR_63 ;
	7'h37 :
		TR_214 = TR_63 ;
	7'h38 :
		TR_214 = TR_63 ;
	7'h39 :
		TR_214 = TR_63 ;
	7'h3a :
		TR_214 = TR_63 ;
	7'h3b :
		TR_214 = TR_63 ;
	7'h3c :
		TR_214 = TR_63 ;
	7'h3d :
		TR_214 = TR_63 ;
	7'h3e :
		TR_214 = TR_63 ;
	7'h3f :
		TR_214 = TR_63 ;
	7'h40 :
		TR_214 = TR_63 ;
	7'h41 :
		TR_214 = TR_63 ;
	7'h42 :
		TR_214 = TR_63 ;
	7'h43 :
		TR_214 = TR_63 ;
	7'h44 :
		TR_214 = TR_63 ;
	7'h45 :
		TR_214 = TR_63 ;
	7'h46 :
		TR_214 = TR_63 ;
	7'h47 :
		TR_214 = TR_63 ;
	7'h48 :
		TR_214 = TR_63 ;
	7'h49 :
		TR_214 = TR_63 ;
	7'h4a :
		TR_214 = TR_63 ;
	7'h4b :
		TR_214 = TR_63 ;
	7'h4c :
		TR_214 = TR_63 ;
	7'h4d :
		TR_214 = TR_63 ;
	7'h4e :
		TR_214 = TR_63 ;
	7'h4f :
		TR_214 = TR_63 ;
	7'h50 :
		TR_214 = TR_63 ;
	7'h51 :
		TR_214 = TR_63 ;
	7'h52 :
		TR_214 = TR_63 ;
	7'h53 :
		TR_214 = TR_63 ;
	7'h54 :
		TR_214 = TR_63 ;
	7'h55 :
		TR_214 = TR_63 ;
	7'h56 :
		TR_214 = TR_63 ;
	7'h57 :
		TR_214 = TR_63 ;
	7'h58 :
		TR_214 = TR_63 ;
	7'h59 :
		TR_214 = TR_63 ;
	7'h5a :
		TR_214 = TR_63 ;
	7'h5b :
		TR_214 = TR_63 ;
	7'h5c :
		TR_214 = TR_63 ;
	7'h5d :
		TR_214 = TR_63 ;
	7'h5e :
		TR_214 = TR_63 ;
	7'h5f :
		TR_214 = TR_63 ;
	7'h60 :
		TR_214 = TR_63 ;
	7'h61 :
		TR_214 = TR_63 ;
	7'h62 :
		TR_214 = TR_63 ;
	7'h63 :
		TR_214 = TR_63 ;
	7'h64 :
		TR_214 = TR_63 ;
	7'h65 :
		TR_214 = TR_63 ;
	7'h66 :
		TR_214 = TR_63 ;
	7'h67 :
		TR_214 = TR_63 ;
	7'h68 :
		TR_214 = TR_63 ;
	7'h69 :
		TR_214 = TR_63 ;
	7'h6a :
		TR_214 = TR_63 ;
	7'h6b :
		TR_214 = TR_63 ;
	7'h6c :
		TR_214 = TR_63 ;
	7'h6d :
		TR_214 = TR_63 ;
	7'h6e :
		TR_214 = TR_63 ;
	7'h6f :
		TR_214 = TR_63 ;
	7'h70 :
		TR_214 = TR_63 ;
	7'h71 :
		TR_214 = TR_63 ;
	7'h72 :
		TR_214 = TR_63 ;
	7'h73 :
		TR_214 = TR_63 ;
	7'h74 :
		TR_214 = TR_63 ;
	7'h75 :
		TR_214 = TR_63 ;
	7'h76 :
		TR_214 = TR_63 ;
	7'h77 :
		TR_214 = TR_63 ;
	7'h78 :
		TR_214 = TR_63 ;
	7'h79 :
		TR_214 = TR_63 ;
	7'h7a :
		TR_214 = TR_63 ;
	7'h7b :
		TR_214 = TR_63 ;
	7'h7c :
		TR_214 = TR_63 ;
	7'h7d :
		TR_214 = TR_63 ;
	7'h7e :
		TR_214 = TR_63 ;
	7'h7f :
		TR_214 = TR_63 ;
	default :
		TR_214 = 9'hx ;
	endcase
always @ ( TR_214 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_23 or 
	U_174 or RG_rl_154 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_51_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h33 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_51_t = ( ( { 9{ ST1_03d } } & RG_rl_154 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_23 )
		| ( { 9{ U_173 } } & TR_214 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_51_en = ( ST1_03d | U_174 | RG_rl_51_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_51_en )
		RG_rl_51 <= RG_rl_51_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_64 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_213 = TR_64 ;
	7'h01 :
		TR_213 = TR_64 ;
	7'h02 :
		TR_213 = TR_64 ;
	7'h03 :
		TR_213 = TR_64 ;
	7'h04 :
		TR_213 = TR_64 ;
	7'h05 :
		TR_213 = TR_64 ;
	7'h06 :
		TR_213 = TR_64 ;
	7'h07 :
		TR_213 = TR_64 ;
	7'h08 :
		TR_213 = TR_64 ;
	7'h09 :
		TR_213 = TR_64 ;
	7'h0a :
		TR_213 = TR_64 ;
	7'h0b :
		TR_213 = TR_64 ;
	7'h0c :
		TR_213 = TR_64 ;
	7'h0d :
		TR_213 = TR_64 ;
	7'h0e :
		TR_213 = TR_64 ;
	7'h0f :
		TR_213 = TR_64 ;
	7'h10 :
		TR_213 = TR_64 ;
	7'h11 :
		TR_213 = TR_64 ;
	7'h12 :
		TR_213 = TR_64 ;
	7'h13 :
		TR_213 = TR_64 ;
	7'h14 :
		TR_213 = TR_64 ;
	7'h15 :
		TR_213 = TR_64 ;
	7'h16 :
		TR_213 = TR_64 ;
	7'h17 :
		TR_213 = TR_64 ;
	7'h18 :
		TR_213 = TR_64 ;
	7'h19 :
		TR_213 = TR_64 ;
	7'h1a :
		TR_213 = TR_64 ;
	7'h1b :
		TR_213 = TR_64 ;
	7'h1c :
		TR_213 = TR_64 ;
	7'h1d :
		TR_213 = TR_64 ;
	7'h1e :
		TR_213 = TR_64 ;
	7'h1f :
		TR_213 = TR_64 ;
	7'h20 :
		TR_213 = TR_64 ;
	7'h21 :
		TR_213 = TR_64 ;
	7'h22 :
		TR_213 = TR_64 ;
	7'h23 :
		TR_213 = TR_64 ;
	7'h24 :
		TR_213 = TR_64 ;
	7'h25 :
		TR_213 = TR_64 ;
	7'h26 :
		TR_213 = TR_64 ;
	7'h27 :
		TR_213 = TR_64 ;
	7'h28 :
		TR_213 = TR_64 ;
	7'h29 :
		TR_213 = TR_64 ;
	7'h2a :
		TR_213 = TR_64 ;
	7'h2b :
		TR_213 = TR_64 ;
	7'h2c :
		TR_213 = TR_64 ;
	7'h2d :
		TR_213 = TR_64 ;
	7'h2e :
		TR_213 = TR_64 ;
	7'h2f :
		TR_213 = TR_64 ;
	7'h30 :
		TR_213 = TR_64 ;
	7'h31 :
		TR_213 = TR_64 ;
	7'h32 :
		TR_213 = TR_64 ;
	7'h33 :
		TR_213 = TR_64 ;
	7'h34 :
		TR_213 = 9'h000 ;	// line#=../rle.cpp:80
	7'h35 :
		TR_213 = TR_64 ;
	7'h36 :
		TR_213 = TR_64 ;
	7'h37 :
		TR_213 = TR_64 ;
	7'h38 :
		TR_213 = TR_64 ;
	7'h39 :
		TR_213 = TR_64 ;
	7'h3a :
		TR_213 = TR_64 ;
	7'h3b :
		TR_213 = TR_64 ;
	7'h3c :
		TR_213 = TR_64 ;
	7'h3d :
		TR_213 = TR_64 ;
	7'h3e :
		TR_213 = TR_64 ;
	7'h3f :
		TR_213 = TR_64 ;
	7'h40 :
		TR_213 = TR_64 ;
	7'h41 :
		TR_213 = TR_64 ;
	7'h42 :
		TR_213 = TR_64 ;
	7'h43 :
		TR_213 = TR_64 ;
	7'h44 :
		TR_213 = TR_64 ;
	7'h45 :
		TR_213 = TR_64 ;
	7'h46 :
		TR_213 = TR_64 ;
	7'h47 :
		TR_213 = TR_64 ;
	7'h48 :
		TR_213 = TR_64 ;
	7'h49 :
		TR_213 = TR_64 ;
	7'h4a :
		TR_213 = TR_64 ;
	7'h4b :
		TR_213 = TR_64 ;
	7'h4c :
		TR_213 = TR_64 ;
	7'h4d :
		TR_213 = TR_64 ;
	7'h4e :
		TR_213 = TR_64 ;
	7'h4f :
		TR_213 = TR_64 ;
	7'h50 :
		TR_213 = TR_64 ;
	7'h51 :
		TR_213 = TR_64 ;
	7'h52 :
		TR_213 = TR_64 ;
	7'h53 :
		TR_213 = TR_64 ;
	7'h54 :
		TR_213 = TR_64 ;
	7'h55 :
		TR_213 = TR_64 ;
	7'h56 :
		TR_213 = TR_64 ;
	7'h57 :
		TR_213 = TR_64 ;
	7'h58 :
		TR_213 = TR_64 ;
	7'h59 :
		TR_213 = TR_64 ;
	7'h5a :
		TR_213 = TR_64 ;
	7'h5b :
		TR_213 = TR_64 ;
	7'h5c :
		TR_213 = TR_64 ;
	7'h5d :
		TR_213 = TR_64 ;
	7'h5e :
		TR_213 = TR_64 ;
	7'h5f :
		TR_213 = TR_64 ;
	7'h60 :
		TR_213 = TR_64 ;
	7'h61 :
		TR_213 = TR_64 ;
	7'h62 :
		TR_213 = TR_64 ;
	7'h63 :
		TR_213 = TR_64 ;
	7'h64 :
		TR_213 = TR_64 ;
	7'h65 :
		TR_213 = TR_64 ;
	7'h66 :
		TR_213 = TR_64 ;
	7'h67 :
		TR_213 = TR_64 ;
	7'h68 :
		TR_213 = TR_64 ;
	7'h69 :
		TR_213 = TR_64 ;
	7'h6a :
		TR_213 = TR_64 ;
	7'h6b :
		TR_213 = TR_64 ;
	7'h6c :
		TR_213 = TR_64 ;
	7'h6d :
		TR_213 = TR_64 ;
	7'h6e :
		TR_213 = TR_64 ;
	7'h6f :
		TR_213 = TR_64 ;
	7'h70 :
		TR_213 = TR_64 ;
	7'h71 :
		TR_213 = TR_64 ;
	7'h72 :
		TR_213 = TR_64 ;
	7'h73 :
		TR_213 = TR_64 ;
	7'h74 :
		TR_213 = TR_64 ;
	7'h75 :
		TR_213 = TR_64 ;
	7'h76 :
		TR_213 = TR_64 ;
	7'h77 :
		TR_213 = TR_64 ;
	7'h78 :
		TR_213 = TR_64 ;
	7'h79 :
		TR_213 = TR_64 ;
	7'h7a :
		TR_213 = TR_64 ;
	7'h7b :
		TR_213 = TR_64 ;
	7'h7c :
		TR_213 = TR_64 ;
	7'h7d :
		TR_213 = TR_64 ;
	7'h7e :
		TR_213 = TR_64 ;
	7'h7f :
		TR_213 = TR_64 ;
	default :
		TR_213 = 9'hx ;
	endcase
always @ ( TR_213 or U_173 or sub8u_71ot or U_183 or RG_rl_155 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_52_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h34 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_52_t = ( ( { 9{ M_180 } } & RG_rl_155 )
		| ( { 9{ U_173 } } & TR_213 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_52_en = ( M_180 | RG_rl_52_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_52_en )
		RG_rl_52 <= RG_rl_52_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_65 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_212 = TR_65 ;
	7'h01 :
		TR_212 = TR_65 ;
	7'h02 :
		TR_212 = TR_65 ;
	7'h03 :
		TR_212 = TR_65 ;
	7'h04 :
		TR_212 = TR_65 ;
	7'h05 :
		TR_212 = TR_65 ;
	7'h06 :
		TR_212 = TR_65 ;
	7'h07 :
		TR_212 = TR_65 ;
	7'h08 :
		TR_212 = TR_65 ;
	7'h09 :
		TR_212 = TR_65 ;
	7'h0a :
		TR_212 = TR_65 ;
	7'h0b :
		TR_212 = TR_65 ;
	7'h0c :
		TR_212 = TR_65 ;
	7'h0d :
		TR_212 = TR_65 ;
	7'h0e :
		TR_212 = TR_65 ;
	7'h0f :
		TR_212 = TR_65 ;
	7'h10 :
		TR_212 = TR_65 ;
	7'h11 :
		TR_212 = TR_65 ;
	7'h12 :
		TR_212 = TR_65 ;
	7'h13 :
		TR_212 = TR_65 ;
	7'h14 :
		TR_212 = TR_65 ;
	7'h15 :
		TR_212 = TR_65 ;
	7'h16 :
		TR_212 = TR_65 ;
	7'h17 :
		TR_212 = TR_65 ;
	7'h18 :
		TR_212 = TR_65 ;
	7'h19 :
		TR_212 = TR_65 ;
	7'h1a :
		TR_212 = TR_65 ;
	7'h1b :
		TR_212 = TR_65 ;
	7'h1c :
		TR_212 = TR_65 ;
	7'h1d :
		TR_212 = TR_65 ;
	7'h1e :
		TR_212 = TR_65 ;
	7'h1f :
		TR_212 = TR_65 ;
	7'h20 :
		TR_212 = TR_65 ;
	7'h21 :
		TR_212 = TR_65 ;
	7'h22 :
		TR_212 = TR_65 ;
	7'h23 :
		TR_212 = TR_65 ;
	7'h24 :
		TR_212 = TR_65 ;
	7'h25 :
		TR_212 = TR_65 ;
	7'h26 :
		TR_212 = TR_65 ;
	7'h27 :
		TR_212 = TR_65 ;
	7'h28 :
		TR_212 = TR_65 ;
	7'h29 :
		TR_212 = TR_65 ;
	7'h2a :
		TR_212 = TR_65 ;
	7'h2b :
		TR_212 = TR_65 ;
	7'h2c :
		TR_212 = TR_65 ;
	7'h2d :
		TR_212 = TR_65 ;
	7'h2e :
		TR_212 = TR_65 ;
	7'h2f :
		TR_212 = TR_65 ;
	7'h30 :
		TR_212 = TR_65 ;
	7'h31 :
		TR_212 = TR_65 ;
	7'h32 :
		TR_212 = TR_65 ;
	7'h33 :
		TR_212 = TR_65 ;
	7'h34 :
		TR_212 = TR_65 ;
	7'h35 :
		TR_212 = 9'h000 ;	// line#=../rle.cpp:80
	7'h36 :
		TR_212 = TR_65 ;
	7'h37 :
		TR_212 = TR_65 ;
	7'h38 :
		TR_212 = TR_65 ;
	7'h39 :
		TR_212 = TR_65 ;
	7'h3a :
		TR_212 = TR_65 ;
	7'h3b :
		TR_212 = TR_65 ;
	7'h3c :
		TR_212 = TR_65 ;
	7'h3d :
		TR_212 = TR_65 ;
	7'h3e :
		TR_212 = TR_65 ;
	7'h3f :
		TR_212 = TR_65 ;
	7'h40 :
		TR_212 = TR_65 ;
	7'h41 :
		TR_212 = TR_65 ;
	7'h42 :
		TR_212 = TR_65 ;
	7'h43 :
		TR_212 = TR_65 ;
	7'h44 :
		TR_212 = TR_65 ;
	7'h45 :
		TR_212 = TR_65 ;
	7'h46 :
		TR_212 = TR_65 ;
	7'h47 :
		TR_212 = TR_65 ;
	7'h48 :
		TR_212 = TR_65 ;
	7'h49 :
		TR_212 = TR_65 ;
	7'h4a :
		TR_212 = TR_65 ;
	7'h4b :
		TR_212 = TR_65 ;
	7'h4c :
		TR_212 = TR_65 ;
	7'h4d :
		TR_212 = TR_65 ;
	7'h4e :
		TR_212 = TR_65 ;
	7'h4f :
		TR_212 = TR_65 ;
	7'h50 :
		TR_212 = TR_65 ;
	7'h51 :
		TR_212 = TR_65 ;
	7'h52 :
		TR_212 = TR_65 ;
	7'h53 :
		TR_212 = TR_65 ;
	7'h54 :
		TR_212 = TR_65 ;
	7'h55 :
		TR_212 = TR_65 ;
	7'h56 :
		TR_212 = TR_65 ;
	7'h57 :
		TR_212 = TR_65 ;
	7'h58 :
		TR_212 = TR_65 ;
	7'h59 :
		TR_212 = TR_65 ;
	7'h5a :
		TR_212 = TR_65 ;
	7'h5b :
		TR_212 = TR_65 ;
	7'h5c :
		TR_212 = TR_65 ;
	7'h5d :
		TR_212 = TR_65 ;
	7'h5e :
		TR_212 = TR_65 ;
	7'h5f :
		TR_212 = TR_65 ;
	7'h60 :
		TR_212 = TR_65 ;
	7'h61 :
		TR_212 = TR_65 ;
	7'h62 :
		TR_212 = TR_65 ;
	7'h63 :
		TR_212 = TR_65 ;
	7'h64 :
		TR_212 = TR_65 ;
	7'h65 :
		TR_212 = TR_65 ;
	7'h66 :
		TR_212 = TR_65 ;
	7'h67 :
		TR_212 = TR_65 ;
	7'h68 :
		TR_212 = TR_65 ;
	7'h69 :
		TR_212 = TR_65 ;
	7'h6a :
		TR_212 = TR_65 ;
	7'h6b :
		TR_212 = TR_65 ;
	7'h6c :
		TR_212 = TR_65 ;
	7'h6d :
		TR_212 = TR_65 ;
	7'h6e :
		TR_212 = TR_65 ;
	7'h6f :
		TR_212 = TR_65 ;
	7'h70 :
		TR_212 = TR_65 ;
	7'h71 :
		TR_212 = TR_65 ;
	7'h72 :
		TR_212 = TR_65 ;
	7'h73 :
		TR_212 = TR_65 ;
	7'h74 :
		TR_212 = TR_65 ;
	7'h75 :
		TR_212 = TR_65 ;
	7'h76 :
		TR_212 = TR_65 ;
	7'h77 :
		TR_212 = TR_65 ;
	7'h78 :
		TR_212 = TR_65 ;
	7'h79 :
		TR_212 = TR_65 ;
	7'h7a :
		TR_212 = TR_65 ;
	7'h7b :
		TR_212 = TR_65 ;
	7'h7c :
		TR_212 = TR_65 ;
	7'h7d :
		TR_212 = TR_65 ;
	7'h7e :
		TR_212 = TR_65 ;
	7'h7f :
		TR_212 = TR_65 ;
	default :
		TR_212 = 9'hx ;
	endcase
always @ ( TR_212 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_24 or 
	U_174 or RG_rl_155 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_53_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h35 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_53_t = ( ( { 9{ ST1_03d } } & RG_rl_155 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_24 )
		| ( { 9{ U_173 } } & TR_212 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_53_en = ( ST1_03d | U_174 | RG_rl_53_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_53_en )
		RG_rl_53 <= RG_rl_53_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_66 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_211 = TR_66 ;
	7'h01 :
		TR_211 = TR_66 ;
	7'h02 :
		TR_211 = TR_66 ;
	7'h03 :
		TR_211 = TR_66 ;
	7'h04 :
		TR_211 = TR_66 ;
	7'h05 :
		TR_211 = TR_66 ;
	7'h06 :
		TR_211 = TR_66 ;
	7'h07 :
		TR_211 = TR_66 ;
	7'h08 :
		TR_211 = TR_66 ;
	7'h09 :
		TR_211 = TR_66 ;
	7'h0a :
		TR_211 = TR_66 ;
	7'h0b :
		TR_211 = TR_66 ;
	7'h0c :
		TR_211 = TR_66 ;
	7'h0d :
		TR_211 = TR_66 ;
	7'h0e :
		TR_211 = TR_66 ;
	7'h0f :
		TR_211 = TR_66 ;
	7'h10 :
		TR_211 = TR_66 ;
	7'h11 :
		TR_211 = TR_66 ;
	7'h12 :
		TR_211 = TR_66 ;
	7'h13 :
		TR_211 = TR_66 ;
	7'h14 :
		TR_211 = TR_66 ;
	7'h15 :
		TR_211 = TR_66 ;
	7'h16 :
		TR_211 = TR_66 ;
	7'h17 :
		TR_211 = TR_66 ;
	7'h18 :
		TR_211 = TR_66 ;
	7'h19 :
		TR_211 = TR_66 ;
	7'h1a :
		TR_211 = TR_66 ;
	7'h1b :
		TR_211 = TR_66 ;
	7'h1c :
		TR_211 = TR_66 ;
	7'h1d :
		TR_211 = TR_66 ;
	7'h1e :
		TR_211 = TR_66 ;
	7'h1f :
		TR_211 = TR_66 ;
	7'h20 :
		TR_211 = TR_66 ;
	7'h21 :
		TR_211 = TR_66 ;
	7'h22 :
		TR_211 = TR_66 ;
	7'h23 :
		TR_211 = TR_66 ;
	7'h24 :
		TR_211 = TR_66 ;
	7'h25 :
		TR_211 = TR_66 ;
	7'h26 :
		TR_211 = TR_66 ;
	7'h27 :
		TR_211 = TR_66 ;
	7'h28 :
		TR_211 = TR_66 ;
	7'h29 :
		TR_211 = TR_66 ;
	7'h2a :
		TR_211 = TR_66 ;
	7'h2b :
		TR_211 = TR_66 ;
	7'h2c :
		TR_211 = TR_66 ;
	7'h2d :
		TR_211 = TR_66 ;
	7'h2e :
		TR_211 = TR_66 ;
	7'h2f :
		TR_211 = TR_66 ;
	7'h30 :
		TR_211 = TR_66 ;
	7'h31 :
		TR_211 = TR_66 ;
	7'h32 :
		TR_211 = TR_66 ;
	7'h33 :
		TR_211 = TR_66 ;
	7'h34 :
		TR_211 = TR_66 ;
	7'h35 :
		TR_211 = TR_66 ;
	7'h36 :
		TR_211 = 9'h000 ;	// line#=../rle.cpp:80
	7'h37 :
		TR_211 = TR_66 ;
	7'h38 :
		TR_211 = TR_66 ;
	7'h39 :
		TR_211 = TR_66 ;
	7'h3a :
		TR_211 = TR_66 ;
	7'h3b :
		TR_211 = TR_66 ;
	7'h3c :
		TR_211 = TR_66 ;
	7'h3d :
		TR_211 = TR_66 ;
	7'h3e :
		TR_211 = TR_66 ;
	7'h3f :
		TR_211 = TR_66 ;
	7'h40 :
		TR_211 = TR_66 ;
	7'h41 :
		TR_211 = TR_66 ;
	7'h42 :
		TR_211 = TR_66 ;
	7'h43 :
		TR_211 = TR_66 ;
	7'h44 :
		TR_211 = TR_66 ;
	7'h45 :
		TR_211 = TR_66 ;
	7'h46 :
		TR_211 = TR_66 ;
	7'h47 :
		TR_211 = TR_66 ;
	7'h48 :
		TR_211 = TR_66 ;
	7'h49 :
		TR_211 = TR_66 ;
	7'h4a :
		TR_211 = TR_66 ;
	7'h4b :
		TR_211 = TR_66 ;
	7'h4c :
		TR_211 = TR_66 ;
	7'h4d :
		TR_211 = TR_66 ;
	7'h4e :
		TR_211 = TR_66 ;
	7'h4f :
		TR_211 = TR_66 ;
	7'h50 :
		TR_211 = TR_66 ;
	7'h51 :
		TR_211 = TR_66 ;
	7'h52 :
		TR_211 = TR_66 ;
	7'h53 :
		TR_211 = TR_66 ;
	7'h54 :
		TR_211 = TR_66 ;
	7'h55 :
		TR_211 = TR_66 ;
	7'h56 :
		TR_211 = TR_66 ;
	7'h57 :
		TR_211 = TR_66 ;
	7'h58 :
		TR_211 = TR_66 ;
	7'h59 :
		TR_211 = TR_66 ;
	7'h5a :
		TR_211 = TR_66 ;
	7'h5b :
		TR_211 = TR_66 ;
	7'h5c :
		TR_211 = TR_66 ;
	7'h5d :
		TR_211 = TR_66 ;
	7'h5e :
		TR_211 = TR_66 ;
	7'h5f :
		TR_211 = TR_66 ;
	7'h60 :
		TR_211 = TR_66 ;
	7'h61 :
		TR_211 = TR_66 ;
	7'h62 :
		TR_211 = TR_66 ;
	7'h63 :
		TR_211 = TR_66 ;
	7'h64 :
		TR_211 = TR_66 ;
	7'h65 :
		TR_211 = TR_66 ;
	7'h66 :
		TR_211 = TR_66 ;
	7'h67 :
		TR_211 = TR_66 ;
	7'h68 :
		TR_211 = TR_66 ;
	7'h69 :
		TR_211 = TR_66 ;
	7'h6a :
		TR_211 = TR_66 ;
	7'h6b :
		TR_211 = TR_66 ;
	7'h6c :
		TR_211 = TR_66 ;
	7'h6d :
		TR_211 = TR_66 ;
	7'h6e :
		TR_211 = TR_66 ;
	7'h6f :
		TR_211 = TR_66 ;
	7'h70 :
		TR_211 = TR_66 ;
	7'h71 :
		TR_211 = TR_66 ;
	7'h72 :
		TR_211 = TR_66 ;
	7'h73 :
		TR_211 = TR_66 ;
	7'h74 :
		TR_211 = TR_66 ;
	7'h75 :
		TR_211 = TR_66 ;
	7'h76 :
		TR_211 = TR_66 ;
	7'h77 :
		TR_211 = TR_66 ;
	7'h78 :
		TR_211 = TR_66 ;
	7'h79 :
		TR_211 = TR_66 ;
	7'h7a :
		TR_211 = TR_66 ;
	7'h7b :
		TR_211 = TR_66 ;
	7'h7c :
		TR_211 = TR_66 ;
	7'h7d :
		TR_211 = TR_66 ;
	7'h7e :
		TR_211 = TR_66 ;
	7'h7f :
		TR_211 = TR_66 ;
	default :
		TR_211 = 9'hx ;
	endcase
always @ ( TR_211 or U_173 or sub8u_71ot or U_183 or RG_rl_156 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_54_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h36 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_54_t = ( ( { 9{ M_180 } } & RG_rl_156 )
		| ( { 9{ U_173 } } & TR_211 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_54_en = ( M_180 | RG_rl_54_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_54_en )
		RG_rl_54 <= RG_rl_54_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_67 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_210 = TR_67 ;
	7'h01 :
		TR_210 = TR_67 ;
	7'h02 :
		TR_210 = TR_67 ;
	7'h03 :
		TR_210 = TR_67 ;
	7'h04 :
		TR_210 = TR_67 ;
	7'h05 :
		TR_210 = TR_67 ;
	7'h06 :
		TR_210 = TR_67 ;
	7'h07 :
		TR_210 = TR_67 ;
	7'h08 :
		TR_210 = TR_67 ;
	7'h09 :
		TR_210 = TR_67 ;
	7'h0a :
		TR_210 = TR_67 ;
	7'h0b :
		TR_210 = TR_67 ;
	7'h0c :
		TR_210 = TR_67 ;
	7'h0d :
		TR_210 = TR_67 ;
	7'h0e :
		TR_210 = TR_67 ;
	7'h0f :
		TR_210 = TR_67 ;
	7'h10 :
		TR_210 = TR_67 ;
	7'h11 :
		TR_210 = TR_67 ;
	7'h12 :
		TR_210 = TR_67 ;
	7'h13 :
		TR_210 = TR_67 ;
	7'h14 :
		TR_210 = TR_67 ;
	7'h15 :
		TR_210 = TR_67 ;
	7'h16 :
		TR_210 = TR_67 ;
	7'h17 :
		TR_210 = TR_67 ;
	7'h18 :
		TR_210 = TR_67 ;
	7'h19 :
		TR_210 = TR_67 ;
	7'h1a :
		TR_210 = TR_67 ;
	7'h1b :
		TR_210 = TR_67 ;
	7'h1c :
		TR_210 = TR_67 ;
	7'h1d :
		TR_210 = TR_67 ;
	7'h1e :
		TR_210 = TR_67 ;
	7'h1f :
		TR_210 = TR_67 ;
	7'h20 :
		TR_210 = TR_67 ;
	7'h21 :
		TR_210 = TR_67 ;
	7'h22 :
		TR_210 = TR_67 ;
	7'h23 :
		TR_210 = TR_67 ;
	7'h24 :
		TR_210 = TR_67 ;
	7'h25 :
		TR_210 = TR_67 ;
	7'h26 :
		TR_210 = TR_67 ;
	7'h27 :
		TR_210 = TR_67 ;
	7'h28 :
		TR_210 = TR_67 ;
	7'h29 :
		TR_210 = TR_67 ;
	7'h2a :
		TR_210 = TR_67 ;
	7'h2b :
		TR_210 = TR_67 ;
	7'h2c :
		TR_210 = TR_67 ;
	7'h2d :
		TR_210 = TR_67 ;
	7'h2e :
		TR_210 = TR_67 ;
	7'h2f :
		TR_210 = TR_67 ;
	7'h30 :
		TR_210 = TR_67 ;
	7'h31 :
		TR_210 = TR_67 ;
	7'h32 :
		TR_210 = TR_67 ;
	7'h33 :
		TR_210 = TR_67 ;
	7'h34 :
		TR_210 = TR_67 ;
	7'h35 :
		TR_210 = TR_67 ;
	7'h36 :
		TR_210 = TR_67 ;
	7'h37 :
		TR_210 = 9'h000 ;	// line#=../rle.cpp:80
	7'h38 :
		TR_210 = TR_67 ;
	7'h39 :
		TR_210 = TR_67 ;
	7'h3a :
		TR_210 = TR_67 ;
	7'h3b :
		TR_210 = TR_67 ;
	7'h3c :
		TR_210 = TR_67 ;
	7'h3d :
		TR_210 = TR_67 ;
	7'h3e :
		TR_210 = TR_67 ;
	7'h3f :
		TR_210 = TR_67 ;
	7'h40 :
		TR_210 = TR_67 ;
	7'h41 :
		TR_210 = TR_67 ;
	7'h42 :
		TR_210 = TR_67 ;
	7'h43 :
		TR_210 = TR_67 ;
	7'h44 :
		TR_210 = TR_67 ;
	7'h45 :
		TR_210 = TR_67 ;
	7'h46 :
		TR_210 = TR_67 ;
	7'h47 :
		TR_210 = TR_67 ;
	7'h48 :
		TR_210 = TR_67 ;
	7'h49 :
		TR_210 = TR_67 ;
	7'h4a :
		TR_210 = TR_67 ;
	7'h4b :
		TR_210 = TR_67 ;
	7'h4c :
		TR_210 = TR_67 ;
	7'h4d :
		TR_210 = TR_67 ;
	7'h4e :
		TR_210 = TR_67 ;
	7'h4f :
		TR_210 = TR_67 ;
	7'h50 :
		TR_210 = TR_67 ;
	7'h51 :
		TR_210 = TR_67 ;
	7'h52 :
		TR_210 = TR_67 ;
	7'h53 :
		TR_210 = TR_67 ;
	7'h54 :
		TR_210 = TR_67 ;
	7'h55 :
		TR_210 = TR_67 ;
	7'h56 :
		TR_210 = TR_67 ;
	7'h57 :
		TR_210 = TR_67 ;
	7'h58 :
		TR_210 = TR_67 ;
	7'h59 :
		TR_210 = TR_67 ;
	7'h5a :
		TR_210 = TR_67 ;
	7'h5b :
		TR_210 = TR_67 ;
	7'h5c :
		TR_210 = TR_67 ;
	7'h5d :
		TR_210 = TR_67 ;
	7'h5e :
		TR_210 = TR_67 ;
	7'h5f :
		TR_210 = TR_67 ;
	7'h60 :
		TR_210 = TR_67 ;
	7'h61 :
		TR_210 = TR_67 ;
	7'h62 :
		TR_210 = TR_67 ;
	7'h63 :
		TR_210 = TR_67 ;
	7'h64 :
		TR_210 = TR_67 ;
	7'h65 :
		TR_210 = TR_67 ;
	7'h66 :
		TR_210 = TR_67 ;
	7'h67 :
		TR_210 = TR_67 ;
	7'h68 :
		TR_210 = TR_67 ;
	7'h69 :
		TR_210 = TR_67 ;
	7'h6a :
		TR_210 = TR_67 ;
	7'h6b :
		TR_210 = TR_67 ;
	7'h6c :
		TR_210 = TR_67 ;
	7'h6d :
		TR_210 = TR_67 ;
	7'h6e :
		TR_210 = TR_67 ;
	7'h6f :
		TR_210 = TR_67 ;
	7'h70 :
		TR_210 = TR_67 ;
	7'h71 :
		TR_210 = TR_67 ;
	7'h72 :
		TR_210 = TR_67 ;
	7'h73 :
		TR_210 = TR_67 ;
	7'h74 :
		TR_210 = TR_67 ;
	7'h75 :
		TR_210 = TR_67 ;
	7'h76 :
		TR_210 = TR_67 ;
	7'h77 :
		TR_210 = TR_67 ;
	7'h78 :
		TR_210 = TR_67 ;
	7'h79 :
		TR_210 = TR_67 ;
	7'h7a :
		TR_210 = TR_67 ;
	7'h7b :
		TR_210 = TR_67 ;
	7'h7c :
		TR_210 = TR_67 ;
	7'h7d :
		TR_210 = TR_67 ;
	7'h7e :
		TR_210 = TR_67 ;
	7'h7f :
		TR_210 = TR_67 ;
	default :
		TR_210 = 9'hx ;
	endcase
always @ ( TR_210 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_25 or 
	U_174 or RG_rl_156 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_55_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h37 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_55_t = ( ( { 9{ ST1_03d } } & RG_rl_156 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_25 )
		| ( { 9{ U_173 } } & TR_210 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_55_en = ( ST1_03d | U_174 | RG_rl_55_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_55_en )
		RG_rl_55 <= RG_rl_55_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_68 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_209 = TR_68 ;
	7'h01 :
		TR_209 = TR_68 ;
	7'h02 :
		TR_209 = TR_68 ;
	7'h03 :
		TR_209 = TR_68 ;
	7'h04 :
		TR_209 = TR_68 ;
	7'h05 :
		TR_209 = TR_68 ;
	7'h06 :
		TR_209 = TR_68 ;
	7'h07 :
		TR_209 = TR_68 ;
	7'h08 :
		TR_209 = TR_68 ;
	7'h09 :
		TR_209 = TR_68 ;
	7'h0a :
		TR_209 = TR_68 ;
	7'h0b :
		TR_209 = TR_68 ;
	7'h0c :
		TR_209 = TR_68 ;
	7'h0d :
		TR_209 = TR_68 ;
	7'h0e :
		TR_209 = TR_68 ;
	7'h0f :
		TR_209 = TR_68 ;
	7'h10 :
		TR_209 = TR_68 ;
	7'h11 :
		TR_209 = TR_68 ;
	7'h12 :
		TR_209 = TR_68 ;
	7'h13 :
		TR_209 = TR_68 ;
	7'h14 :
		TR_209 = TR_68 ;
	7'h15 :
		TR_209 = TR_68 ;
	7'h16 :
		TR_209 = TR_68 ;
	7'h17 :
		TR_209 = TR_68 ;
	7'h18 :
		TR_209 = TR_68 ;
	7'h19 :
		TR_209 = TR_68 ;
	7'h1a :
		TR_209 = TR_68 ;
	7'h1b :
		TR_209 = TR_68 ;
	7'h1c :
		TR_209 = TR_68 ;
	7'h1d :
		TR_209 = TR_68 ;
	7'h1e :
		TR_209 = TR_68 ;
	7'h1f :
		TR_209 = TR_68 ;
	7'h20 :
		TR_209 = TR_68 ;
	7'h21 :
		TR_209 = TR_68 ;
	7'h22 :
		TR_209 = TR_68 ;
	7'h23 :
		TR_209 = TR_68 ;
	7'h24 :
		TR_209 = TR_68 ;
	7'h25 :
		TR_209 = TR_68 ;
	7'h26 :
		TR_209 = TR_68 ;
	7'h27 :
		TR_209 = TR_68 ;
	7'h28 :
		TR_209 = TR_68 ;
	7'h29 :
		TR_209 = TR_68 ;
	7'h2a :
		TR_209 = TR_68 ;
	7'h2b :
		TR_209 = TR_68 ;
	7'h2c :
		TR_209 = TR_68 ;
	7'h2d :
		TR_209 = TR_68 ;
	7'h2e :
		TR_209 = TR_68 ;
	7'h2f :
		TR_209 = TR_68 ;
	7'h30 :
		TR_209 = TR_68 ;
	7'h31 :
		TR_209 = TR_68 ;
	7'h32 :
		TR_209 = TR_68 ;
	7'h33 :
		TR_209 = TR_68 ;
	7'h34 :
		TR_209 = TR_68 ;
	7'h35 :
		TR_209 = TR_68 ;
	7'h36 :
		TR_209 = TR_68 ;
	7'h37 :
		TR_209 = TR_68 ;
	7'h38 :
		TR_209 = 9'h000 ;	// line#=../rle.cpp:80
	7'h39 :
		TR_209 = TR_68 ;
	7'h3a :
		TR_209 = TR_68 ;
	7'h3b :
		TR_209 = TR_68 ;
	7'h3c :
		TR_209 = TR_68 ;
	7'h3d :
		TR_209 = TR_68 ;
	7'h3e :
		TR_209 = TR_68 ;
	7'h3f :
		TR_209 = TR_68 ;
	7'h40 :
		TR_209 = TR_68 ;
	7'h41 :
		TR_209 = TR_68 ;
	7'h42 :
		TR_209 = TR_68 ;
	7'h43 :
		TR_209 = TR_68 ;
	7'h44 :
		TR_209 = TR_68 ;
	7'h45 :
		TR_209 = TR_68 ;
	7'h46 :
		TR_209 = TR_68 ;
	7'h47 :
		TR_209 = TR_68 ;
	7'h48 :
		TR_209 = TR_68 ;
	7'h49 :
		TR_209 = TR_68 ;
	7'h4a :
		TR_209 = TR_68 ;
	7'h4b :
		TR_209 = TR_68 ;
	7'h4c :
		TR_209 = TR_68 ;
	7'h4d :
		TR_209 = TR_68 ;
	7'h4e :
		TR_209 = TR_68 ;
	7'h4f :
		TR_209 = TR_68 ;
	7'h50 :
		TR_209 = TR_68 ;
	7'h51 :
		TR_209 = TR_68 ;
	7'h52 :
		TR_209 = TR_68 ;
	7'h53 :
		TR_209 = TR_68 ;
	7'h54 :
		TR_209 = TR_68 ;
	7'h55 :
		TR_209 = TR_68 ;
	7'h56 :
		TR_209 = TR_68 ;
	7'h57 :
		TR_209 = TR_68 ;
	7'h58 :
		TR_209 = TR_68 ;
	7'h59 :
		TR_209 = TR_68 ;
	7'h5a :
		TR_209 = TR_68 ;
	7'h5b :
		TR_209 = TR_68 ;
	7'h5c :
		TR_209 = TR_68 ;
	7'h5d :
		TR_209 = TR_68 ;
	7'h5e :
		TR_209 = TR_68 ;
	7'h5f :
		TR_209 = TR_68 ;
	7'h60 :
		TR_209 = TR_68 ;
	7'h61 :
		TR_209 = TR_68 ;
	7'h62 :
		TR_209 = TR_68 ;
	7'h63 :
		TR_209 = TR_68 ;
	7'h64 :
		TR_209 = TR_68 ;
	7'h65 :
		TR_209 = TR_68 ;
	7'h66 :
		TR_209 = TR_68 ;
	7'h67 :
		TR_209 = TR_68 ;
	7'h68 :
		TR_209 = TR_68 ;
	7'h69 :
		TR_209 = TR_68 ;
	7'h6a :
		TR_209 = TR_68 ;
	7'h6b :
		TR_209 = TR_68 ;
	7'h6c :
		TR_209 = TR_68 ;
	7'h6d :
		TR_209 = TR_68 ;
	7'h6e :
		TR_209 = TR_68 ;
	7'h6f :
		TR_209 = TR_68 ;
	7'h70 :
		TR_209 = TR_68 ;
	7'h71 :
		TR_209 = TR_68 ;
	7'h72 :
		TR_209 = TR_68 ;
	7'h73 :
		TR_209 = TR_68 ;
	7'h74 :
		TR_209 = TR_68 ;
	7'h75 :
		TR_209 = TR_68 ;
	7'h76 :
		TR_209 = TR_68 ;
	7'h77 :
		TR_209 = TR_68 ;
	7'h78 :
		TR_209 = TR_68 ;
	7'h79 :
		TR_209 = TR_68 ;
	7'h7a :
		TR_209 = TR_68 ;
	7'h7b :
		TR_209 = TR_68 ;
	7'h7c :
		TR_209 = TR_68 ;
	7'h7d :
		TR_209 = TR_68 ;
	7'h7e :
		TR_209 = TR_68 ;
	7'h7f :
		TR_209 = TR_68 ;
	default :
		TR_209 = 9'hx ;
	endcase
always @ ( TR_209 or U_173 or sub8u_71ot or U_183 or RG_rl_157 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_56_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h38 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_56_t = ( ( { 9{ M_180 } } & RG_rl_157 )
		| ( { 9{ U_173 } } & TR_209 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_56_en = ( M_180 | RG_rl_56_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_56_en )
		RG_rl_56 <= RG_rl_56_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_69 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_208 = TR_69 ;
	7'h01 :
		TR_208 = TR_69 ;
	7'h02 :
		TR_208 = TR_69 ;
	7'h03 :
		TR_208 = TR_69 ;
	7'h04 :
		TR_208 = TR_69 ;
	7'h05 :
		TR_208 = TR_69 ;
	7'h06 :
		TR_208 = TR_69 ;
	7'h07 :
		TR_208 = TR_69 ;
	7'h08 :
		TR_208 = TR_69 ;
	7'h09 :
		TR_208 = TR_69 ;
	7'h0a :
		TR_208 = TR_69 ;
	7'h0b :
		TR_208 = TR_69 ;
	7'h0c :
		TR_208 = TR_69 ;
	7'h0d :
		TR_208 = TR_69 ;
	7'h0e :
		TR_208 = TR_69 ;
	7'h0f :
		TR_208 = TR_69 ;
	7'h10 :
		TR_208 = TR_69 ;
	7'h11 :
		TR_208 = TR_69 ;
	7'h12 :
		TR_208 = TR_69 ;
	7'h13 :
		TR_208 = TR_69 ;
	7'h14 :
		TR_208 = TR_69 ;
	7'h15 :
		TR_208 = TR_69 ;
	7'h16 :
		TR_208 = TR_69 ;
	7'h17 :
		TR_208 = TR_69 ;
	7'h18 :
		TR_208 = TR_69 ;
	7'h19 :
		TR_208 = TR_69 ;
	7'h1a :
		TR_208 = TR_69 ;
	7'h1b :
		TR_208 = TR_69 ;
	7'h1c :
		TR_208 = TR_69 ;
	7'h1d :
		TR_208 = TR_69 ;
	7'h1e :
		TR_208 = TR_69 ;
	7'h1f :
		TR_208 = TR_69 ;
	7'h20 :
		TR_208 = TR_69 ;
	7'h21 :
		TR_208 = TR_69 ;
	7'h22 :
		TR_208 = TR_69 ;
	7'h23 :
		TR_208 = TR_69 ;
	7'h24 :
		TR_208 = TR_69 ;
	7'h25 :
		TR_208 = TR_69 ;
	7'h26 :
		TR_208 = TR_69 ;
	7'h27 :
		TR_208 = TR_69 ;
	7'h28 :
		TR_208 = TR_69 ;
	7'h29 :
		TR_208 = TR_69 ;
	7'h2a :
		TR_208 = TR_69 ;
	7'h2b :
		TR_208 = TR_69 ;
	7'h2c :
		TR_208 = TR_69 ;
	7'h2d :
		TR_208 = TR_69 ;
	7'h2e :
		TR_208 = TR_69 ;
	7'h2f :
		TR_208 = TR_69 ;
	7'h30 :
		TR_208 = TR_69 ;
	7'h31 :
		TR_208 = TR_69 ;
	7'h32 :
		TR_208 = TR_69 ;
	7'h33 :
		TR_208 = TR_69 ;
	7'h34 :
		TR_208 = TR_69 ;
	7'h35 :
		TR_208 = TR_69 ;
	7'h36 :
		TR_208 = TR_69 ;
	7'h37 :
		TR_208 = TR_69 ;
	7'h38 :
		TR_208 = TR_69 ;
	7'h39 :
		TR_208 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3a :
		TR_208 = TR_69 ;
	7'h3b :
		TR_208 = TR_69 ;
	7'h3c :
		TR_208 = TR_69 ;
	7'h3d :
		TR_208 = TR_69 ;
	7'h3e :
		TR_208 = TR_69 ;
	7'h3f :
		TR_208 = TR_69 ;
	7'h40 :
		TR_208 = TR_69 ;
	7'h41 :
		TR_208 = TR_69 ;
	7'h42 :
		TR_208 = TR_69 ;
	7'h43 :
		TR_208 = TR_69 ;
	7'h44 :
		TR_208 = TR_69 ;
	7'h45 :
		TR_208 = TR_69 ;
	7'h46 :
		TR_208 = TR_69 ;
	7'h47 :
		TR_208 = TR_69 ;
	7'h48 :
		TR_208 = TR_69 ;
	7'h49 :
		TR_208 = TR_69 ;
	7'h4a :
		TR_208 = TR_69 ;
	7'h4b :
		TR_208 = TR_69 ;
	7'h4c :
		TR_208 = TR_69 ;
	7'h4d :
		TR_208 = TR_69 ;
	7'h4e :
		TR_208 = TR_69 ;
	7'h4f :
		TR_208 = TR_69 ;
	7'h50 :
		TR_208 = TR_69 ;
	7'h51 :
		TR_208 = TR_69 ;
	7'h52 :
		TR_208 = TR_69 ;
	7'h53 :
		TR_208 = TR_69 ;
	7'h54 :
		TR_208 = TR_69 ;
	7'h55 :
		TR_208 = TR_69 ;
	7'h56 :
		TR_208 = TR_69 ;
	7'h57 :
		TR_208 = TR_69 ;
	7'h58 :
		TR_208 = TR_69 ;
	7'h59 :
		TR_208 = TR_69 ;
	7'h5a :
		TR_208 = TR_69 ;
	7'h5b :
		TR_208 = TR_69 ;
	7'h5c :
		TR_208 = TR_69 ;
	7'h5d :
		TR_208 = TR_69 ;
	7'h5e :
		TR_208 = TR_69 ;
	7'h5f :
		TR_208 = TR_69 ;
	7'h60 :
		TR_208 = TR_69 ;
	7'h61 :
		TR_208 = TR_69 ;
	7'h62 :
		TR_208 = TR_69 ;
	7'h63 :
		TR_208 = TR_69 ;
	7'h64 :
		TR_208 = TR_69 ;
	7'h65 :
		TR_208 = TR_69 ;
	7'h66 :
		TR_208 = TR_69 ;
	7'h67 :
		TR_208 = TR_69 ;
	7'h68 :
		TR_208 = TR_69 ;
	7'h69 :
		TR_208 = TR_69 ;
	7'h6a :
		TR_208 = TR_69 ;
	7'h6b :
		TR_208 = TR_69 ;
	7'h6c :
		TR_208 = TR_69 ;
	7'h6d :
		TR_208 = TR_69 ;
	7'h6e :
		TR_208 = TR_69 ;
	7'h6f :
		TR_208 = TR_69 ;
	7'h70 :
		TR_208 = TR_69 ;
	7'h71 :
		TR_208 = TR_69 ;
	7'h72 :
		TR_208 = TR_69 ;
	7'h73 :
		TR_208 = TR_69 ;
	7'h74 :
		TR_208 = TR_69 ;
	7'h75 :
		TR_208 = TR_69 ;
	7'h76 :
		TR_208 = TR_69 ;
	7'h77 :
		TR_208 = TR_69 ;
	7'h78 :
		TR_208 = TR_69 ;
	7'h79 :
		TR_208 = TR_69 ;
	7'h7a :
		TR_208 = TR_69 ;
	7'h7b :
		TR_208 = TR_69 ;
	7'h7c :
		TR_208 = TR_69 ;
	7'h7d :
		TR_208 = TR_69 ;
	7'h7e :
		TR_208 = TR_69 ;
	7'h7f :
		TR_208 = TR_69 ;
	default :
		TR_208 = 9'hx ;
	endcase
always @ ( TR_208 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_26 or 
	U_174 or RG_rl_157 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_57_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h39 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_57_t = ( ( { 9{ ST1_03d } } & RG_rl_157 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_26 )
		| ( { 9{ U_173 } } & TR_208 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_57_en = ( ST1_03d | U_174 | RG_rl_57_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_57_en )
		RG_rl_57 <= RG_rl_57_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_70 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_207 = TR_70 ;
	7'h01 :
		TR_207 = TR_70 ;
	7'h02 :
		TR_207 = TR_70 ;
	7'h03 :
		TR_207 = TR_70 ;
	7'h04 :
		TR_207 = TR_70 ;
	7'h05 :
		TR_207 = TR_70 ;
	7'h06 :
		TR_207 = TR_70 ;
	7'h07 :
		TR_207 = TR_70 ;
	7'h08 :
		TR_207 = TR_70 ;
	7'h09 :
		TR_207 = TR_70 ;
	7'h0a :
		TR_207 = TR_70 ;
	7'h0b :
		TR_207 = TR_70 ;
	7'h0c :
		TR_207 = TR_70 ;
	7'h0d :
		TR_207 = TR_70 ;
	7'h0e :
		TR_207 = TR_70 ;
	7'h0f :
		TR_207 = TR_70 ;
	7'h10 :
		TR_207 = TR_70 ;
	7'h11 :
		TR_207 = TR_70 ;
	7'h12 :
		TR_207 = TR_70 ;
	7'h13 :
		TR_207 = TR_70 ;
	7'h14 :
		TR_207 = TR_70 ;
	7'h15 :
		TR_207 = TR_70 ;
	7'h16 :
		TR_207 = TR_70 ;
	7'h17 :
		TR_207 = TR_70 ;
	7'h18 :
		TR_207 = TR_70 ;
	7'h19 :
		TR_207 = TR_70 ;
	7'h1a :
		TR_207 = TR_70 ;
	7'h1b :
		TR_207 = TR_70 ;
	7'h1c :
		TR_207 = TR_70 ;
	7'h1d :
		TR_207 = TR_70 ;
	7'h1e :
		TR_207 = TR_70 ;
	7'h1f :
		TR_207 = TR_70 ;
	7'h20 :
		TR_207 = TR_70 ;
	7'h21 :
		TR_207 = TR_70 ;
	7'h22 :
		TR_207 = TR_70 ;
	7'h23 :
		TR_207 = TR_70 ;
	7'h24 :
		TR_207 = TR_70 ;
	7'h25 :
		TR_207 = TR_70 ;
	7'h26 :
		TR_207 = TR_70 ;
	7'h27 :
		TR_207 = TR_70 ;
	7'h28 :
		TR_207 = TR_70 ;
	7'h29 :
		TR_207 = TR_70 ;
	7'h2a :
		TR_207 = TR_70 ;
	7'h2b :
		TR_207 = TR_70 ;
	7'h2c :
		TR_207 = TR_70 ;
	7'h2d :
		TR_207 = TR_70 ;
	7'h2e :
		TR_207 = TR_70 ;
	7'h2f :
		TR_207 = TR_70 ;
	7'h30 :
		TR_207 = TR_70 ;
	7'h31 :
		TR_207 = TR_70 ;
	7'h32 :
		TR_207 = TR_70 ;
	7'h33 :
		TR_207 = TR_70 ;
	7'h34 :
		TR_207 = TR_70 ;
	7'h35 :
		TR_207 = TR_70 ;
	7'h36 :
		TR_207 = TR_70 ;
	7'h37 :
		TR_207 = TR_70 ;
	7'h38 :
		TR_207 = TR_70 ;
	7'h39 :
		TR_207 = TR_70 ;
	7'h3a :
		TR_207 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3b :
		TR_207 = TR_70 ;
	7'h3c :
		TR_207 = TR_70 ;
	7'h3d :
		TR_207 = TR_70 ;
	7'h3e :
		TR_207 = TR_70 ;
	7'h3f :
		TR_207 = TR_70 ;
	7'h40 :
		TR_207 = TR_70 ;
	7'h41 :
		TR_207 = TR_70 ;
	7'h42 :
		TR_207 = TR_70 ;
	7'h43 :
		TR_207 = TR_70 ;
	7'h44 :
		TR_207 = TR_70 ;
	7'h45 :
		TR_207 = TR_70 ;
	7'h46 :
		TR_207 = TR_70 ;
	7'h47 :
		TR_207 = TR_70 ;
	7'h48 :
		TR_207 = TR_70 ;
	7'h49 :
		TR_207 = TR_70 ;
	7'h4a :
		TR_207 = TR_70 ;
	7'h4b :
		TR_207 = TR_70 ;
	7'h4c :
		TR_207 = TR_70 ;
	7'h4d :
		TR_207 = TR_70 ;
	7'h4e :
		TR_207 = TR_70 ;
	7'h4f :
		TR_207 = TR_70 ;
	7'h50 :
		TR_207 = TR_70 ;
	7'h51 :
		TR_207 = TR_70 ;
	7'h52 :
		TR_207 = TR_70 ;
	7'h53 :
		TR_207 = TR_70 ;
	7'h54 :
		TR_207 = TR_70 ;
	7'h55 :
		TR_207 = TR_70 ;
	7'h56 :
		TR_207 = TR_70 ;
	7'h57 :
		TR_207 = TR_70 ;
	7'h58 :
		TR_207 = TR_70 ;
	7'h59 :
		TR_207 = TR_70 ;
	7'h5a :
		TR_207 = TR_70 ;
	7'h5b :
		TR_207 = TR_70 ;
	7'h5c :
		TR_207 = TR_70 ;
	7'h5d :
		TR_207 = TR_70 ;
	7'h5e :
		TR_207 = TR_70 ;
	7'h5f :
		TR_207 = TR_70 ;
	7'h60 :
		TR_207 = TR_70 ;
	7'h61 :
		TR_207 = TR_70 ;
	7'h62 :
		TR_207 = TR_70 ;
	7'h63 :
		TR_207 = TR_70 ;
	7'h64 :
		TR_207 = TR_70 ;
	7'h65 :
		TR_207 = TR_70 ;
	7'h66 :
		TR_207 = TR_70 ;
	7'h67 :
		TR_207 = TR_70 ;
	7'h68 :
		TR_207 = TR_70 ;
	7'h69 :
		TR_207 = TR_70 ;
	7'h6a :
		TR_207 = TR_70 ;
	7'h6b :
		TR_207 = TR_70 ;
	7'h6c :
		TR_207 = TR_70 ;
	7'h6d :
		TR_207 = TR_70 ;
	7'h6e :
		TR_207 = TR_70 ;
	7'h6f :
		TR_207 = TR_70 ;
	7'h70 :
		TR_207 = TR_70 ;
	7'h71 :
		TR_207 = TR_70 ;
	7'h72 :
		TR_207 = TR_70 ;
	7'h73 :
		TR_207 = TR_70 ;
	7'h74 :
		TR_207 = TR_70 ;
	7'h75 :
		TR_207 = TR_70 ;
	7'h76 :
		TR_207 = TR_70 ;
	7'h77 :
		TR_207 = TR_70 ;
	7'h78 :
		TR_207 = TR_70 ;
	7'h79 :
		TR_207 = TR_70 ;
	7'h7a :
		TR_207 = TR_70 ;
	7'h7b :
		TR_207 = TR_70 ;
	7'h7c :
		TR_207 = TR_70 ;
	7'h7d :
		TR_207 = TR_70 ;
	7'h7e :
		TR_207 = TR_70 ;
	7'h7f :
		TR_207 = TR_70 ;
	default :
		TR_207 = 9'hx ;
	endcase
always @ ( TR_207 or U_173 or sub8u_71ot or U_183 or RG_rl_158 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_58_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h3a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_58_t = ( ( { 9{ M_180 } } & RG_rl_158 )
		| ( { 9{ U_173 } } & TR_207 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_58_en = ( M_180 | RG_rl_58_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_58_en )
		RG_rl_58 <= RG_rl_58_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_71 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_206 = TR_71 ;
	7'h01 :
		TR_206 = TR_71 ;
	7'h02 :
		TR_206 = TR_71 ;
	7'h03 :
		TR_206 = TR_71 ;
	7'h04 :
		TR_206 = TR_71 ;
	7'h05 :
		TR_206 = TR_71 ;
	7'h06 :
		TR_206 = TR_71 ;
	7'h07 :
		TR_206 = TR_71 ;
	7'h08 :
		TR_206 = TR_71 ;
	7'h09 :
		TR_206 = TR_71 ;
	7'h0a :
		TR_206 = TR_71 ;
	7'h0b :
		TR_206 = TR_71 ;
	7'h0c :
		TR_206 = TR_71 ;
	7'h0d :
		TR_206 = TR_71 ;
	7'h0e :
		TR_206 = TR_71 ;
	7'h0f :
		TR_206 = TR_71 ;
	7'h10 :
		TR_206 = TR_71 ;
	7'h11 :
		TR_206 = TR_71 ;
	7'h12 :
		TR_206 = TR_71 ;
	7'h13 :
		TR_206 = TR_71 ;
	7'h14 :
		TR_206 = TR_71 ;
	7'h15 :
		TR_206 = TR_71 ;
	7'h16 :
		TR_206 = TR_71 ;
	7'h17 :
		TR_206 = TR_71 ;
	7'h18 :
		TR_206 = TR_71 ;
	7'h19 :
		TR_206 = TR_71 ;
	7'h1a :
		TR_206 = TR_71 ;
	7'h1b :
		TR_206 = TR_71 ;
	7'h1c :
		TR_206 = TR_71 ;
	7'h1d :
		TR_206 = TR_71 ;
	7'h1e :
		TR_206 = TR_71 ;
	7'h1f :
		TR_206 = TR_71 ;
	7'h20 :
		TR_206 = TR_71 ;
	7'h21 :
		TR_206 = TR_71 ;
	7'h22 :
		TR_206 = TR_71 ;
	7'h23 :
		TR_206 = TR_71 ;
	7'h24 :
		TR_206 = TR_71 ;
	7'h25 :
		TR_206 = TR_71 ;
	7'h26 :
		TR_206 = TR_71 ;
	7'h27 :
		TR_206 = TR_71 ;
	7'h28 :
		TR_206 = TR_71 ;
	7'h29 :
		TR_206 = TR_71 ;
	7'h2a :
		TR_206 = TR_71 ;
	7'h2b :
		TR_206 = TR_71 ;
	7'h2c :
		TR_206 = TR_71 ;
	7'h2d :
		TR_206 = TR_71 ;
	7'h2e :
		TR_206 = TR_71 ;
	7'h2f :
		TR_206 = TR_71 ;
	7'h30 :
		TR_206 = TR_71 ;
	7'h31 :
		TR_206 = TR_71 ;
	7'h32 :
		TR_206 = TR_71 ;
	7'h33 :
		TR_206 = TR_71 ;
	7'h34 :
		TR_206 = TR_71 ;
	7'h35 :
		TR_206 = TR_71 ;
	7'h36 :
		TR_206 = TR_71 ;
	7'h37 :
		TR_206 = TR_71 ;
	7'h38 :
		TR_206 = TR_71 ;
	7'h39 :
		TR_206 = TR_71 ;
	7'h3a :
		TR_206 = TR_71 ;
	7'h3b :
		TR_206 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3c :
		TR_206 = TR_71 ;
	7'h3d :
		TR_206 = TR_71 ;
	7'h3e :
		TR_206 = TR_71 ;
	7'h3f :
		TR_206 = TR_71 ;
	7'h40 :
		TR_206 = TR_71 ;
	7'h41 :
		TR_206 = TR_71 ;
	7'h42 :
		TR_206 = TR_71 ;
	7'h43 :
		TR_206 = TR_71 ;
	7'h44 :
		TR_206 = TR_71 ;
	7'h45 :
		TR_206 = TR_71 ;
	7'h46 :
		TR_206 = TR_71 ;
	7'h47 :
		TR_206 = TR_71 ;
	7'h48 :
		TR_206 = TR_71 ;
	7'h49 :
		TR_206 = TR_71 ;
	7'h4a :
		TR_206 = TR_71 ;
	7'h4b :
		TR_206 = TR_71 ;
	7'h4c :
		TR_206 = TR_71 ;
	7'h4d :
		TR_206 = TR_71 ;
	7'h4e :
		TR_206 = TR_71 ;
	7'h4f :
		TR_206 = TR_71 ;
	7'h50 :
		TR_206 = TR_71 ;
	7'h51 :
		TR_206 = TR_71 ;
	7'h52 :
		TR_206 = TR_71 ;
	7'h53 :
		TR_206 = TR_71 ;
	7'h54 :
		TR_206 = TR_71 ;
	7'h55 :
		TR_206 = TR_71 ;
	7'h56 :
		TR_206 = TR_71 ;
	7'h57 :
		TR_206 = TR_71 ;
	7'h58 :
		TR_206 = TR_71 ;
	7'h59 :
		TR_206 = TR_71 ;
	7'h5a :
		TR_206 = TR_71 ;
	7'h5b :
		TR_206 = TR_71 ;
	7'h5c :
		TR_206 = TR_71 ;
	7'h5d :
		TR_206 = TR_71 ;
	7'h5e :
		TR_206 = TR_71 ;
	7'h5f :
		TR_206 = TR_71 ;
	7'h60 :
		TR_206 = TR_71 ;
	7'h61 :
		TR_206 = TR_71 ;
	7'h62 :
		TR_206 = TR_71 ;
	7'h63 :
		TR_206 = TR_71 ;
	7'h64 :
		TR_206 = TR_71 ;
	7'h65 :
		TR_206 = TR_71 ;
	7'h66 :
		TR_206 = TR_71 ;
	7'h67 :
		TR_206 = TR_71 ;
	7'h68 :
		TR_206 = TR_71 ;
	7'h69 :
		TR_206 = TR_71 ;
	7'h6a :
		TR_206 = TR_71 ;
	7'h6b :
		TR_206 = TR_71 ;
	7'h6c :
		TR_206 = TR_71 ;
	7'h6d :
		TR_206 = TR_71 ;
	7'h6e :
		TR_206 = TR_71 ;
	7'h6f :
		TR_206 = TR_71 ;
	7'h70 :
		TR_206 = TR_71 ;
	7'h71 :
		TR_206 = TR_71 ;
	7'h72 :
		TR_206 = TR_71 ;
	7'h73 :
		TR_206 = TR_71 ;
	7'h74 :
		TR_206 = TR_71 ;
	7'h75 :
		TR_206 = TR_71 ;
	7'h76 :
		TR_206 = TR_71 ;
	7'h77 :
		TR_206 = TR_71 ;
	7'h78 :
		TR_206 = TR_71 ;
	7'h79 :
		TR_206 = TR_71 ;
	7'h7a :
		TR_206 = TR_71 ;
	7'h7b :
		TR_206 = TR_71 ;
	7'h7c :
		TR_206 = TR_71 ;
	7'h7d :
		TR_206 = TR_71 ;
	7'h7e :
		TR_206 = TR_71 ;
	7'h7f :
		TR_206 = TR_71 ;
	default :
		TR_206 = 9'hx ;
	endcase
always @ ( TR_206 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_27 or 
	U_174 or RG_rl_158 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_59_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h3b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_59_t = ( ( { 9{ ST1_03d } } & RG_rl_158 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_27 )
		| ( { 9{ U_173 } } & TR_206 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_59_en = ( ST1_03d | U_174 | RG_rl_59_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_59_en )
		RG_rl_59 <= RG_rl_59_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_72 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_205 = TR_72 ;
	7'h01 :
		TR_205 = TR_72 ;
	7'h02 :
		TR_205 = TR_72 ;
	7'h03 :
		TR_205 = TR_72 ;
	7'h04 :
		TR_205 = TR_72 ;
	7'h05 :
		TR_205 = TR_72 ;
	7'h06 :
		TR_205 = TR_72 ;
	7'h07 :
		TR_205 = TR_72 ;
	7'h08 :
		TR_205 = TR_72 ;
	7'h09 :
		TR_205 = TR_72 ;
	7'h0a :
		TR_205 = TR_72 ;
	7'h0b :
		TR_205 = TR_72 ;
	7'h0c :
		TR_205 = TR_72 ;
	7'h0d :
		TR_205 = TR_72 ;
	7'h0e :
		TR_205 = TR_72 ;
	7'h0f :
		TR_205 = TR_72 ;
	7'h10 :
		TR_205 = TR_72 ;
	7'h11 :
		TR_205 = TR_72 ;
	7'h12 :
		TR_205 = TR_72 ;
	7'h13 :
		TR_205 = TR_72 ;
	7'h14 :
		TR_205 = TR_72 ;
	7'h15 :
		TR_205 = TR_72 ;
	7'h16 :
		TR_205 = TR_72 ;
	7'h17 :
		TR_205 = TR_72 ;
	7'h18 :
		TR_205 = TR_72 ;
	7'h19 :
		TR_205 = TR_72 ;
	7'h1a :
		TR_205 = TR_72 ;
	7'h1b :
		TR_205 = TR_72 ;
	7'h1c :
		TR_205 = TR_72 ;
	7'h1d :
		TR_205 = TR_72 ;
	7'h1e :
		TR_205 = TR_72 ;
	7'h1f :
		TR_205 = TR_72 ;
	7'h20 :
		TR_205 = TR_72 ;
	7'h21 :
		TR_205 = TR_72 ;
	7'h22 :
		TR_205 = TR_72 ;
	7'h23 :
		TR_205 = TR_72 ;
	7'h24 :
		TR_205 = TR_72 ;
	7'h25 :
		TR_205 = TR_72 ;
	7'h26 :
		TR_205 = TR_72 ;
	7'h27 :
		TR_205 = TR_72 ;
	7'h28 :
		TR_205 = TR_72 ;
	7'h29 :
		TR_205 = TR_72 ;
	7'h2a :
		TR_205 = TR_72 ;
	7'h2b :
		TR_205 = TR_72 ;
	7'h2c :
		TR_205 = TR_72 ;
	7'h2d :
		TR_205 = TR_72 ;
	7'h2e :
		TR_205 = TR_72 ;
	7'h2f :
		TR_205 = TR_72 ;
	7'h30 :
		TR_205 = TR_72 ;
	7'h31 :
		TR_205 = TR_72 ;
	7'h32 :
		TR_205 = TR_72 ;
	7'h33 :
		TR_205 = TR_72 ;
	7'h34 :
		TR_205 = TR_72 ;
	7'h35 :
		TR_205 = TR_72 ;
	7'h36 :
		TR_205 = TR_72 ;
	7'h37 :
		TR_205 = TR_72 ;
	7'h38 :
		TR_205 = TR_72 ;
	7'h39 :
		TR_205 = TR_72 ;
	7'h3a :
		TR_205 = TR_72 ;
	7'h3b :
		TR_205 = TR_72 ;
	7'h3c :
		TR_205 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3d :
		TR_205 = TR_72 ;
	7'h3e :
		TR_205 = TR_72 ;
	7'h3f :
		TR_205 = TR_72 ;
	7'h40 :
		TR_205 = TR_72 ;
	7'h41 :
		TR_205 = TR_72 ;
	7'h42 :
		TR_205 = TR_72 ;
	7'h43 :
		TR_205 = TR_72 ;
	7'h44 :
		TR_205 = TR_72 ;
	7'h45 :
		TR_205 = TR_72 ;
	7'h46 :
		TR_205 = TR_72 ;
	7'h47 :
		TR_205 = TR_72 ;
	7'h48 :
		TR_205 = TR_72 ;
	7'h49 :
		TR_205 = TR_72 ;
	7'h4a :
		TR_205 = TR_72 ;
	7'h4b :
		TR_205 = TR_72 ;
	7'h4c :
		TR_205 = TR_72 ;
	7'h4d :
		TR_205 = TR_72 ;
	7'h4e :
		TR_205 = TR_72 ;
	7'h4f :
		TR_205 = TR_72 ;
	7'h50 :
		TR_205 = TR_72 ;
	7'h51 :
		TR_205 = TR_72 ;
	7'h52 :
		TR_205 = TR_72 ;
	7'h53 :
		TR_205 = TR_72 ;
	7'h54 :
		TR_205 = TR_72 ;
	7'h55 :
		TR_205 = TR_72 ;
	7'h56 :
		TR_205 = TR_72 ;
	7'h57 :
		TR_205 = TR_72 ;
	7'h58 :
		TR_205 = TR_72 ;
	7'h59 :
		TR_205 = TR_72 ;
	7'h5a :
		TR_205 = TR_72 ;
	7'h5b :
		TR_205 = TR_72 ;
	7'h5c :
		TR_205 = TR_72 ;
	7'h5d :
		TR_205 = TR_72 ;
	7'h5e :
		TR_205 = TR_72 ;
	7'h5f :
		TR_205 = TR_72 ;
	7'h60 :
		TR_205 = TR_72 ;
	7'h61 :
		TR_205 = TR_72 ;
	7'h62 :
		TR_205 = TR_72 ;
	7'h63 :
		TR_205 = TR_72 ;
	7'h64 :
		TR_205 = TR_72 ;
	7'h65 :
		TR_205 = TR_72 ;
	7'h66 :
		TR_205 = TR_72 ;
	7'h67 :
		TR_205 = TR_72 ;
	7'h68 :
		TR_205 = TR_72 ;
	7'h69 :
		TR_205 = TR_72 ;
	7'h6a :
		TR_205 = TR_72 ;
	7'h6b :
		TR_205 = TR_72 ;
	7'h6c :
		TR_205 = TR_72 ;
	7'h6d :
		TR_205 = TR_72 ;
	7'h6e :
		TR_205 = TR_72 ;
	7'h6f :
		TR_205 = TR_72 ;
	7'h70 :
		TR_205 = TR_72 ;
	7'h71 :
		TR_205 = TR_72 ;
	7'h72 :
		TR_205 = TR_72 ;
	7'h73 :
		TR_205 = TR_72 ;
	7'h74 :
		TR_205 = TR_72 ;
	7'h75 :
		TR_205 = TR_72 ;
	7'h76 :
		TR_205 = TR_72 ;
	7'h77 :
		TR_205 = TR_72 ;
	7'h78 :
		TR_205 = TR_72 ;
	7'h79 :
		TR_205 = TR_72 ;
	7'h7a :
		TR_205 = TR_72 ;
	7'h7b :
		TR_205 = TR_72 ;
	7'h7c :
		TR_205 = TR_72 ;
	7'h7d :
		TR_205 = TR_72 ;
	7'h7e :
		TR_205 = TR_72 ;
	7'h7f :
		TR_205 = TR_72 ;
	default :
		TR_205 = 9'hx ;
	endcase
always @ ( TR_205 or U_173 or sub8u_71ot or U_183 or RG_rl_159 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_60_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h3c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_60_t = ( ( { 9{ M_180 } } & RG_rl_159 )
		| ( { 9{ U_173 } } & TR_205 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_60_en = ( M_180 | RG_rl_60_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_60_en )
		RG_rl_60 <= RG_rl_60_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_73 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_204 = TR_73 ;
	7'h01 :
		TR_204 = TR_73 ;
	7'h02 :
		TR_204 = TR_73 ;
	7'h03 :
		TR_204 = TR_73 ;
	7'h04 :
		TR_204 = TR_73 ;
	7'h05 :
		TR_204 = TR_73 ;
	7'h06 :
		TR_204 = TR_73 ;
	7'h07 :
		TR_204 = TR_73 ;
	7'h08 :
		TR_204 = TR_73 ;
	7'h09 :
		TR_204 = TR_73 ;
	7'h0a :
		TR_204 = TR_73 ;
	7'h0b :
		TR_204 = TR_73 ;
	7'h0c :
		TR_204 = TR_73 ;
	7'h0d :
		TR_204 = TR_73 ;
	7'h0e :
		TR_204 = TR_73 ;
	7'h0f :
		TR_204 = TR_73 ;
	7'h10 :
		TR_204 = TR_73 ;
	7'h11 :
		TR_204 = TR_73 ;
	7'h12 :
		TR_204 = TR_73 ;
	7'h13 :
		TR_204 = TR_73 ;
	7'h14 :
		TR_204 = TR_73 ;
	7'h15 :
		TR_204 = TR_73 ;
	7'h16 :
		TR_204 = TR_73 ;
	7'h17 :
		TR_204 = TR_73 ;
	7'h18 :
		TR_204 = TR_73 ;
	7'h19 :
		TR_204 = TR_73 ;
	7'h1a :
		TR_204 = TR_73 ;
	7'h1b :
		TR_204 = TR_73 ;
	7'h1c :
		TR_204 = TR_73 ;
	7'h1d :
		TR_204 = TR_73 ;
	7'h1e :
		TR_204 = TR_73 ;
	7'h1f :
		TR_204 = TR_73 ;
	7'h20 :
		TR_204 = TR_73 ;
	7'h21 :
		TR_204 = TR_73 ;
	7'h22 :
		TR_204 = TR_73 ;
	7'h23 :
		TR_204 = TR_73 ;
	7'h24 :
		TR_204 = TR_73 ;
	7'h25 :
		TR_204 = TR_73 ;
	7'h26 :
		TR_204 = TR_73 ;
	7'h27 :
		TR_204 = TR_73 ;
	7'h28 :
		TR_204 = TR_73 ;
	7'h29 :
		TR_204 = TR_73 ;
	7'h2a :
		TR_204 = TR_73 ;
	7'h2b :
		TR_204 = TR_73 ;
	7'h2c :
		TR_204 = TR_73 ;
	7'h2d :
		TR_204 = TR_73 ;
	7'h2e :
		TR_204 = TR_73 ;
	7'h2f :
		TR_204 = TR_73 ;
	7'h30 :
		TR_204 = TR_73 ;
	7'h31 :
		TR_204 = TR_73 ;
	7'h32 :
		TR_204 = TR_73 ;
	7'h33 :
		TR_204 = TR_73 ;
	7'h34 :
		TR_204 = TR_73 ;
	7'h35 :
		TR_204 = TR_73 ;
	7'h36 :
		TR_204 = TR_73 ;
	7'h37 :
		TR_204 = TR_73 ;
	7'h38 :
		TR_204 = TR_73 ;
	7'h39 :
		TR_204 = TR_73 ;
	7'h3a :
		TR_204 = TR_73 ;
	7'h3b :
		TR_204 = TR_73 ;
	7'h3c :
		TR_204 = TR_73 ;
	7'h3d :
		TR_204 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3e :
		TR_204 = TR_73 ;
	7'h3f :
		TR_204 = TR_73 ;
	7'h40 :
		TR_204 = TR_73 ;
	7'h41 :
		TR_204 = TR_73 ;
	7'h42 :
		TR_204 = TR_73 ;
	7'h43 :
		TR_204 = TR_73 ;
	7'h44 :
		TR_204 = TR_73 ;
	7'h45 :
		TR_204 = TR_73 ;
	7'h46 :
		TR_204 = TR_73 ;
	7'h47 :
		TR_204 = TR_73 ;
	7'h48 :
		TR_204 = TR_73 ;
	7'h49 :
		TR_204 = TR_73 ;
	7'h4a :
		TR_204 = TR_73 ;
	7'h4b :
		TR_204 = TR_73 ;
	7'h4c :
		TR_204 = TR_73 ;
	7'h4d :
		TR_204 = TR_73 ;
	7'h4e :
		TR_204 = TR_73 ;
	7'h4f :
		TR_204 = TR_73 ;
	7'h50 :
		TR_204 = TR_73 ;
	7'h51 :
		TR_204 = TR_73 ;
	7'h52 :
		TR_204 = TR_73 ;
	7'h53 :
		TR_204 = TR_73 ;
	7'h54 :
		TR_204 = TR_73 ;
	7'h55 :
		TR_204 = TR_73 ;
	7'h56 :
		TR_204 = TR_73 ;
	7'h57 :
		TR_204 = TR_73 ;
	7'h58 :
		TR_204 = TR_73 ;
	7'h59 :
		TR_204 = TR_73 ;
	7'h5a :
		TR_204 = TR_73 ;
	7'h5b :
		TR_204 = TR_73 ;
	7'h5c :
		TR_204 = TR_73 ;
	7'h5d :
		TR_204 = TR_73 ;
	7'h5e :
		TR_204 = TR_73 ;
	7'h5f :
		TR_204 = TR_73 ;
	7'h60 :
		TR_204 = TR_73 ;
	7'h61 :
		TR_204 = TR_73 ;
	7'h62 :
		TR_204 = TR_73 ;
	7'h63 :
		TR_204 = TR_73 ;
	7'h64 :
		TR_204 = TR_73 ;
	7'h65 :
		TR_204 = TR_73 ;
	7'h66 :
		TR_204 = TR_73 ;
	7'h67 :
		TR_204 = TR_73 ;
	7'h68 :
		TR_204 = TR_73 ;
	7'h69 :
		TR_204 = TR_73 ;
	7'h6a :
		TR_204 = TR_73 ;
	7'h6b :
		TR_204 = TR_73 ;
	7'h6c :
		TR_204 = TR_73 ;
	7'h6d :
		TR_204 = TR_73 ;
	7'h6e :
		TR_204 = TR_73 ;
	7'h6f :
		TR_204 = TR_73 ;
	7'h70 :
		TR_204 = TR_73 ;
	7'h71 :
		TR_204 = TR_73 ;
	7'h72 :
		TR_204 = TR_73 ;
	7'h73 :
		TR_204 = TR_73 ;
	7'h74 :
		TR_204 = TR_73 ;
	7'h75 :
		TR_204 = TR_73 ;
	7'h76 :
		TR_204 = TR_73 ;
	7'h77 :
		TR_204 = TR_73 ;
	7'h78 :
		TR_204 = TR_73 ;
	7'h79 :
		TR_204 = TR_73 ;
	7'h7a :
		TR_204 = TR_73 ;
	7'h7b :
		TR_204 = TR_73 ;
	7'h7c :
		TR_204 = TR_73 ;
	7'h7d :
		TR_204 = TR_73 ;
	7'h7e :
		TR_204 = TR_73 ;
	7'h7f :
		TR_204 = TR_73 ;
	default :
		TR_204 = 9'hx ;
	endcase
always @ ( TR_204 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_28 or 
	U_174 or RG_rl_159 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_61_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h3d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_61_t = ( ( { 9{ ST1_03d } } & RG_rl_159 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_28 )
		| ( { 9{ U_173 } } & TR_204 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_61_en = ( ST1_03d | U_174 | RG_rl_61_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_61_en )
		RG_rl_61 <= RG_rl_61_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_74 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_203 = TR_74 ;
	7'h01 :
		TR_203 = TR_74 ;
	7'h02 :
		TR_203 = TR_74 ;
	7'h03 :
		TR_203 = TR_74 ;
	7'h04 :
		TR_203 = TR_74 ;
	7'h05 :
		TR_203 = TR_74 ;
	7'h06 :
		TR_203 = TR_74 ;
	7'h07 :
		TR_203 = TR_74 ;
	7'h08 :
		TR_203 = TR_74 ;
	7'h09 :
		TR_203 = TR_74 ;
	7'h0a :
		TR_203 = TR_74 ;
	7'h0b :
		TR_203 = TR_74 ;
	7'h0c :
		TR_203 = TR_74 ;
	7'h0d :
		TR_203 = TR_74 ;
	7'h0e :
		TR_203 = TR_74 ;
	7'h0f :
		TR_203 = TR_74 ;
	7'h10 :
		TR_203 = TR_74 ;
	7'h11 :
		TR_203 = TR_74 ;
	7'h12 :
		TR_203 = TR_74 ;
	7'h13 :
		TR_203 = TR_74 ;
	7'h14 :
		TR_203 = TR_74 ;
	7'h15 :
		TR_203 = TR_74 ;
	7'h16 :
		TR_203 = TR_74 ;
	7'h17 :
		TR_203 = TR_74 ;
	7'h18 :
		TR_203 = TR_74 ;
	7'h19 :
		TR_203 = TR_74 ;
	7'h1a :
		TR_203 = TR_74 ;
	7'h1b :
		TR_203 = TR_74 ;
	7'h1c :
		TR_203 = TR_74 ;
	7'h1d :
		TR_203 = TR_74 ;
	7'h1e :
		TR_203 = TR_74 ;
	7'h1f :
		TR_203 = TR_74 ;
	7'h20 :
		TR_203 = TR_74 ;
	7'h21 :
		TR_203 = TR_74 ;
	7'h22 :
		TR_203 = TR_74 ;
	7'h23 :
		TR_203 = TR_74 ;
	7'h24 :
		TR_203 = TR_74 ;
	7'h25 :
		TR_203 = TR_74 ;
	7'h26 :
		TR_203 = TR_74 ;
	7'h27 :
		TR_203 = TR_74 ;
	7'h28 :
		TR_203 = TR_74 ;
	7'h29 :
		TR_203 = TR_74 ;
	7'h2a :
		TR_203 = TR_74 ;
	7'h2b :
		TR_203 = TR_74 ;
	7'h2c :
		TR_203 = TR_74 ;
	7'h2d :
		TR_203 = TR_74 ;
	7'h2e :
		TR_203 = TR_74 ;
	7'h2f :
		TR_203 = TR_74 ;
	7'h30 :
		TR_203 = TR_74 ;
	7'h31 :
		TR_203 = TR_74 ;
	7'h32 :
		TR_203 = TR_74 ;
	7'h33 :
		TR_203 = TR_74 ;
	7'h34 :
		TR_203 = TR_74 ;
	7'h35 :
		TR_203 = TR_74 ;
	7'h36 :
		TR_203 = TR_74 ;
	7'h37 :
		TR_203 = TR_74 ;
	7'h38 :
		TR_203 = TR_74 ;
	7'h39 :
		TR_203 = TR_74 ;
	7'h3a :
		TR_203 = TR_74 ;
	7'h3b :
		TR_203 = TR_74 ;
	7'h3c :
		TR_203 = TR_74 ;
	7'h3d :
		TR_203 = TR_74 ;
	7'h3e :
		TR_203 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3f :
		TR_203 = TR_74 ;
	7'h40 :
		TR_203 = TR_74 ;
	7'h41 :
		TR_203 = TR_74 ;
	7'h42 :
		TR_203 = TR_74 ;
	7'h43 :
		TR_203 = TR_74 ;
	7'h44 :
		TR_203 = TR_74 ;
	7'h45 :
		TR_203 = TR_74 ;
	7'h46 :
		TR_203 = TR_74 ;
	7'h47 :
		TR_203 = TR_74 ;
	7'h48 :
		TR_203 = TR_74 ;
	7'h49 :
		TR_203 = TR_74 ;
	7'h4a :
		TR_203 = TR_74 ;
	7'h4b :
		TR_203 = TR_74 ;
	7'h4c :
		TR_203 = TR_74 ;
	7'h4d :
		TR_203 = TR_74 ;
	7'h4e :
		TR_203 = TR_74 ;
	7'h4f :
		TR_203 = TR_74 ;
	7'h50 :
		TR_203 = TR_74 ;
	7'h51 :
		TR_203 = TR_74 ;
	7'h52 :
		TR_203 = TR_74 ;
	7'h53 :
		TR_203 = TR_74 ;
	7'h54 :
		TR_203 = TR_74 ;
	7'h55 :
		TR_203 = TR_74 ;
	7'h56 :
		TR_203 = TR_74 ;
	7'h57 :
		TR_203 = TR_74 ;
	7'h58 :
		TR_203 = TR_74 ;
	7'h59 :
		TR_203 = TR_74 ;
	7'h5a :
		TR_203 = TR_74 ;
	7'h5b :
		TR_203 = TR_74 ;
	7'h5c :
		TR_203 = TR_74 ;
	7'h5d :
		TR_203 = TR_74 ;
	7'h5e :
		TR_203 = TR_74 ;
	7'h5f :
		TR_203 = TR_74 ;
	7'h60 :
		TR_203 = TR_74 ;
	7'h61 :
		TR_203 = TR_74 ;
	7'h62 :
		TR_203 = TR_74 ;
	7'h63 :
		TR_203 = TR_74 ;
	7'h64 :
		TR_203 = TR_74 ;
	7'h65 :
		TR_203 = TR_74 ;
	7'h66 :
		TR_203 = TR_74 ;
	7'h67 :
		TR_203 = TR_74 ;
	7'h68 :
		TR_203 = TR_74 ;
	7'h69 :
		TR_203 = TR_74 ;
	7'h6a :
		TR_203 = TR_74 ;
	7'h6b :
		TR_203 = TR_74 ;
	7'h6c :
		TR_203 = TR_74 ;
	7'h6d :
		TR_203 = TR_74 ;
	7'h6e :
		TR_203 = TR_74 ;
	7'h6f :
		TR_203 = TR_74 ;
	7'h70 :
		TR_203 = TR_74 ;
	7'h71 :
		TR_203 = TR_74 ;
	7'h72 :
		TR_203 = TR_74 ;
	7'h73 :
		TR_203 = TR_74 ;
	7'h74 :
		TR_203 = TR_74 ;
	7'h75 :
		TR_203 = TR_74 ;
	7'h76 :
		TR_203 = TR_74 ;
	7'h77 :
		TR_203 = TR_74 ;
	7'h78 :
		TR_203 = TR_74 ;
	7'h79 :
		TR_203 = TR_74 ;
	7'h7a :
		TR_203 = TR_74 ;
	7'h7b :
		TR_203 = TR_74 ;
	7'h7c :
		TR_203 = TR_74 ;
	7'h7d :
		TR_203 = TR_74 ;
	7'h7e :
		TR_203 = TR_74 ;
	7'h7f :
		TR_203 = TR_74 ;
	default :
		TR_203 = 9'hx ;
	endcase
always @ ( TR_203 or U_173 or sub8u_71ot or U_183 or RG_rl_160 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_62_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h3e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_62_t = ( ( { 9{ M_180 } } & RG_rl_160 )
		| ( { 9{ U_173 } } & TR_203 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_62_en = ( M_180 | RG_rl_62_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_62_en )
		RG_rl_62 <= RG_rl_62_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_75 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_202 = TR_75 ;
	7'h01 :
		TR_202 = TR_75 ;
	7'h02 :
		TR_202 = TR_75 ;
	7'h03 :
		TR_202 = TR_75 ;
	7'h04 :
		TR_202 = TR_75 ;
	7'h05 :
		TR_202 = TR_75 ;
	7'h06 :
		TR_202 = TR_75 ;
	7'h07 :
		TR_202 = TR_75 ;
	7'h08 :
		TR_202 = TR_75 ;
	7'h09 :
		TR_202 = TR_75 ;
	7'h0a :
		TR_202 = TR_75 ;
	7'h0b :
		TR_202 = TR_75 ;
	7'h0c :
		TR_202 = TR_75 ;
	7'h0d :
		TR_202 = TR_75 ;
	7'h0e :
		TR_202 = TR_75 ;
	7'h0f :
		TR_202 = TR_75 ;
	7'h10 :
		TR_202 = TR_75 ;
	7'h11 :
		TR_202 = TR_75 ;
	7'h12 :
		TR_202 = TR_75 ;
	7'h13 :
		TR_202 = TR_75 ;
	7'h14 :
		TR_202 = TR_75 ;
	7'h15 :
		TR_202 = TR_75 ;
	7'h16 :
		TR_202 = TR_75 ;
	7'h17 :
		TR_202 = TR_75 ;
	7'h18 :
		TR_202 = TR_75 ;
	7'h19 :
		TR_202 = TR_75 ;
	7'h1a :
		TR_202 = TR_75 ;
	7'h1b :
		TR_202 = TR_75 ;
	7'h1c :
		TR_202 = TR_75 ;
	7'h1d :
		TR_202 = TR_75 ;
	7'h1e :
		TR_202 = TR_75 ;
	7'h1f :
		TR_202 = TR_75 ;
	7'h20 :
		TR_202 = TR_75 ;
	7'h21 :
		TR_202 = TR_75 ;
	7'h22 :
		TR_202 = TR_75 ;
	7'h23 :
		TR_202 = TR_75 ;
	7'h24 :
		TR_202 = TR_75 ;
	7'h25 :
		TR_202 = TR_75 ;
	7'h26 :
		TR_202 = TR_75 ;
	7'h27 :
		TR_202 = TR_75 ;
	7'h28 :
		TR_202 = TR_75 ;
	7'h29 :
		TR_202 = TR_75 ;
	7'h2a :
		TR_202 = TR_75 ;
	7'h2b :
		TR_202 = TR_75 ;
	7'h2c :
		TR_202 = TR_75 ;
	7'h2d :
		TR_202 = TR_75 ;
	7'h2e :
		TR_202 = TR_75 ;
	7'h2f :
		TR_202 = TR_75 ;
	7'h30 :
		TR_202 = TR_75 ;
	7'h31 :
		TR_202 = TR_75 ;
	7'h32 :
		TR_202 = TR_75 ;
	7'h33 :
		TR_202 = TR_75 ;
	7'h34 :
		TR_202 = TR_75 ;
	7'h35 :
		TR_202 = TR_75 ;
	7'h36 :
		TR_202 = TR_75 ;
	7'h37 :
		TR_202 = TR_75 ;
	7'h38 :
		TR_202 = TR_75 ;
	7'h39 :
		TR_202 = TR_75 ;
	7'h3a :
		TR_202 = TR_75 ;
	7'h3b :
		TR_202 = TR_75 ;
	7'h3c :
		TR_202 = TR_75 ;
	7'h3d :
		TR_202 = TR_75 ;
	7'h3e :
		TR_202 = TR_75 ;
	7'h3f :
		TR_202 = 9'h000 ;	// line#=../rle.cpp:80
	7'h40 :
		TR_202 = TR_75 ;
	7'h41 :
		TR_202 = TR_75 ;
	7'h42 :
		TR_202 = TR_75 ;
	7'h43 :
		TR_202 = TR_75 ;
	7'h44 :
		TR_202 = TR_75 ;
	7'h45 :
		TR_202 = TR_75 ;
	7'h46 :
		TR_202 = TR_75 ;
	7'h47 :
		TR_202 = TR_75 ;
	7'h48 :
		TR_202 = TR_75 ;
	7'h49 :
		TR_202 = TR_75 ;
	7'h4a :
		TR_202 = TR_75 ;
	7'h4b :
		TR_202 = TR_75 ;
	7'h4c :
		TR_202 = TR_75 ;
	7'h4d :
		TR_202 = TR_75 ;
	7'h4e :
		TR_202 = TR_75 ;
	7'h4f :
		TR_202 = TR_75 ;
	7'h50 :
		TR_202 = TR_75 ;
	7'h51 :
		TR_202 = TR_75 ;
	7'h52 :
		TR_202 = TR_75 ;
	7'h53 :
		TR_202 = TR_75 ;
	7'h54 :
		TR_202 = TR_75 ;
	7'h55 :
		TR_202 = TR_75 ;
	7'h56 :
		TR_202 = TR_75 ;
	7'h57 :
		TR_202 = TR_75 ;
	7'h58 :
		TR_202 = TR_75 ;
	7'h59 :
		TR_202 = TR_75 ;
	7'h5a :
		TR_202 = TR_75 ;
	7'h5b :
		TR_202 = TR_75 ;
	7'h5c :
		TR_202 = TR_75 ;
	7'h5d :
		TR_202 = TR_75 ;
	7'h5e :
		TR_202 = TR_75 ;
	7'h5f :
		TR_202 = TR_75 ;
	7'h60 :
		TR_202 = TR_75 ;
	7'h61 :
		TR_202 = TR_75 ;
	7'h62 :
		TR_202 = TR_75 ;
	7'h63 :
		TR_202 = TR_75 ;
	7'h64 :
		TR_202 = TR_75 ;
	7'h65 :
		TR_202 = TR_75 ;
	7'h66 :
		TR_202 = TR_75 ;
	7'h67 :
		TR_202 = TR_75 ;
	7'h68 :
		TR_202 = TR_75 ;
	7'h69 :
		TR_202 = TR_75 ;
	7'h6a :
		TR_202 = TR_75 ;
	7'h6b :
		TR_202 = TR_75 ;
	7'h6c :
		TR_202 = TR_75 ;
	7'h6d :
		TR_202 = TR_75 ;
	7'h6e :
		TR_202 = TR_75 ;
	7'h6f :
		TR_202 = TR_75 ;
	7'h70 :
		TR_202 = TR_75 ;
	7'h71 :
		TR_202 = TR_75 ;
	7'h72 :
		TR_202 = TR_75 ;
	7'h73 :
		TR_202 = TR_75 ;
	7'h74 :
		TR_202 = TR_75 ;
	7'h75 :
		TR_202 = TR_75 ;
	7'h76 :
		TR_202 = TR_75 ;
	7'h77 :
		TR_202 = TR_75 ;
	7'h78 :
		TR_202 = TR_75 ;
	7'h79 :
		TR_202 = TR_75 ;
	7'h7a :
		TR_202 = TR_75 ;
	7'h7b :
		TR_202 = TR_75 ;
	7'h7c :
		TR_202 = TR_75 ;
	7'h7d :
		TR_202 = TR_75 ;
	7'h7e :
		TR_202 = TR_75 ;
	7'h7f :
		TR_202 = TR_75 ;
	default :
		TR_202 = 9'hx ;
	endcase
always @ ( TR_202 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_29 or 
	U_174 or RG_rl_160 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_63_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h3f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_63_t = ( ( { 9{ ST1_03d } } & RG_rl_160 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_29 )
		| ( { 9{ U_173 } } & TR_202 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_63_en = ( ST1_03d | U_174 | RG_rl_63_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_63_en )
		RG_rl_63 <= RG_rl_63_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_76 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_201 = TR_76 ;
	7'h01 :
		TR_201 = TR_76 ;
	7'h02 :
		TR_201 = TR_76 ;
	7'h03 :
		TR_201 = TR_76 ;
	7'h04 :
		TR_201 = TR_76 ;
	7'h05 :
		TR_201 = TR_76 ;
	7'h06 :
		TR_201 = TR_76 ;
	7'h07 :
		TR_201 = TR_76 ;
	7'h08 :
		TR_201 = TR_76 ;
	7'h09 :
		TR_201 = TR_76 ;
	7'h0a :
		TR_201 = TR_76 ;
	7'h0b :
		TR_201 = TR_76 ;
	7'h0c :
		TR_201 = TR_76 ;
	7'h0d :
		TR_201 = TR_76 ;
	7'h0e :
		TR_201 = TR_76 ;
	7'h0f :
		TR_201 = TR_76 ;
	7'h10 :
		TR_201 = TR_76 ;
	7'h11 :
		TR_201 = TR_76 ;
	7'h12 :
		TR_201 = TR_76 ;
	7'h13 :
		TR_201 = TR_76 ;
	7'h14 :
		TR_201 = TR_76 ;
	7'h15 :
		TR_201 = TR_76 ;
	7'h16 :
		TR_201 = TR_76 ;
	7'h17 :
		TR_201 = TR_76 ;
	7'h18 :
		TR_201 = TR_76 ;
	7'h19 :
		TR_201 = TR_76 ;
	7'h1a :
		TR_201 = TR_76 ;
	7'h1b :
		TR_201 = TR_76 ;
	7'h1c :
		TR_201 = TR_76 ;
	7'h1d :
		TR_201 = TR_76 ;
	7'h1e :
		TR_201 = TR_76 ;
	7'h1f :
		TR_201 = TR_76 ;
	7'h20 :
		TR_201 = TR_76 ;
	7'h21 :
		TR_201 = TR_76 ;
	7'h22 :
		TR_201 = TR_76 ;
	7'h23 :
		TR_201 = TR_76 ;
	7'h24 :
		TR_201 = TR_76 ;
	7'h25 :
		TR_201 = TR_76 ;
	7'h26 :
		TR_201 = TR_76 ;
	7'h27 :
		TR_201 = TR_76 ;
	7'h28 :
		TR_201 = TR_76 ;
	7'h29 :
		TR_201 = TR_76 ;
	7'h2a :
		TR_201 = TR_76 ;
	7'h2b :
		TR_201 = TR_76 ;
	7'h2c :
		TR_201 = TR_76 ;
	7'h2d :
		TR_201 = TR_76 ;
	7'h2e :
		TR_201 = TR_76 ;
	7'h2f :
		TR_201 = TR_76 ;
	7'h30 :
		TR_201 = TR_76 ;
	7'h31 :
		TR_201 = TR_76 ;
	7'h32 :
		TR_201 = TR_76 ;
	7'h33 :
		TR_201 = TR_76 ;
	7'h34 :
		TR_201 = TR_76 ;
	7'h35 :
		TR_201 = TR_76 ;
	7'h36 :
		TR_201 = TR_76 ;
	7'h37 :
		TR_201 = TR_76 ;
	7'h38 :
		TR_201 = TR_76 ;
	7'h39 :
		TR_201 = TR_76 ;
	7'h3a :
		TR_201 = TR_76 ;
	7'h3b :
		TR_201 = TR_76 ;
	7'h3c :
		TR_201 = TR_76 ;
	7'h3d :
		TR_201 = TR_76 ;
	7'h3e :
		TR_201 = TR_76 ;
	7'h3f :
		TR_201 = TR_76 ;
	7'h40 :
		TR_201 = 9'h000 ;	// line#=../rle.cpp:80
	7'h41 :
		TR_201 = TR_76 ;
	7'h42 :
		TR_201 = TR_76 ;
	7'h43 :
		TR_201 = TR_76 ;
	7'h44 :
		TR_201 = TR_76 ;
	7'h45 :
		TR_201 = TR_76 ;
	7'h46 :
		TR_201 = TR_76 ;
	7'h47 :
		TR_201 = TR_76 ;
	7'h48 :
		TR_201 = TR_76 ;
	7'h49 :
		TR_201 = TR_76 ;
	7'h4a :
		TR_201 = TR_76 ;
	7'h4b :
		TR_201 = TR_76 ;
	7'h4c :
		TR_201 = TR_76 ;
	7'h4d :
		TR_201 = TR_76 ;
	7'h4e :
		TR_201 = TR_76 ;
	7'h4f :
		TR_201 = TR_76 ;
	7'h50 :
		TR_201 = TR_76 ;
	7'h51 :
		TR_201 = TR_76 ;
	7'h52 :
		TR_201 = TR_76 ;
	7'h53 :
		TR_201 = TR_76 ;
	7'h54 :
		TR_201 = TR_76 ;
	7'h55 :
		TR_201 = TR_76 ;
	7'h56 :
		TR_201 = TR_76 ;
	7'h57 :
		TR_201 = TR_76 ;
	7'h58 :
		TR_201 = TR_76 ;
	7'h59 :
		TR_201 = TR_76 ;
	7'h5a :
		TR_201 = TR_76 ;
	7'h5b :
		TR_201 = TR_76 ;
	7'h5c :
		TR_201 = TR_76 ;
	7'h5d :
		TR_201 = TR_76 ;
	7'h5e :
		TR_201 = TR_76 ;
	7'h5f :
		TR_201 = TR_76 ;
	7'h60 :
		TR_201 = TR_76 ;
	7'h61 :
		TR_201 = TR_76 ;
	7'h62 :
		TR_201 = TR_76 ;
	7'h63 :
		TR_201 = TR_76 ;
	7'h64 :
		TR_201 = TR_76 ;
	7'h65 :
		TR_201 = TR_76 ;
	7'h66 :
		TR_201 = TR_76 ;
	7'h67 :
		TR_201 = TR_76 ;
	7'h68 :
		TR_201 = TR_76 ;
	7'h69 :
		TR_201 = TR_76 ;
	7'h6a :
		TR_201 = TR_76 ;
	7'h6b :
		TR_201 = TR_76 ;
	7'h6c :
		TR_201 = TR_76 ;
	7'h6d :
		TR_201 = TR_76 ;
	7'h6e :
		TR_201 = TR_76 ;
	7'h6f :
		TR_201 = TR_76 ;
	7'h70 :
		TR_201 = TR_76 ;
	7'h71 :
		TR_201 = TR_76 ;
	7'h72 :
		TR_201 = TR_76 ;
	7'h73 :
		TR_201 = TR_76 ;
	7'h74 :
		TR_201 = TR_76 ;
	7'h75 :
		TR_201 = TR_76 ;
	7'h76 :
		TR_201 = TR_76 ;
	7'h77 :
		TR_201 = TR_76 ;
	7'h78 :
		TR_201 = TR_76 ;
	7'h79 :
		TR_201 = TR_76 ;
	7'h7a :
		TR_201 = TR_76 ;
	7'h7b :
		TR_201 = TR_76 ;
	7'h7c :
		TR_201 = TR_76 ;
	7'h7d :
		TR_201 = TR_76 ;
	7'h7e :
		TR_201 = TR_76 ;
	7'h7f :
		TR_201 = TR_76 ;
	default :
		TR_201 = 9'hx ;
	endcase
always @ ( TR_201 or U_173 or sub8u_71ot or U_183 or RG_rl_161 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_64_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h40 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_64_t = ( ( { 9{ M_180 } } & RG_rl_161 )
		| ( { 9{ U_173 } } & TR_201 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_64_en = ( M_180 | RG_rl_64_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_64_en )
		RG_rl_64 <= RG_rl_64_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_77 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_200 = TR_77 ;
	7'h01 :
		TR_200 = TR_77 ;
	7'h02 :
		TR_200 = TR_77 ;
	7'h03 :
		TR_200 = TR_77 ;
	7'h04 :
		TR_200 = TR_77 ;
	7'h05 :
		TR_200 = TR_77 ;
	7'h06 :
		TR_200 = TR_77 ;
	7'h07 :
		TR_200 = TR_77 ;
	7'h08 :
		TR_200 = TR_77 ;
	7'h09 :
		TR_200 = TR_77 ;
	7'h0a :
		TR_200 = TR_77 ;
	7'h0b :
		TR_200 = TR_77 ;
	7'h0c :
		TR_200 = TR_77 ;
	7'h0d :
		TR_200 = TR_77 ;
	7'h0e :
		TR_200 = TR_77 ;
	7'h0f :
		TR_200 = TR_77 ;
	7'h10 :
		TR_200 = TR_77 ;
	7'h11 :
		TR_200 = TR_77 ;
	7'h12 :
		TR_200 = TR_77 ;
	7'h13 :
		TR_200 = TR_77 ;
	7'h14 :
		TR_200 = TR_77 ;
	7'h15 :
		TR_200 = TR_77 ;
	7'h16 :
		TR_200 = TR_77 ;
	7'h17 :
		TR_200 = TR_77 ;
	7'h18 :
		TR_200 = TR_77 ;
	7'h19 :
		TR_200 = TR_77 ;
	7'h1a :
		TR_200 = TR_77 ;
	7'h1b :
		TR_200 = TR_77 ;
	7'h1c :
		TR_200 = TR_77 ;
	7'h1d :
		TR_200 = TR_77 ;
	7'h1e :
		TR_200 = TR_77 ;
	7'h1f :
		TR_200 = TR_77 ;
	7'h20 :
		TR_200 = TR_77 ;
	7'h21 :
		TR_200 = TR_77 ;
	7'h22 :
		TR_200 = TR_77 ;
	7'h23 :
		TR_200 = TR_77 ;
	7'h24 :
		TR_200 = TR_77 ;
	7'h25 :
		TR_200 = TR_77 ;
	7'h26 :
		TR_200 = TR_77 ;
	7'h27 :
		TR_200 = TR_77 ;
	7'h28 :
		TR_200 = TR_77 ;
	7'h29 :
		TR_200 = TR_77 ;
	7'h2a :
		TR_200 = TR_77 ;
	7'h2b :
		TR_200 = TR_77 ;
	7'h2c :
		TR_200 = TR_77 ;
	7'h2d :
		TR_200 = TR_77 ;
	7'h2e :
		TR_200 = TR_77 ;
	7'h2f :
		TR_200 = TR_77 ;
	7'h30 :
		TR_200 = TR_77 ;
	7'h31 :
		TR_200 = TR_77 ;
	7'h32 :
		TR_200 = TR_77 ;
	7'h33 :
		TR_200 = TR_77 ;
	7'h34 :
		TR_200 = TR_77 ;
	7'h35 :
		TR_200 = TR_77 ;
	7'h36 :
		TR_200 = TR_77 ;
	7'h37 :
		TR_200 = TR_77 ;
	7'h38 :
		TR_200 = TR_77 ;
	7'h39 :
		TR_200 = TR_77 ;
	7'h3a :
		TR_200 = TR_77 ;
	7'h3b :
		TR_200 = TR_77 ;
	7'h3c :
		TR_200 = TR_77 ;
	7'h3d :
		TR_200 = TR_77 ;
	7'h3e :
		TR_200 = TR_77 ;
	7'h3f :
		TR_200 = TR_77 ;
	7'h40 :
		TR_200 = TR_77 ;
	7'h41 :
		TR_200 = 9'h000 ;	// line#=../rle.cpp:80
	7'h42 :
		TR_200 = TR_77 ;
	7'h43 :
		TR_200 = TR_77 ;
	7'h44 :
		TR_200 = TR_77 ;
	7'h45 :
		TR_200 = TR_77 ;
	7'h46 :
		TR_200 = TR_77 ;
	7'h47 :
		TR_200 = TR_77 ;
	7'h48 :
		TR_200 = TR_77 ;
	7'h49 :
		TR_200 = TR_77 ;
	7'h4a :
		TR_200 = TR_77 ;
	7'h4b :
		TR_200 = TR_77 ;
	7'h4c :
		TR_200 = TR_77 ;
	7'h4d :
		TR_200 = TR_77 ;
	7'h4e :
		TR_200 = TR_77 ;
	7'h4f :
		TR_200 = TR_77 ;
	7'h50 :
		TR_200 = TR_77 ;
	7'h51 :
		TR_200 = TR_77 ;
	7'h52 :
		TR_200 = TR_77 ;
	7'h53 :
		TR_200 = TR_77 ;
	7'h54 :
		TR_200 = TR_77 ;
	7'h55 :
		TR_200 = TR_77 ;
	7'h56 :
		TR_200 = TR_77 ;
	7'h57 :
		TR_200 = TR_77 ;
	7'h58 :
		TR_200 = TR_77 ;
	7'h59 :
		TR_200 = TR_77 ;
	7'h5a :
		TR_200 = TR_77 ;
	7'h5b :
		TR_200 = TR_77 ;
	7'h5c :
		TR_200 = TR_77 ;
	7'h5d :
		TR_200 = TR_77 ;
	7'h5e :
		TR_200 = TR_77 ;
	7'h5f :
		TR_200 = TR_77 ;
	7'h60 :
		TR_200 = TR_77 ;
	7'h61 :
		TR_200 = TR_77 ;
	7'h62 :
		TR_200 = TR_77 ;
	7'h63 :
		TR_200 = TR_77 ;
	7'h64 :
		TR_200 = TR_77 ;
	7'h65 :
		TR_200 = TR_77 ;
	7'h66 :
		TR_200 = TR_77 ;
	7'h67 :
		TR_200 = TR_77 ;
	7'h68 :
		TR_200 = TR_77 ;
	7'h69 :
		TR_200 = TR_77 ;
	7'h6a :
		TR_200 = TR_77 ;
	7'h6b :
		TR_200 = TR_77 ;
	7'h6c :
		TR_200 = TR_77 ;
	7'h6d :
		TR_200 = TR_77 ;
	7'h6e :
		TR_200 = TR_77 ;
	7'h6f :
		TR_200 = TR_77 ;
	7'h70 :
		TR_200 = TR_77 ;
	7'h71 :
		TR_200 = TR_77 ;
	7'h72 :
		TR_200 = TR_77 ;
	7'h73 :
		TR_200 = TR_77 ;
	7'h74 :
		TR_200 = TR_77 ;
	7'h75 :
		TR_200 = TR_77 ;
	7'h76 :
		TR_200 = TR_77 ;
	7'h77 :
		TR_200 = TR_77 ;
	7'h78 :
		TR_200 = TR_77 ;
	7'h79 :
		TR_200 = TR_77 ;
	7'h7a :
		TR_200 = TR_77 ;
	7'h7b :
		TR_200 = TR_77 ;
	7'h7c :
		TR_200 = TR_77 ;
	7'h7d :
		TR_200 = TR_77 ;
	7'h7e :
		TR_200 = TR_77 ;
	7'h7f :
		TR_200 = TR_77 ;
	default :
		TR_200 = 9'hx ;
	endcase
always @ ( TR_200 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_30 or 
	U_174 or RG_rl_161 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_65_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h41 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_65_t = ( ( { 9{ ST1_03d } } & RG_rl_161 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_30 )
		| ( { 9{ U_173 } } & TR_200 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_65_en = ( ST1_03d | U_174 | RG_rl_65_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_65_en )
		RG_rl_65 <= RG_rl_65_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_78 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_199 = TR_78 ;
	7'h01 :
		TR_199 = TR_78 ;
	7'h02 :
		TR_199 = TR_78 ;
	7'h03 :
		TR_199 = TR_78 ;
	7'h04 :
		TR_199 = TR_78 ;
	7'h05 :
		TR_199 = TR_78 ;
	7'h06 :
		TR_199 = TR_78 ;
	7'h07 :
		TR_199 = TR_78 ;
	7'h08 :
		TR_199 = TR_78 ;
	7'h09 :
		TR_199 = TR_78 ;
	7'h0a :
		TR_199 = TR_78 ;
	7'h0b :
		TR_199 = TR_78 ;
	7'h0c :
		TR_199 = TR_78 ;
	7'h0d :
		TR_199 = TR_78 ;
	7'h0e :
		TR_199 = TR_78 ;
	7'h0f :
		TR_199 = TR_78 ;
	7'h10 :
		TR_199 = TR_78 ;
	7'h11 :
		TR_199 = TR_78 ;
	7'h12 :
		TR_199 = TR_78 ;
	7'h13 :
		TR_199 = TR_78 ;
	7'h14 :
		TR_199 = TR_78 ;
	7'h15 :
		TR_199 = TR_78 ;
	7'h16 :
		TR_199 = TR_78 ;
	7'h17 :
		TR_199 = TR_78 ;
	7'h18 :
		TR_199 = TR_78 ;
	7'h19 :
		TR_199 = TR_78 ;
	7'h1a :
		TR_199 = TR_78 ;
	7'h1b :
		TR_199 = TR_78 ;
	7'h1c :
		TR_199 = TR_78 ;
	7'h1d :
		TR_199 = TR_78 ;
	7'h1e :
		TR_199 = TR_78 ;
	7'h1f :
		TR_199 = TR_78 ;
	7'h20 :
		TR_199 = TR_78 ;
	7'h21 :
		TR_199 = TR_78 ;
	7'h22 :
		TR_199 = TR_78 ;
	7'h23 :
		TR_199 = TR_78 ;
	7'h24 :
		TR_199 = TR_78 ;
	7'h25 :
		TR_199 = TR_78 ;
	7'h26 :
		TR_199 = TR_78 ;
	7'h27 :
		TR_199 = TR_78 ;
	7'h28 :
		TR_199 = TR_78 ;
	7'h29 :
		TR_199 = TR_78 ;
	7'h2a :
		TR_199 = TR_78 ;
	7'h2b :
		TR_199 = TR_78 ;
	7'h2c :
		TR_199 = TR_78 ;
	7'h2d :
		TR_199 = TR_78 ;
	7'h2e :
		TR_199 = TR_78 ;
	7'h2f :
		TR_199 = TR_78 ;
	7'h30 :
		TR_199 = TR_78 ;
	7'h31 :
		TR_199 = TR_78 ;
	7'h32 :
		TR_199 = TR_78 ;
	7'h33 :
		TR_199 = TR_78 ;
	7'h34 :
		TR_199 = TR_78 ;
	7'h35 :
		TR_199 = TR_78 ;
	7'h36 :
		TR_199 = TR_78 ;
	7'h37 :
		TR_199 = TR_78 ;
	7'h38 :
		TR_199 = TR_78 ;
	7'h39 :
		TR_199 = TR_78 ;
	7'h3a :
		TR_199 = TR_78 ;
	7'h3b :
		TR_199 = TR_78 ;
	7'h3c :
		TR_199 = TR_78 ;
	7'h3d :
		TR_199 = TR_78 ;
	7'h3e :
		TR_199 = TR_78 ;
	7'h3f :
		TR_199 = TR_78 ;
	7'h40 :
		TR_199 = TR_78 ;
	7'h41 :
		TR_199 = TR_78 ;
	7'h42 :
		TR_199 = 9'h000 ;	// line#=../rle.cpp:80
	7'h43 :
		TR_199 = TR_78 ;
	7'h44 :
		TR_199 = TR_78 ;
	7'h45 :
		TR_199 = TR_78 ;
	7'h46 :
		TR_199 = TR_78 ;
	7'h47 :
		TR_199 = TR_78 ;
	7'h48 :
		TR_199 = TR_78 ;
	7'h49 :
		TR_199 = TR_78 ;
	7'h4a :
		TR_199 = TR_78 ;
	7'h4b :
		TR_199 = TR_78 ;
	7'h4c :
		TR_199 = TR_78 ;
	7'h4d :
		TR_199 = TR_78 ;
	7'h4e :
		TR_199 = TR_78 ;
	7'h4f :
		TR_199 = TR_78 ;
	7'h50 :
		TR_199 = TR_78 ;
	7'h51 :
		TR_199 = TR_78 ;
	7'h52 :
		TR_199 = TR_78 ;
	7'h53 :
		TR_199 = TR_78 ;
	7'h54 :
		TR_199 = TR_78 ;
	7'h55 :
		TR_199 = TR_78 ;
	7'h56 :
		TR_199 = TR_78 ;
	7'h57 :
		TR_199 = TR_78 ;
	7'h58 :
		TR_199 = TR_78 ;
	7'h59 :
		TR_199 = TR_78 ;
	7'h5a :
		TR_199 = TR_78 ;
	7'h5b :
		TR_199 = TR_78 ;
	7'h5c :
		TR_199 = TR_78 ;
	7'h5d :
		TR_199 = TR_78 ;
	7'h5e :
		TR_199 = TR_78 ;
	7'h5f :
		TR_199 = TR_78 ;
	7'h60 :
		TR_199 = TR_78 ;
	7'h61 :
		TR_199 = TR_78 ;
	7'h62 :
		TR_199 = TR_78 ;
	7'h63 :
		TR_199 = TR_78 ;
	7'h64 :
		TR_199 = TR_78 ;
	7'h65 :
		TR_199 = TR_78 ;
	7'h66 :
		TR_199 = TR_78 ;
	7'h67 :
		TR_199 = TR_78 ;
	7'h68 :
		TR_199 = TR_78 ;
	7'h69 :
		TR_199 = TR_78 ;
	7'h6a :
		TR_199 = TR_78 ;
	7'h6b :
		TR_199 = TR_78 ;
	7'h6c :
		TR_199 = TR_78 ;
	7'h6d :
		TR_199 = TR_78 ;
	7'h6e :
		TR_199 = TR_78 ;
	7'h6f :
		TR_199 = TR_78 ;
	7'h70 :
		TR_199 = TR_78 ;
	7'h71 :
		TR_199 = TR_78 ;
	7'h72 :
		TR_199 = TR_78 ;
	7'h73 :
		TR_199 = TR_78 ;
	7'h74 :
		TR_199 = TR_78 ;
	7'h75 :
		TR_199 = TR_78 ;
	7'h76 :
		TR_199 = TR_78 ;
	7'h77 :
		TR_199 = TR_78 ;
	7'h78 :
		TR_199 = TR_78 ;
	7'h79 :
		TR_199 = TR_78 ;
	7'h7a :
		TR_199 = TR_78 ;
	7'h7b :
		TR_199 = TR_78 ;
	7'h7c :
		TR_199 = TR_78 ;
	7'h7d :
		TR_199 = TR_78 ;
	7'h7e :
		TR_199 = TR_78 ;
	7'h7f :
		TR_199 = TR_78 ;
	default :
		TR_199 = 9'hx ;
	endcase
always @ ( TR_199 or U_173 or sub8u_71ot or U_183 or RG_rl_162 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_66_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h42 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_66_t = ( ( { 9{ M_180 } } & RG_rl_162 )
		| ( { 9{ U_173 } } & TR_199 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_66_en = ( M_180 | RG_rl_66_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_66_en )
		RG_rl_66 <= RG_rl_66_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_79 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_198 = TR_79 ;
	7'h01 :
		TR_198 = TR_79 ;
	7'h02 :
		TR_198 = TR_79 ;
	7'h03 :
		TR_198 = TR_79 ;
	7'h04 :
		TR_198 = TR_79 ;
	7'h05 :
		TR_198 = TR_79 ;
	7'h06 :
		TR_198 = TR_79 ;
	7'h07 :
		TR_198 = TR_79 ;
	7'h08 :
		TR_198 = TR_79 ;
	7'h09 :
		TR_198 = TR_79 ;
	7'h0a :
		TR_198 = TR_79 ;
	7'h0b :
		TR_198 = TR_79 ;
	7'h0c :
		TR_198 = TR_79 ;
	7'h0d :
		TR_198 = TR_79 ;
	7'h0e :
		TR_198 = TR_79 ;
	7'h0f :
		TR_198 = TR_79 ;
	7'h10 :
		TR_198 = TR_79 ;
	7'h11 :
		TR_198 = TR_79 ;
	7'h12 :
		TR_198 = TR_79 ;
	7'h13 :
		TR_198 = TR_79 ;
	7'h14 :
		TR_198 = TR_79 ;
	7'h15 :
		TR_198 = TR_79 ;
	7'h16 :
		TR_198 = TR_79 ;
	7'h17 :
		TR_198 = TR_79 ;
	7'h18 :
		TR_198 = TR_79 ;
	7'h19 :
		TR_198 = TR_79 ;
	7'h1a :
		TR_198 = TR_79 ;
	7'h1b :
		TR_198 = TR_79 ;
	7'h1c :
		TR_198 = TR_79 ;
	7'h1d :
		TR_198 = TR_79 ;
	7'h1e :
		TR_198 = TR_79 ;
	7'h1f :
		TR_198 = TR_79 ;
	7'h20 :
		TR_198 = TR_79 ;
	7'h21 :
		TR_198 = TR_79 ;
	7'h22 :
		TR_198 = TR_79 ;
	7'h23 :
		TR_198 = TR_79 ;
	7'h24 :
		TR_198 = TR_79 ;
	7'h25 :
		TR_198 = TR_79 ;
	7'h26 :
		TR_198 = TR_79 ;
	7'h27 :
		TR_198 = TR_79 ;
	7'h28 :
		TR_198 = TR_79 ;
	7'h29 :
		TR_198 = TR_79 ;
	7'h2a :
		TR_198 = TR_79 ;
	7'h2b :
		TR_198 = TR_79 ;
	7'h2c :
		TR_198 = TR_79 ;
	7'h2d :
		TR_198 = TR_79 ;
	7'h2e :
		TR_198 = TR_79 ;
	7'h2f :
		TR_198 = TR_79 ;
	7'h30 :
		TR_198 = TR_79 ;
	7'h31 :
		TR_198 = TR_79 ;
	7'h32 :
		TR_198 = TR_79 ;
	7'h33 :
		TR_198 = TR_79 ;
	7'h34 :
		TR_198 = TR_79 ;
	7'h35 :
		TR_198 = TR_79 ;
	7'h36 :
		TR_198 = TR_79 ;
	7'h37 :
		TR_198 = TR_79 ;
	7'h38 :
		TR_198 = TR_79 ;
	7'h39 :
		TR_198 = TR_79 ;
	7'h3a :
		TR_198 = TR_79 ;
	7'h3b :
		TR_198 = TR_79 ;
	7'h3c :
		TR_198 = TR_79 ;
	7'h3d :
		TR_198 = TR_79 ;
	7'h3e :
		TR_198 = TR_79 ;
	7'h3f :
		TR_198 = TR_79 ;
	7'h40 :
		TR_198 = TR_79 ;
	7'h41 :
		TR_198 = TR_79 ;
	7'h42 :
		TR_198 = TR_79 ;
	7'h43 :
		TR_198 = 9'h000 ;	// line#=../rle.cpp:80
	7'h44 :
		TR_198 = TR_79 ;
	7'h45 :
		TR_198 = TR_79 ;
	7'h46 :
		TR_198 = TR_79 ;
	7'h47 :
		TR_198 = TR_79 ;
	7'h48 :
		TR_198 = TR_79 ;
	7'h49 :
		TR_198 = TR_79 ;
	7'h4a :
		TR_198 = TR_79 ;
	7'h4b :
		TR_198 = TR_79 ;
	7'h4c :
		TR_198 = TR_79 ;
	7'h4d :
		TR_198 = TR_79 ;
	7'h4e :
		TR_198 = TR_79 ;
	7'h4f :
		TR_198 = TR_79 ;
	7'h50 :
		TR_198 = TR_79 ;
	7'h51 :
		TR_198 = TR_79 ;
	7'h52 :
		TR_198 = TR_79 ;
	7'h53 :
		TR_198 = TR_79 ;
	7'h54 :
		TR_198 = TR_79 ;
	7'h55 :
		TR_198 = TR_79 ;
	7'h56 :
		TR_198 = TR_79 ;
	7'h57 :
		TR_198 = TR_79 ;
	7'h58 :
		TR_198 = TR_79 ;
	7'h59 :
		TR_198 = TR_79 ;
	7'h5a :
		TR_198 = TR_79 ;
	7'h5b :
		TR_198 = TR_79 ;
	7'h5c :
		TR_198 = TR_79 ;
	7'h5d :
		TR_198 = TR_79 ;
	7'h5e :
		TR_198 = TR_79 ;
	7'h5f :
		TR_198 = TR_79 ;
	7'h60 :
		TR_198 = TR_79 ;
	7'h61 :
		TR_198 = TR_79 ;
	7'h62 :
		TR_198 = TR_79 ;
	7'h63 :
		TR_198 = TR_79 ;
	7'h64 :
		TR_198 = TR_79 ;
	7'h65 :
		TR_198 = TR_79 ;
	7'h66 :
		TR_198 = TR_79 ;
	7'h67 :
		TR_198 = TR_79 ;
	7'h68 :
		TR_198 = TR_79 ;
	7'h69 :
		TR_198 = TR_79 ;
	7'h6a :
		TR_198 = TR_79 ;
	7'h6b :
		TR_198 = TR_79 ;
	7'h6c :
		TR_198 = TR_79 ;
	7'h6d :
		TR_198 = TR_79 ;
	7'h6e :
		TR_198 = TR_79 ;
	7'h6f :
		TR_198 = TR_79 ;
	7'h70 :
		TR_198 = TR_79 ;
	7'h71 :
		TR_198 = TR_79 ;
	7'h72 :
		TR_198 = TR_79 ;
	7'h73 :
		TR_198 = TR_79 ;
	7'h74 :
		TR_198 = TR_79 ;
	7'h75 :
		TR_198 = TR_79 ;
	7'h76 :
		TR_198 = TR_79 ;
	7'h77 :
		TR_198 = TR_79 ;
	7'h78 :
		TR_198 = TR_79 ;
	7'h79 :
		TR_198 = TR_79 ;
	7'h7a :
		TR_198 = TR_79 ;
	7'h7b :
		TR_198 = TR_79 ;
	7'h7c :
		TR_198 = TR_79 ;
	7'h7d :
		TR_198 = TR_79 ;
	7'h7e :
		TR_198 = TR_79 ;
	7'h7f :
		TR_198 = TR_79 ;
	default :
		TR_198 = 9'hx ;
	endcase
always @ ( TR_198 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_31 or 
	U_174 or RG_rl_162 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_67_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h43 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_67_t = ( ( { 9{ ST1_03d } } & RG_rl_162 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_31 )
		| ( { 9{ U_173 } } & TR_198 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_67_en = ( ST1_03d | U_174 | RG_rl_67_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_67_en )
		RG_rl_67 <= RG_rl_67_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_80 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_197 = TR_80 ;
	7'h01 :
		TR_197 = TR_80 ;
	7'h02 :
		TR_197 = TR_80 ;
	7'h03 :
		TR_197 = TR_80 ;
	7'h04 :
		TR_197 = TR_80 ;
	7'h05 :
		TR_197 = TR_80 ;
	7'h06 :
		TR_197 = TR_80 ;
	7'h07 :
		TR_197 = TR_80 ;
	7'h08 :
		TR_197 = TR_80 ;
	7'h09 :
		TR_197 = TR_80 ;
	7'h0a :
		TR_197 = TR_80 ;
	7'h0b :
		TR_197 = TR_80 ;
	7'h0c :
		TR_197 = TR_80 ;
	7'h0d :
		TR_197 = TR_80 ;
	7'h0e :
		TR_197 = TR_80 ;
	7'h0f :
		TR_197 = TR_80 ;
	7'h10 :
		TR_197 = TR_80 ;
	7'h11 :
		TR_197 = TR_80 ;
	7'h12 :
		TR_197 = TR_80 ;
	7'h13 :
		TR_197 = TR_80 ;
	7'h14 :
		TR_197 = TR_80 ;
	7'h15 :
		TR_197 = TR_80 ;
	7'h16 :
		TR_197 = TR_80 ;
	7'h17 :
		TR_197 = TR_80 ;
	7'h18 :
		TR_197 = TR_80 ;
	7'h19 :
		TR_197 = TR_80 ;
	7'h1a :
		TR_197 = TR_80 ;
	7'h1b :
		TR_197 = TR_80 ;
	7'h1c :
		TR_197 = TR_80 ;
	7'h1d :
		TR_197 = TR_80 ;
	7'h1e :
		TR_197 = TR_80 ;
	7'h1f :
		TR_197 = TR_80 ;
	7'h20 :
		TR_197 = TR_80 ;
	7'h21 :
		TR_197 = TR_80 ;
	7'h22 :
		TR_197 = TR_80 ;
	7'h23 :
		TR_197 = TR_80 ;
	7'h24 :
		TR_197 = TR_80 ;
	7'h25 :
		TR_197 = TR_80 ;
	7'h26 :
		TR_197 = TR_80 ;
	7'h27 :
		TR_197 = TR_80 ;
	7'h28 :
		TR_197 = TR_80 ;
	7'h29 :
		TR_197 = TR_80 ;
	7'h2a :
		TR_197 = TR_80 ;
	7'h2b :
		TR_197 = TR_80 ;
	7'h2c :
		TR_197 = TR_80 ;
	7'h2d :
		TR_197 = TR_80 ;
	7'h2e :
		TR_197 = TR_80 ;
	7'h2f :
		TR_197 = TR_80 ;
	7'h30 :
		TR_197 = TR_80 ;
	7'h31 :
		TR_197 = TR_80 ;
	7'h32 :
		TR_197 = TR_80 ;
	7'h33 :
		TR_197 = TR_80 ;
	7'h34 :
		TR_197 = TR_80 ;
	7'h35 :
		TR_197 = TR_80 ;
	7'h36 :
		TR_197 = TR_80 ;
	7'h37 :
		TR_197 = TR_80 ;
	7'h38 :
		TR_197 = TR_80 ;
	7'h39 :
		TR_197 = TR_80 ;
	7'h3a :
		TR_197 = TR_80 ;
	7'h3b :
		TR_197 = TR_80 ;
	7'h3c :
		TR_197 = TR_80 ;
	7'h3d :
		TR_197 = TR_80 ;
	7'h3e :
		TR_197 = TR_80 ;
	7'h3f :
		TR_197 = TR_80 ;
	7'h40 :
		TR_197 = TR_80 ;
	7'h41 :
		TR_197 = TR_80 ;
	7'h42 :
		TR_197 = TR_80 ;
	7'h43 :
		TR_197 = TR_80 ;
	7'h44 :
		TR_197 = 9'h000 ;	// line#=../rle.cpp:80
	7'h45 :
		TR_197 = TR_80 ;
	7'h46 :
		TR_197 = TR_80 ;
	7'h47 :
		TR_197 = TR_80 ;
	7'h48 :
		TR_197 = TR_80 ;
	7'h49 :
		TR_197 = TR_80 ;
	7'h4a :
		TR_197 = TR_80 ;
	7'h4b :
		TR_197 = TR_80 ;
	7'h4c :
		TR_197 = TR_80 ;
	7'h4d :
		TR_197 = TR_80 ;
	7'h4e :
		TR_197 = TR_80 ;
	7'h4f :
		TR_197 = TR_80 ;
	7'h50 :
		TR_197 = TR_80 ;
	7'h51 :
		TR_197 = TR_80 ;
	7'h52 :
		TR_197 = TR_80 ;
	7'h53 :
		TR_197 = TR_80 ;
	7'h54 :
		TR_197 = TR_80 ;
	7'h55 :
		TR_197 = TR_80 ;
	7'h56 :
		TR_197 = TR_80 ;
	7'h57 :
		TR_197 = TR_80 ;
	7'h58 :
		TR_197 = TR_80 ;
	7'h59 :
		TR_197 = TR_80 ;
	7'h5a :
		TR_197 = TR_80 ;
	7'h5b :
		TR_197 = TR_80 ;
	7'h5c :
		TR_197 = TR_80 ;
	7'h5d :
		TR_197 = TR_80 ;
	7'h5e :
		TR_197 = TR_80 ;
	7'h5f :
		TR_197 = TR_80 ;
	7'h60 :
		TR_197 = TR_80 ;
	7'h61 :
		TR_197 = TR_80 ;
	7'h62 :
		TR_197 = TR_80 ;
	7'h63 :
		TR_197 = TR_80 ;
	7'h64 :
		TR_197 = TR_80 ;
	7'h65 :
		TR_197 = TR_80 ;
	7'h66 :
		TR_197 = TR_80 ;
	7'h67 :
		TR_197 = TR_80 ;
	7'h68 :
		TR_197 = TR_80 ;
	7'h69 :
		TR_197 = TR_80 ;
	7'h6a :
		TR_197 = TR_80 ;
	7'h6b :
		TR_197 = TR_80 ;
	7'h6c :
		TR_197 = TR_80 ;
	7'h6d :
		TR_197 = TR_80 ;
	7'h6e :
		TR_197 = TR_80 ;
	7'h6f :
		TR_197 = TR_80 ;
	7'h70 :
		TR_197 = TR_80 ;
	7'h71 :
		TR_197 = TR_80 ;
	7'h72 :
		TR_197 = TR_80 ;
	7'h73 :
		TR_197 = TR_80 ;
	7'h74 :
		TR_197 = TR_80 ;
	7'h75 :
		TR_197 = TR_80 ;
	7'h76 :
		TR_197 = TR_80 ;
	7'h77 :
		TR_197 = TR_80 ;
	7'h78 :
		TR_197 = TR_80 ;
	7'h79 :
		TR_197 = TR_80 ;
	7'h7a :
		TR_197 = TR_80 ;
	7'h7b :
		TR_197 = TR_80 ;
	7'h7c :
		TR_197 = TR_80 ;
	7'h7d :
		TR_197 = TR_80 ;
	7'h7e :
		TR_197 = TR_80 ;
	7'h7f :
		TR_197 = TR_80 ;
	default :
		TR_197 = 9'hx ;
	endcase
always @ ( TR_197 or U_173 or sub8u_71ot or U_183 or RG_rl_163 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_68_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h44 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_68_t = ( ( { 9{ M_180 } } & RG_rl_163 )
		| ( { 9{ U_173 } } & TR_197 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_68_en = ( M_180 | RG_rl_68_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_68_en )
		RG_rl_68 <= RG_rl_68_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_81 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_196 = TR_81 ;
	7'h01 :
		TR_196 = TR_81 ;
	7'h02 :
		TR_196 = TR_81 ;
	7'h03 :
		TR_196 = TR_81 ;
	7'h04 :
		TR_196 = TR_81 ;
	7'h05 :
		TR_196 = TR_81 ;
	7'h06 :
		TR_196 = TR_81 ;
	7'h07 :
		TR_196 = TR_81 ;
	7'h08 :
		TR_196 = TR_81 ;
	7'h09 :
		TR_196 = TR_81 ;
	7'h0a :
		TR_196 = TR_81 ;
	7'h0b :
		TR_196 = TR_81 ;
	7'h0c :
		TR_196 = TR_81 ;
	7'h0d :
		TR_196 = TR_81 ;
	7'h0e :
		TR_196 = TR_81 ;
	7'h0f :
		TR_196 = TR_81 ;
	7'h10 :
		TR_196 = TR_81 ;
	7'h11 :
		TR_196 = TR_81 ;
	7'h12 :
		TR_196 = TR_81 ;
	7'h13 :
		TR_196 = TR_81 ;
	7'h14 :
		TR_196 = TR_81 ;
	7'h15 :
		TR_196 = TR_81 ;
	7'h16 :
		TR_196 = TR_81 ;
	7'h17 :
		TR_196 = TR_81 ;
	7'h18 :
		TR_196 = TR_81 ;
	7'h19 :
		TR_196 = TR_81 ;
	7'h1a :
		TR_196 = TR_81 ;
	7'h1b :
		TR_196 = TR_81 ;
	7'h1c :
		TR_196 = TR_81 ;
	7'h1d :
		TR_196 = TR_81 ;
	7'h1e :
		TR_196 = TR_81 ;
	7'h1f :
		TR_196 = TR_81 ;
	7'h20 :
		TR_196 = TR_81 ;
	7'h21 :
		TR_196 = TR_81 ;
	7'h22 :
		TR_196 = TR_81 ;
	7'h23 :
		TR_196 = TR_81 ;
	7'h24 :
		TR_196 = TR_81 ;
	7'h25 :
		TR_196 = TR_81 ;
	7'h26 :
		TR_196 = TR_81 ;
	7'h27 :
		TR_196 = TR_81 ;
	7'h28 :
		TR_196 = TR_81 ;
	7'h29 :
		TR_196 = TR_81 ;
	7'h2a :
		TR_196 = TR_81 ;
	7'h2b :
		TR_196 = TR_81 ;
	7'h2c :
		TR_196 = TR_81 ;
	7'h2d :
		TR_196 = TR_81 ;
	7'h2e :
		TR_196 = TR_81 ;
	7'h2f :
		TR_196 = TR_81 ;
	7'h30 :
		TR_196 = TR_81 ;
	7'h31 :
		TR_196 = TR_81 ;
	7'h32 :
		TR_196 = TR_81 ;
	7'h33 :
		TR_196 = TR_81 ;
	7'h34 :
		TR_196 = TR_81 ;
	7'h35 :
		TR_196 = TR_81 ;
	7'h36 :
		TR_196 = TR_81 ;
	7'h37 :
		TR_196 = TR_81 ;
	7'h38 :
		TR_196 = TR_81 ;
	7'h39 :
		TR_196 = TR_81 ;
	7'h3a :
		TR_196 = TR_81 ;
	7'h3b :
		TR_196 = TR_81 ;
	7'h3c :
		TR_196 = TR_81 ;
	7'h3d :
		TR_196 = TR_81 ;
	7'h3e :
		TR_196 = TR_81 ;
	7'h3f :
		TR_196 = TR_81 ;
	7'h40 :
		TR_196 = TR_81 ;
	7'h41 :
		TR_196 = TR_81 ;
	7'h42 :
		TR_196 = TR_81 ;
	7'h43 :
		TR_196 = TR_81 ;
	7'h44 :
		TR_196 = TR_81 ;
	7'h45 :
		TR_196 = 9'h000 ;	// line#=../rle.cpp:80
	7'h46 :
		TR_196 = TR_81 ;
	7'h47 :
		TR_196 = TR_81 ;
	7'h48 :
		TR_196 = TR_81 ;
	7'h49 :
		TR_196 = TR_81 ;
	7'h4a :
		TR_196 = TR_81 ;
	7'h4b :
		TR_196 = TR_81 ;
	7'h4c :
		TR_196 = TR_81 ;
	7'h4d :
		TR_196 = TR_81 ;
	7'h4e :
		TR_196 = TR_81 ;
	7'h4f :
		TR_196 = TR_81 ;
	7'h50 :
		TR_196 = TR_81 ;
	7'h51 :
		TR_196 = TR_81 ;
	7'h52 :
		TR_196 = TR_81 ;
	7'h53 :
		TR_196 = TR_81 ;
	7'h54 :
		TR_196 = TR_81 ;
	7'h55 :
		TR_196 = TR_81 ;
	7'h56 :
		TR_196 = TR_81 ;
	7'h57 :
		TR_196 = TR_81 ;
	7'h58 :
		TR_196 = TR_81 ;
	7'h59 :
		TR_196 = TR_81 ;
	7'h5a :
		TR_196 = TR_81 ;
	7'h5b :
		TR_196 = TR_81 ;
	7'h5c :
		TR_196 = TR_81 ;
	7'h5d :
		TR_196 = TR_81 ;
	7'h5e :
		TR_196 = TR_81 ;
	7'h5f :
		TR_196 = TR_81 ;
	7'h60 :
		TR_196 = TR_81 ;
	7'h61 :
		TR_196 = TR_81 ;
	7'h62 :
		TR_196 = TR_81 ;
	7'h63 :
		TR_196 = TR_81 ;
	7'h64 :
		TR_196 = TR_81 ;
	7'h65 :
		TR_196 = TR_81 ;
	7'h66 :
		TR_196 = TR_81 ;
	7'h67 :
		TR_196 = TR_81 ;
	7'h68 :
		TR_196 = TR_81 ;
	7'h69 :
		TR_196 = TR_81 ;
	7'h6a :
		TR_196 = TR_81 ;
	7'h6b :
		TR_196 = TR_81 ;
	7'h6c :
		TR_196 = TR_81 ;
	7'h6d :
		TR_196 = TR_81 ;
	7'h6e :
		TR_196 = TR_81 ;
	7'h6f :
		TR_196 = TR_81 ;
	7'h70 :
		TR_196 = TR_81 ;
	7'h71 :
		TR_196 = TR_81 ;
	7'h72 :
		TR_196 = TR_81 ;
	7'h73 :
		TR_196 = TR_81 ;
	7'h74 :
		TR_196 = TR_81 ;
	7'h75 :
		TR_196 = TR_81 ;
	7'h76 :
		TR_196 = TR_81 ;
	7'h77 :
		TR_196 = TR_81 ;
	7'h78 :
		TR_196 = TR_81 ;
	7'h79 :
		TR_196 = TR_81 ;
	7'h7a :
		TR_196 = TR_81 ;
	7'h7b :
		TR_196 = TR_81 ;
	7'h7c :
		TR_196 = TR_81 ;
	7'h7d :
		TR_196 = TR_81 ;
	7'h7e :
		TR_196 = TR_81 ;
	7'h7f :
		TR_196 = TR_81 ;
	default :
		TR_196 = 9'hx ;
	endcase
always @ ( TR_196 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_32 or 
	U_174 or RG_rl_163 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_69_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h45 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_69_t = ( ( { 9{ ST1_03d } } & RG_rl_163 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_32 )
		| ( { 9{ U_173 } } & TR_196 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_69_en = ( ST1_03d | U_174 | RG_rl_69_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_69_en )
		RG_rl_69 <= RG_rl_69_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_82 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_195 = TR_82 ;
	7'h01 :
		TR_195 = TR_82 ;
	7'h02 :
		TR_195 = TR_82 ;
	7'h03 :
		TR_195 = TR_82 ;
	7'h04 :
		TR_195 = TR_82 ;
	7'h05 :
		TR_195 = TR_82 ;
	7'h06 :
		TR_195 = TR_82 ;
	7'h07 :
		TR_195 = TR_82 ;
	7'h08 :
		TR_195 = TR_82 ;
	7'h09 :
		TR_195 = TR_82 ;
	7'h0a :
		TR_195 = TR_82 ;
	7'h0b :
		TR_195 = TR_82 ;
	7'h0c :
		TR_195 = TR_82 ;
	7'h0d :
		TR_195 = TR_82 ;
	7'h0e :
		TR_195 = TR_82 ;
	7'h0f :
		TR_195 = TR_82 ;
	7'h10 :
		TR_195 = TR_82 ;
	7'h11 :
		TR_195 = TR_82 ;
	7'h12 :
		TR_195 = TR_82 ;
	7'h13 :
		TR_195 = TR_82 ;
	7'h14 :
		TR_195 = TR_82 ;
	7'h15 :
		TR_195 = TR_82 ;
	7'h16 :
		TR_195 = TR_82 ;
	7'h17 :
		TR_195 = TR_82 ;
	7'h18 :
		TR_195 = TR_82 ;
	7'h19 :
		TR_195 = TR_82 ;
	7'h1a :
		TR_195 = TR_82 ;
	7'h1b :
		TR_195 = TR_82 ;
	7'h1c :
		TR_195 = TR_82 ;
	7'h1d :
		TR_195 = TR_82 ;
	7'h1e :
		TR_195 = TR_82 ;
	7'h1f :
		TR_195 = TR_82 ;
	7'h20 :
		TR_195 = TR_82 ;
	7'h21 :
		TR_195 = TR_82 ;
	7'h22 :
		TR_195 = TR_82 ;
	7'h23 :
		TR_195 = TR_82 ;
	7'h24 :
		TR_195 = TR_82 ;
	7'h25 :
		TR_195 = TR_82 ;
	7'h26 :
		TR_195 = TR_82 ;
	7'h27 :
		TR_195 = TR_82 ;
	7'h28 :
		TR_195 = TR_82 ;
	7'h29 :
		TR_195 = TR_82 ;
	7'h2a :
		TR_195 = TR_82 ;
	7'h2b :
		TR_195 = TR_82 ;
	7'h2c :
		TR_195 = TR_82 ;
	7'h2d :
		TR_195 = TR_82 ;
	7'h2e :
		TR_195 = TR_82 ;
	7'h2f :
		TR_195 = TR_82 ;
	7'h30 :
		TR_195 = TR_82 ;
	7'h31 :
		TR_195 = TR_82 ;
	7'h32 :
		TR_195 = TR_82 ;
	7'h33 :
		TR_195 = TR_82 ;
	7'h34 :
		TR_195 = TR_82 ;
	7'h35 :
		TR_195 = TR_82 ;
	7'h36 :
		TR_195 = TR_82 ;
	7'h37 :
		TR_195 = TR_82 ;
	7'h38 :
		TR_195 = TR_82 ;
	7'h39 :
		TR_195 = TR_82 ;
	7'h3a :
		TR_195 = TR_82 ;
	7'h3b :
		TR_195 = TR_82 ;
	7'h3c :
		TR_195 = TR_82 ;
	7'h3d :
		TR_195 = TR_82 ;
	7'h3e :
		TR_195 = TR_82 ;
	7'h3f :
		TR_195 = TR_82 ;
	7'h40 :
		TR_195 = TR_82 ;
	7'h41 :
		TR_195 = TR_82 ;
	7'h42 :
		TR_195 = TR_82 ;
	7'h43 :
		TR_195 = TR_82 ;
	7'h44 :
		TR_195 = TR_82 ;
	7'h45 :
		TR_195 = TR_82 ;
	7'h46 :
		TR_195 = 9'h000 ;	// line#=../rle.cpp:80
	7'h47 :
		TR_195 = TR_82 ;
	7'h48 :
		TR_195 = TR_82 ;
	7'h49 :
		TR_195 = TR_82 ;
	7'h4a :
		TR_195 = TR_82 ;
	7'h4b :
		TR_195 = TR_82 ;
	7'h4c :
		TR_195 = TR_82 ;
	7'h4d :
		TR_195 = TR_82 ;
	7'h4e :
		TR_195 = TR_82 ;
	7'h4f :
		TR_195 = TR_82 ;
	7'h50 :
		TR_195 = TR_82 ;
	7'h51 :
		TR_195 = TR_82 ;
	7'h52 :
		TR_195 = TR_82 ;
	7'h53 :
		TR_195 = TR_82 ;
	7'h54 :
		TR_195 = TR_82 ;
	7'h55 :
		TR_195 = TR_82 ;
	7'h56 :
		TR_195 = TR_82 ;
	7'h57 :
		TR_195 = TR_82 ;
	7'h58 :
		TR_195 = TR_82 ;
	7'h59 :
		TR_195 = TR_82 ;
	7'h5a :
		TR_195 = TR_82 ;
	7'h5b :
		TR_195 = TR_82 ;
	7'h5c :
		TR_195 = TR_82 ;
	7'h5d :
		TR_195 = TR_82 ;
	7'h5e :
		TR_195 = TR_82 ;
	7'h5f :
		TR_195 = TR_82 ;
	7'h60 :
		TR_195 = TR_82 ;
	7'h61 :
		TR_195 = TR_82 ;
	7'h62 :
		TR_195 = TR_82 ;
	7'h63 :
		TR_195 = TR_82 ;
	7'h64 :
		TR_195 = TR_82 ;
	7'h65 :
		TR_195 = TR_82 ;
	7'h66 :
		TR_195 = TR_82 ;
	7'h67 :
		TR_195 = TR_82 ;
	7'h68 :
		TR_195 = TR_82 ;
	7'h69 :
		TR_195 = TR_82 ;
	7'h6a :
		TR_195 = TR_82 ;
	7'h6b :
		TR_195 = TR_82 ;
	7'h6c :
		TR_195 = TR_82 ;
	7'h6d :
		TR_195 = TR_82 ;
	7'h6e :
		TR_195 = TR_82 ;
	7'h6f :
		TR_195 = TR_82 ;
	7'h70 :
		TR_195 = TR_82 ;
	7'h71 :
		TR_195 = TR_82 ;
	7'h72 :
		TR_195 = TR_82 ;
	7'h73 :
		TR_195 = TR_82 ;
	7'h74 :
		TR_195 = TR_82 ;
	7'h75 :
		TR_195 = TR_82 ;
	7'h76 :
		TR_195 = TR_82 ;
	7'h77 :
		TR_195 = TR_82 ;
	7'h78 :
		TR_195 = TR_82 ;
	7'h79 :
		TR_195 = TR_82 ;
	7'h7a :
		TR_195 = TR_82 ;
	7'h7b :
		TR_195 = TR_82 ;
	7'h7c :
		TR_195 = TR_82 ;
	7'h7d :
		TR_195 = TR_82 ;
	7'h7e :
		TR_195 = TR_82 ;
	7'h7f :
		TR_195 = TR_82 ;
	default :
		TR_195 = 9'hx ;
	endcase
always @ ( TR_195 or U_173 or sub8u_71ot or U_183 or RG_rl_164 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_70_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h46 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_70_t = ( ( { 9{ M_180 } } & RG_rl_164 )
		| ( { 9{ U_173 } } & TR_195 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_70_en = ( M_180 | RG_rl_70_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_70_en )
		RG_rl_70 <= RG_rl_70_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_83 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_194 = TR_83 ;
	7'h01 :
		TR_194 = TR_83 ;
	7'h02 :
		TR_194 = TR_83 ;
	7'h03 :
		TR_194 = TR_83 ;
	7'h04 :
		TR_194 = TR_83 ;
	7'h05 :
		TR_194 = TR_83 ;
	7'h06 :
		TR_194 = TR_83 ;
	7'h07 :
		TR_194 = TR_83 ;
	7'h08 :
		TR_194 = TR_83 ;
	7'h09 :
		TR_194 = TR_83 ;
	7'h0a :
		TR_194 = TR_83 ;
	7'h0b :
		TR_194 = TR_83 ;
	7'h0c :
		TR_194 = TR_83 ;
	7'h0d :
		TR_194 = TR_83 ;
	7'h0e :
		TR_194 = TR_83 ;
	7'h0f :
		TR_194 = TR_83 ;
	7'h10 :
		TR_194 = TR_83 ;
	7'h11 :
		TR_194 = TR_83 ;
	7'h12 :
		TR_194 = TR_83 ;
	7'h13 :
		TR_194 = TR_83 ;
	7'h14 :
		TR_194 = TR_83 ;
	7'h15 :
		TR_194 = TR_83 ;
	7'h16 :
		TR_194 = TR_83 ;
	7'h17 :
		TR_194 = TR_83 ;
	7'h18 :
		TR_194 = TR_83 ;
	7'h19 :
		TR_194 = TR_83 ;
	7'h1a :
		TR_194 = TR_83 ;
	7'h1b :
		TR_194 = TR_83 ;
	7'h1c :
		TR_194 = TR_83 ;
	7'h1d :
		TR_194 = TR_83 ;
	7'h1e :
		TR_194 = TR_83 ;
	7'h1f :
		TR_194 = TR_83 ;
	7'h20 :
		TR_194 = TR_83 ;
	7'h21 :
		TR_194 = TR_83 ;
	7'h22 :
		TR_194 = TR_83 ;
	7'h23 :
		TR_194 = TR_83 ;
	7'h24 :
		TR_194 = TR_83 ;
	7'h25 :
		TR_194 = TR_83 ;
	7'h26 :
		TR_194 = TR_83 ;
	7'h27 :
		TR_194 = TR_83 ;
	7'h28 :
		TR_194 = TR_83 ;
	7'h29 :
		TR_194 = TR_83 ;
	7'h2a :
		TR_194 = TR_83 ;
	7'h2b :
		TR_194 = TR_83 ;
	7'h2c :
		TR_194 = TR_83 ;
	7'h2d :
		TR_194 = TR_83 ;
	7'h2e :
		TR_194 = TR_83 ;
	7'h2f :
		TR_194 = TR_83 ;
	7'h30 :
		TR_194 = TR_83 ;
	7'h31 :
		TR_194 = TR_83 ;
	7'h32 :
		TR_194 = TR_83 ;
	7'h33 :
		TR_194 = TR_83 ;
	7'h34 :
		TR_194 = TR_83 ;
	7'h35 :
		TR_194 = TR_83 ;
	7'h36 :
		TR_194 = TR_83 ;
	7'h37 :
		TR_194 = TR_83 ;
	7'h38 :
		TR_194 = TR_83 ;
	7'h39 :
		TR_194 = TR_83 ;
	7'h3a :
		TR_194 = TR_83 ;
	7'h3b :
		TR_194 = TR_83 ;
	7'h3c :
		TR_194 = TR_83 ;
	7'h3d :
		TR_194 = TR_83 ;
	7'h3e :
		TR_194 = TR_83 ;
	7'h3f :
		TR_194 = TR_83 ;
	7'h40 :
		TR_194 = TR_83 ;
	7'h41 :
		TR_194 = TR_83 ;
	7'h42 :
		TR_194 = TR_83 ;
	7'h43 :
		TR_194 = TR_83 ;
	7'h44 :
		TR_194 = TR_83 ;
	7'h45 :
		TR_194 = TR_83 ;
	7'h46 :
		TR_194 = TR_83 ;
	7'h47 :
		TR_194 = 9'h000 ;	// line#=../rle.cpp:80
	7'h48 :
		TR_194 = TR_83 ;
	7'h49 :
		TR_194 = TR_83 ;
	7'h4a :
		TR_194 = TR_83 ;
	7'h4b :
		TR_194 = TR_83 ;
	7'h4c :
		TR_194 = TR_83 ;
	7'h4d :
		TR_194 = TR_83 ;
	7'h4e :
		TR_194 = TR_83 ;
	7'h4f :
		TR_194 = TR_83 ;
	7'h50 :
		TR_194 = TR_83 ;
	7'h51 :
		TR_194 = TR_83 ;
	7'h52 :
		TR_194 = TR_83 ;
	7'h53 :
		TR_194 = TR_83 ;
	7'h54 :
		TR_194 = TR_83 ;
	7'h55 :
		TR_194 = TR_83 ;
	7'h56 :
		TR_194 = TR_83 ;
	7'h57 :
		TR_194 = TR_83 ;
	7'h58 :
		TR_194 = TR_83 ;
	7'h59 :
		TR_194 = TR_83 ;
	7'h5a :
		TR_194 = TR_83 ;
	7'h5b :
		TR_194 = TR_83 ;
	7'h5c :
		TR_194 = TR_83 ;
	7'h5d :
		TR_194 = TR_83 ;
	7'h5e :
		TR_194 = TR_83 ;
	7'h5f :
		TR_194 = TR_83 ;
	7'h60 :
		TR_194 = TR_83 ;
	7'h61 :
		TR_194 = TR_83 ;
	7'h62 :
		TR_194 = TR_83 ;
	7'h63 :
		TR_194 = TR_83 ;
	7'h64 :
		TR_194 = TR_83 ;
	7'h65 :
		TR_194 = TR_83 ;
	7'h66 :
		TR_194 = TR_83 ;
	7'h67 :
		TR_194 = TR_83 ;
	7'h68 :
		TR_194 = TR_83 ;
	7'h69 :
		TR_194 = TR_83 ;
	7'h6a :
		TR_194 = TR_83 ;
	7'h6b :
		TR_194 = TR_83 ;
	7'h6c :
		TR_194 = TR_83 ;
	7'h6d :
		TR_194 = TR_83 ;
	7'h6e :
		TR_194 = TR_83 ;
	7'h6f :
		TR_194 = TR_83 ;
	7'h70 :
		TR_194 = TR_83 ;
	7'h71 :
		TR_194 = TR_83 ;
	7'h72 :
		TR_194 = TR_83 ;
	7'h73 :
		TR_194 = TR_83 ;
	7'h74 :
		TR_194 = TR_83 ;
	7'h75 :
		TR_194 = TR_83 ;
	7'h76 :
		TR_194 = TR_83 ;
	7'h77 :
		TR_194 = TR_83 ;
	7'h78 :
		TR_194 = TR_83 ;
	7'h79 :
		TR_194 = TR_83 ;
	7'h7a :
		TR_194 = TR_83 ;
	7'h7b :
		TR_194 = TR_83 ;
	7'h7c :
		TR_194 = TR_83 ;
	7'h7d :
		TR_194 = TR_83 ;
	7'h7e :
		TR_194 = TR_83 ;
	7'h7f :
		TR_194 = TR_83 ;
	default :
		TR_194 = 9'hx ;
	endcase
always @ ( TR_194 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_33 or 
	U_174 or RG_rl_164 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_71_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h47 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_71_t = ( ( { 9{ ST1_03d } } & RG_rl_164 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_33 )
		| ( { 9{ U_173 } } & TR_194 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_71_en = ( ST1_03d | U_174 | RG_rl_71_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_71_en )
		RG_rl_71 <= RG_rl_71_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_84 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_193 = TR_84 ;
	7'h01 :
		TR_193 = TR_84 ;
	7'h02 :
		TR_193 = TR_84 ;
	7'h03 :
		TR_193 = TR_84 ;
	7'h04 :
		TR_193 = TR_84 ;
	7'h05 :
		TR_193 = TR_84 ;
	7'h06 :
		TR_193 = TR_84 ;
	7'h07 :
		TR_193 = TR_84 ;
	7'h08 :
		TR_193 = TR_84 ;
	7'h09 :
		TR_193 = TR_84 ;
	7'h0a :
		TR_193 = TR_84 ;
	7'h0b :
		TR_193 = TR_84 ;
	7'h0c :
		TR_193 = TR_84 ;
	7'h0d :
		TR_193 = TR_84 ;
	7'h0e :
		TR_193 = TR_84 ;
	7'h0f :
		TR_193 = TR_84 ;
	7'h10 :
		TR_193 = TR_84 ;
	7'h11 :
		TR_193 = TR_84 ;
	7'h12 :
		TR_193 = TR_84 ;
	7'h13 :
		TR_193 = TR_84 ;
	7'h14 :
		TR_193 = TR_84 ;
	7'h15 :
		TR_193 = TR_84 ;
	7'h16 :
		TR_193 = TR_84 ;
	7'h17 :
		TR_193 = TR_84 ;
	7'h18 :
		TR_193 = TR_84 ;
	7'h19 :
		TR_193 = TR_84 ;
	7'h1a :
		TR_193 = TR_84 ;
	7'h1b :
		TR_193 = TR_84 ;
	7'h1c :
		TR_193 = TR_84 ;
	7'h1d :
		TR_193 = TR_84 ;
	7'h1e :
		TR_193 = TR_84 ;
	7'h1f :
		TR_193 = TR_84 ;
	7'h20 :
		TR_193 = TR_84 ;
	7'h21 :
		TR_193 = TR_84 ;
	7'h22 :
		TR_193 = TR_84 ;
	7'h23 :
		TR_193 = TR_84 ;
	7'h24 :
		TR_193 = TR_84 ;
	7'h25 :
		TR_193 = TR_84 ;
	7'h26 :
		TR_193 = TR_84 ;
	7'h27 :
		TR_193 = TR_84 ;
	7'h28 :
		TR_193 = TR_84 ;
	7'h29 :
		TR_193 = TR_84 ;
	7'h2a :
		TR_193 = TR_84 ;
	7'h2b :
		TR_193 = TR_84 ;
	7'h2c :
		TR_193 = TR_84 ;
	7'h2d :
		TR_193 = TR_84 ;
	7'h2e :
		TR_193 = TR_84 ;
	7'h2f :
		TR_193 = TR_84 ;
	7'h30 :
		TR_193 = TR_84 ;
	7'h31 :
		TR_193 = TR_84 ;
	7'h32 :
		TR_193 = TR_84 ;
	7'h33 :
		TR_193 = TR_84 ;
	7'h34 :
		TR_193 = TR_84 ;
	7'h35 :
		TR_193 = TR_84 ;
	7'h36 :
		TR_193 = TR_84 ;
	7'h37 :
		TR_193 = TR_84 ;
	7'h38 :
		TR_193 = TR_84 ;
	7'h39 :
		TR_193 = TR_84 ;
	7'h3a :
		TR_193 = TR_84 ;
	7'h3b :
		TR_193 = TR_84 ;
	7'h3c :
		TR_193 = TR_84 ;
	7'h3d :
		TR_193 = TR_84 ;
	7'h3e :
		TR_193 = TR_84 ;
	7'h3f :
		TR_193 = TR_84 ;
	7'h40 :
		TR_193 = TR_84 ;
	7'h41 :
		TR_193 = TR_84 ;
	7'h42 :
		TR_193 = TR_84 ;
	7'h43 :
		TR_193 = TR_84 ;
	7'h44 :
		TR_193 = TR_84 ;
	7'h45 :
		TR_193 = TR_84 ;
	7'h46 :
		TR_193 = TR_84 ;
	7'h47 :
		TR_193 = TR_84 ;
	7'h48 :
		TR_193 = 9'h000 ;	// line#=../rle.cpp:80
	7'h49 :
		TR_193 = TR_84 ;
	7'h4a :
		TR_193 = TR_84 ;
	7'h4b :
		TR_193 = TR_84 ;
	7'h4c :
		TR_193 = TR_84 ;
	7'h4d :
		TR_193 = TR_84 ;
	7'h4e :
		TR_193 = TR_84 ;
	7'h4f :
		TR_193 = TR_84 ;
	7'h50 :
		TR_193 = TR_84 ;
	7'h51 :
		TR_193 = TR_84 ;
	7'h52 :
		TR_193 = TR_84 ;
	7'h53 :
		TR_193 = TR_84 ;
	7'h54 :
		TR_193 = TR_84 ;
	7'h55 :
		TR_193 = TR_84 ;
	7'h56 :
		TR_193 = TR_84 ;
	7'h57 :
		TR_193 = TR_84 ;
	7'h58 :
		TR_193 = TR_84 ;
	7'h59 :
		TR_193 = TR_84 ;
	7'h5a :
		TR_193 = TR_84 ;
	7'h5b :
		TR_193 = TR_84 ;
	7'h5c :
		TR_193 = TR_84 ;
	7'h5d :
		TR_193 = TR_84 ;
	7'h5e :
		TR_193 = TR_84 ;
	7'h5f :
		TR_193 = TR_84 ;
	7'h60 :
		TR_193 = TR_84 ;
	7'h61 :
		TR_193 = TR_84 ;
	7'h62 :
		TR_193 = TR_84 ;
	7'h63 :
		TR_193 = TR_84 ;
	7'h64 :
		TR_193 = TR_84 ;
	7'h65 :
		TR_193 = TR_84 ;
	7'h66 :
		TR_193 = TR_84 ;
	7'h67 :
		TR_193 = TR_84 ;
	7'h68 :
		TR_193 = TR_84 ;
	7'h69 :
		TR_193 = TR_84 ;
	7'h6a :
		TR_193 = TR_84 ;
	7'h6b :
		TR_193 = TR_84 ;
	7'h6c :
		TR_193 = TR_84 ;
	7'h6d :
		TR_193 = TR_84 ;
	7'h6e :
		TR_193 = TR_84 ;
	7'h6f :
		TR_193 = TR_84 ;
	7'h70 :
		TR_193 = TR_84 ;
	7'h71 :
		TR_193 = TR_84 ;
	7'h72 :
		TR_193 = TR_84 ;
	7'h73 :
		TR_193 = TR_84 ;
	7'h74 :
		TR_193 = TR_84 ;
	7'h75 :
		TR_193 = TR_84 ;
	7'h76 :
		TR_193 = TR_84 ;
	7'h77 :
		TR_193 = TR_84 ;
	7'h78 :
		TR_193 = TR_84 ;
	7'h79 :
		TR_193 = TR_84 ;
	7'h7a :
		TR_193 = TR_84 ;
	7'h7b :
		TR_193 = TR_84 ;
	7'h7c :
		TR_193 = TR_84 ;
	7'h7d :
		TR_193 = TR_84 ;
	7'h7e :
		TR_193 = TR_84 ;
	7'h7f :
		TR_193 = TR_84 ;
	default :
		TR_193 = 9'hx ;
	endcase
always @ ( TR_193 or U_173 or sub8u_71ot or U_183 or RG_rl_165 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_72_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h48 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_72_t = ( ( { 9{ M_180 } } & RG_rl_165 )
		| ( { 9{ U_173 } } & TR_193 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_72_en = ( M_180 | RG_rl_72_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_72_en )
		RG_rl_72 <= RG_rl_72_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_85 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_192 = TR_85 ;
	7'h01 :
		TR_192 = TR_85 ;
	7'h02 :
		TR_192 = TR_85 ;
	7'h03 :
		TR_192 = TR_85 ;
	7'h04 :
		TR_192 = TR_85 ;
	7'h05 :
		TR_192 = TR_85 ;
	7'h06 :
		TR_192 = TR_85 ;
	7'h07 :
		TR_192 = TR_85 ;
	7'h08 :
		TR_192 = TR_85 ;
	7'h09 :
		TR_192 = TR_85 ;
	7'h0a :
		TR_192 = TR_85 ;
	7'h0b :
		TR_192 = TR_85 ;
	7'h0c :
		TR_192 = TR_85 ;
	7'h0d :
		TR_192 = TR_85 ;
	7'h0e :
		TR_192 = TR_85 ;
	7'h0f :
		TR_192 = TR_85 ;
	7'h10 :
		TR_192 = TR_85 ;
	7'h11 :
		TR_192 = TR_85 ;
	7'h12 :
		TR_192 = TR_85 ;
	7'h13 :
		TR_192 = TR_85 ;
	7'h14 :
		TR_192 = TR_85 ;
	7'h15 :
		TR_192 = TR_85 ;
	7'h16 :
		TR_192 = TR_85 ;
	7'h17 :
		TR_192 = TR_85 ;
	7'h18 :
		TR_192 = TR_85 ;
	7'h19 :
		TR_192 = TR_85 ;
	7'h1a :
		TR_192 = TR_85 ;
	7'h1b :
		TR_192 = TR_85 ;
	7'h1c :
		TR_192 = TR_85 ;
	7'h1d :
		TR_192 = TR_85 ;
	7'h1e :
		TR_192 = TR_85 ;
	7'h1f :
		TR_192 = TR_85 ;
	7'h20 :
		TR_192 = TR_85 ;
	7'h21 :
		TR_192 = TR_85 ;
	7'h22 :
		TR_192 = TR_85 ;
	7'h23 :
		TR_192 = TR_85 ;
	7'h24 :
		TR_192 = TR_85 ;
	7'h25 :
		TR_192 = TR_85 ;
	7'h26 :
		TR_192 = TR_85 ;
	7'h27 :
		TR_192 = TR_85 ;
	7'h28 :
		TR_192 = TR_85 ;
	7'h29 :
		TR_192 = TR_85 ;
	7'h2a :
		TR_192 = TR_85 ;
	7'h2b :
		TR_192 = TR_85 ;
	7'h2c :
		TR_192 = TR_85 ;
	7'h2d :
		TR_192 = TR_85 ;
	7'h2e :
		TR_192 = TR_85 ;
	7'h2f :
		TR_192 = TR_85 ;
	7'h30 :
		TR_192 = TR_85 ;
	7'h31 :
		TR_192 = TR_85 ;
	7'h32 :
		TR_192 = TR_85 ;
	7'h33 :
		TR_192 = TR_85 ;
	7'h34 :
		TR_192 = TR_85 ;
	7'h35 :
		TR_192 = TR_85 ;
	7'h36 :
		TR_192 = TR_85 ;
	7'h37 :
		TR_192 = TR_85 ;
	7'h38 :
		TR_192 = TR_85 ;
	7'h39 :
		TR_192 = TR_85 ;
	7'h3a :
		TR_192 = TR_85 ;
	7'h3b :
		TR_192 = TR_85 ;
	7'h3c :
		TR_192 = TR_85 ;
	7'h3d :
		TR_192 = TR_85 ;
	7'h3e :
		TR_192 = TR_85 ;
	7'h3f :
		TR_192 = TR_85 ;
	7'h40 :
		TR_192 = TR_85 ;
	7'h41 :
		TR_192 = TR_85 ;
	7'h42 :
		TR_192 = TR_85 ;
	7'h43 :
		TR_192 = TR_85 ;
	7'h44 :
		TR_192 = TR_85 ;
	7'h45 :
		TR_192 = TR_85 ;
	7'h46 :
		TR_192 = TR_85 ;
	7'h47 :
		TR_192 = TR_85 ;
	7'h48 :
		TR_192 = TR_85 ;
	7'h49 :
		TR_192 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4a :
		TR_192 = TR_85 ;
	7'h4b :
		TR_192 = TR_85 ;
	7'h4c :
		TR_192 = TR_85 ;
	7'h4d :
		TR_192 = TR_85 ;
	7'h4e :
		TR_192 = TR_85 ;
	7'h4f :
		TR_192 = TR_85 ;
	7'h50 :
		TR_192 = TR_85 ;
	7'h51 :
		TR_192 = TR_85 ;
	7'h52 :
		TR_192 = TR_85 ;
	7'h53 :
		TR_192 = TR_85 ;
	7'h54 :
		TR_192 = TR_85 ;
	7'h55 :
		TR_192 = TR_85 ;
	7'h56 :
		TR_192 = TR_85 ;
	7'h57 :
		TR_192 = TR_85 ;
	7'h58 :
		TR_192 = TR_85 ;
	7'h59 :
		TR_192 = TR_85 ;
	7'h5a :
		TR_192 = TR_85 ;
	7'h5b :
		TR_192 = TR_85 ;
	7'h5c :
		TR_192 = TR_85 ;
	7'h5d :
		TR_192 = TR_85 ;
	7'h5e :
		TR_192 = TR_85 ;
	7'h5f :
		TR_192 = TR_85 ;
	7'h60 :
		TR_192 = TR_85 ;
	7'h61 :
		TR_192 = TR_85 ;
	7'h62 :
		TR_192 = TR_85 ;
	7'h63 :
		TR_192 = TR_85 ;
	7'h64 :
		TR_192 = TR_85 ;
	7'h65 :
		TR_192 = TR_85 ;
	7'h66 :
		TR_192 = TR_85 ;
	7'h67 :
		TR_192 = TR_85 ;
	7'h68 :
		TR_192 = TR_85 ;
	7'h69 :
		TR_192 = TR_85 ;
	7'h6a :
		TR_192 = TR_85 ;
	7'h6b :
		TR_192 = TR_85 ;
	7'h6c :
		TR_192 = TR_85 ;
	7'h6d :
		TR_192 = TR_85 ;
	7'h6e :
		TR_192 = TR_85 ;
	7'h6f :
		TR_192 = TR_85 ;
	7'h70 :
		TR_192 = TR_85 ;
	7'h71 :
		TR_192 = TR_85 ;
	7'h72 :
		TR_192 = TR_85 ;
	7'h73 :
		TR_192 = TR_85 ;
	7'h74 :
		TR_192 = TR_85 ;
	7'h75 :
		TR_192 = TR_85 ;
	7'h76 :
		TR_192 = TR_85 ;
	7'h77 :
		TR_192 = TR_85 ;
	7'h78 :
		TR_192 = TR_85 ;
	7'h79 :
		TR_192 = TR_85 ;
	7'h7a :
		TR_192 = TR_85 ;
	7'h7b :
		TR_192 = TR_85 ;
	7'h7c :
		TR_192 = TR_85 ;
	7'h7d :
		TR_192 = TR_85 ;
	7'h7e :
		TR_192 = TR_85 ;
	7'h7f :
		TR_192 = TR_85 ;
	default :
		TR_192 = 9'hx ;
	endcase
always @ ( TR_192 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_34 or 
	U_174 or RG_rl_165 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_73_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h49 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_73_t = ( ( { 9{ ST1_03d } } & RG_rl_165 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_34 )
		| ( { 9{ U_173 } } & TR_192 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_73_en = ( ST1_03d | U_174 | RG_rl_73_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_73_en )
		RG_rl_73 <= RG_rl_73_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_86 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_191 = TR_86 ;
	7'h01 :
		TR_191 = TR_86 ;
	7'h02 :
		TR_191 = TR_86 ;
	7'h03 :
		TR_191 = TR_86 ;
	7'h04 :
		TR_191 = TR_86 ;
	7'h05 :
		TR_191 = TR_86 ;
	7'h06 :
		TR_191 = TR_86 ;
	7'h07 :
		TR_191 = TR_86 ;
	7'h08 :
		TR_191 = TR_86 ;
	7'h09 :
		TR_191 = TR_86 ;
	7'h0a :
		TR_191 = TR_86 ;
	7'h0b :
		TR_191 = TR_86 ;
	7'h0c :
		TR_191 = TR_86 ;
	7'h0d :
		TR_191 = TR_86 ;
	7'h0e :
		TR_191 = TR_86 ;
	7'h0f :
		TR_191 = TR_86 ;
	7'h10 :
		TR_191 = TR_86 ;
	7'h11 :
		TR_191 = TR_86 ;
	7'h12 :
		TR_191 = TR_86 ;
	7'h13 :
		TR_191 = TR_86 ;
	7'h14 :
		TR_191 = TR_86 ;
	7'h15 :
		TR_191 = TR_86 ;
	7'h16 :
		TR_191 = TR_86 ;
	7'h17 :
		TR_191 = TR_86 ;
	7'h18 :
		TR_191 = TR_86 ;
	7'h19 :
		TR_191 = TR_86 ;
	7'h1a :
		TR_191 = TR_86 ;
	7'h1b :
		TR_191 = TR_86 ;
	7'h1c :
		TR_191 = TR_86 ;
	7'h1d :
		TR_191 = TR_86 ;
	7'h1e :
		TR_191 = TR_86 ;
	7'h1f :
		TR_191 = TR_86 ;
	7'h20 :
		TR_191 = TR_86 ;
	7'h21 :
		TR_191 = TR_86 ;
	7'h22 :
		TR_191 = TR_86 ;
	7'h23 :
		TR_191 = TR_86 ;
	7'h24 :
		TR_191 = TR_86 ;
	7'h25 :
		TR_191 = TR_86 ;
	7'h26 :
		TR_191 = TR_86 ;
	7'h27 :
		TR_191 = TR_86 ;
	7'h28 :
		TR_191 = TR_86 ;
	7'h29 :
		TR_191 = TR_86 ;
	7'h2a :
		TR_191 = TR_86 ;
	7'h2b :
		TR_191 = TR_86 ;
	7'h2c :
		TR_191 = TR_86 ;
	7'h2d :
		TR_191 = TR_86 ;
	7'h2e :
		TR_191 = TR_86 ;
	7'h2f :
		TR_191 = TR_86 ;
	7'h30 :
		TR_191 = TR_86 ;
	7'h31 :
		TR_191 = TR_86 ;
	7'h32 :
		TR_191 = TR_86 ;
	7'h33 :
		TR_191 = TR_86 ;
	7'h34 :
		TR_191 = TR_86 ;
	7'h35 :
		TR_191 = TR_86 ;
	7'h36 :
		TR_191 = TR_86 ;
	7'h37 :
		TR_191 = TR_86 ;
	7'h38 :
		TR_191 = TR_86 ;
	7'h39 :
		TR_191 = TR_86 ;
	7'h3a :
		TR_191 = TR_86 ;
	7'h3b :
		TR_191 = TR_86 ;
	7'h3c :
		TR_191 = TR_86 ;
	7'h3d :
		TR_191 = TR_86 ;
	7'h3e :
		TR_191 = TR_86 ;
	7'h3f :
		TR_191 = TR_86 ;
	7'h40 :
		TR_191 = TR_86 ;
	7'h41 :
		TR_191 = TR_86 ;
	7'h42 :
		TR_191 = TR_86 ;
	7'h43 :
		TR_191 = TR_86 ;
	7'h44 :
		TR_191 = TR_86 ;
	7'h45 :
		TR_191 = TR_86 ;
	7'h46 :
		TR_191 = TR_86 ;
	7'h47 :
		TR_191 = TR_86 ;
	7'h48 :
		TR_191 = TR_86 ;
	7'h49 :
		TR_191 = TR_86 ;
	7'h4a :
		TR_191 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4b :
		TR_191 = TR_86 ;
	7'h4c :
		TR_191 = TR_86 ;
	7'h4d :
		TR_191 = TR_86 ;
	7'h4e :
		TR_191 = TR_86 ;
	7'h4f :
		TR_191 = TR_86 ;
	7'h50 :
		TR_191 = TR_86 ;
	7'h51 :
		TR_191 = TR_86 ;
	7'h52 :
		TR_191 = TR_86 ;
	7'h53 :
		TR_191 = TR_86 ;
	7'h54 :
		TR_191 = TR_86 ;
	7'h55 :
		TR_191 = TR_86 ;
	7'h56 :
		TR_191 = TR_86 ;
	7'h57 :
		TR_191 = TR_86 ;
	7'h58 :
		TR_191 = TR_86 ;
	7'h59 :
		TR_191 = TR_86 ;
	7'h5a :
		TR_191 = TR_86 ;
	7'h5b :
		TR_191 = TR_86 ;
	7'h5c :
		TR_191 = TR_86 ;
	7'h5d :
		TR_191 = TR_86 ;
	7'h5e :
		TR_191 = TR_86 ;
	7'h5f :
		TR_191 = TR_86 ;
	7'h60 :
		TR_191 = TR_86 ;
	7'h61 :
		TR_191 = TR_86 ;
	7'h62 :
		TR_191 = TR_86 ;
	7'h63 :
		TR_191 = TR_86 ;
	7'h64 :
		TR_191 = TR_86 ;
	7'h65 :
		TR_191 = TR_86 ;
	7'h66 :
		TR_191 = TR_86 ;
	7'h67 :
		TR_191 = TR_86 ;
	7'h68 :
		TR_191 = TR_86 ;
	7'h69 :
		TR_191 = TR_86 ;
	7'h6a :
		TR_191 = TR_86 ;
	7'h6b :
		TR_191 = TR_86 ;
	7'h6c :
		TR_191 = TR_86 ;
	7'h6d :
		TR_191 = TR_86 ;
	7'h6e :
		TR_191 = TR_86 ;
	7'h6f :
		TR_191 = TR_86 ;
	7'h70 :
		TR_191 = TR_86 ;
	7'h71 :
		TR_191 = TR_86 ;
	7'h72 :
		TR_191 = TR_86 ;
	7'h73 :
		TR_191 = TR_86 ;
	7'h74 :
		TR_191 = TR_86 ;
	7'h75 :
		TR_191 = TR_86 ;
	7'h76 :
		TR_191 = TR_86 ;
	7'h77 :
		TR_191 = TR_86 ;
	7'h78 :
		TR_191 = TR_86 ;
	7'h79 :
		TR_191 = TR_86 ;
	7'h7a :
		TR_191 = TR_86 ;
	7'h7b :
		TR_191 = TR_86 ;
	7'h7c :
		TR_191 = TR_86 ;
	7'h7d :
		TR_191 = TR_86 ;
	7'h7e :
		TR_191 = TR_86 ;
	7'h7f :
		TR_191 = TR_86 ;
	default :
		TR_191 = 9'hx ;
	endcase
always @ ( TR_191 or U_173 or sub8u_71ot or U_183 or RG_rl_166 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_74_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h4a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_74_t = ( ( { 9{ M_180 } } & RG_rl_166 )
		| ( { 9{ U_173 } } & TR_191 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_74_en = ( M_180 | RG_rl_74_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_74_en )
		RG_rl_74 <= RG_rl_74_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_87 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_190 = TR_87 ;
	7'h01 :
		TR_190 = TR_87 ;
	7'h02 :
		TR_190 = TR_87 ;
	7'h03 :
		TR_190 = TR_87 ;
	7'h04 :
		TR_190 = TR_87 ;
	7'h05 :
		TR_190 = TR_87 ;
	7'h06 :
		TR_190 = TR_87 ;
	7'h07 :
		TR_190 = TR_87 ;
	7'h08 :
		TR_190 = TR_87 ;
	7'h09 :
		TR_190 = TR_87 ;
	7'h0a :
		TR_190 = TR_87 ;
	7'h0b :
		TR_190 = TR_87 ;
	7'h0c :
		TR_190 = TR_87 ;
	7'h0d :
		TR_190 = TR_87 ;
	7'h0e :
		TR_190 = TR_87 ;
	7'h0f :
		TR_190 = TR_87 ;
	7'h10 :
		TR_190 = TR_87 ;
	7'h11 :
		TR_190 = TR_87 ;
	7'h12 :
		TR_190 = TR_87 ;
	7'h13 :
		TR_190 = TR_87 ;
	7'h14 :
		TR_190 = TR_87 ;
	7'h15 :
		TR_190 = TR_87 ;
	7'h16 :
		TR_190 = TR_87 ;
	7'h17 :
		TR_190 = TR_87 ;
	7'h18 :
		TR_190 = TR_87 ;
	7'h19 :
		TR_190 = TR_87 ;
	7'h1a :
		TR_190 = TR_87 ;
	7'h1b :
		TR_190 = TR_87 ;
	7'h1c :
		TR_190 = TR_87 ;
	7'h1d :
		TR_190 = TR_87 ;
	7'h1e :
		TR_190 = TR_87 ;
	7'h1f :
		TR_190 = TR_87 ;
	7'h20 :
		TR_190 = TR_87 ;
	7'h21 :
		TR_190 = TR_87 ;
	7'h22 :
		TR_190 = TR_87 ;
	7'h23 :
		TR_190 = TR_87 ;
	7'h24 :
		TR_190 = TR_87 ;
	7'h25 :
		TR_190 = TR_87 ;
	7'h26 :
		TR_190 = TR_87 ;
	7'h27 :
		TR_190 = TR_87 ;
	7'h28 :
		TR_190 = TR_87 ;
	7'h29 :
		TR_190 = TR_87 ;
	7'h2a :
		TR_190 = TR_87 ;
	7'h2b :
		TR_190 = TR_87 ;
	7'h2c :
		TR_190 = TR_87 ;
	7'h2d :
		TR_190 = TR_87 ;
	7'h2e :
		TR_190 = TR_87 ;
	7'h2f :
		TR_190 = TR_87 ;
	7'h30 :
		TR_190 = TR_87 ;
	7'h31 :
		TR_190 = TR_87 ;
	7'h32 :
		TR_190 = TR_87 ;
	7'h33 :
		TR_190 = TR_87 ;
	7'h34 :
		TR_190 = TR_87 ;
	7'h35 :
		TR_190 = TR_87 ;
	7'h36 :
		TR_190 = TR_87 ;
	7'h37 :
		TR_190 = TR_87 ;
	7'h38 :
		TR_190 = TR_87 ;
	7'h39 :
		TR_190 = TR_87 ;
	7'h3a :
		TR_190 = TR_87 ;
	7'h3b :
		TR_190 = TR_87 ;
	7'h3c :
		TR_190 = TR_87 ;
	7'h3d :
		TR_190 = TR_87 ;
	7'h3e :
		TR_190 = TR_87 ;
	7'h3f :
		TR_190 = TR_87 ;
	7'h40 :
		TR_190 = TR_87 ;
	7'h41 :
		TR_190 = TR_87 ;
	7'h42 :
		TR_190 = TR_87 ;
	7'h43 :
		TR_190 = TR_87 ;
	7'h44 :
		TR_190 = TR_87 ;
	7'h45 :
		TR_190 = TR_87 ;
	7'h46 :
		TR_190 = TR_87 ;
	7'h47 :
		TR_190 = TR_87 ;
	7'h48 :
		TR_190 = TR_87 ;
	7'h49 :
		TR_190 = TR_87 ;
	7'h4a :
		TR_190 = TR_87 ;
	7'h4b :
		TR_190 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4c :
		TR_190 = TR_87 ;
	7'h4d :
		TR_190 = TR_87 ;
	7'h4e :
		TR_190 = TR_87 ;
	7'h4f :
		TR_190 = TR_87 ;
	7'h50 :
		TR_190 = TR_87 ;
	7'h51 :
		TR_190 = TR_87 ;
	7'h52 :
		TR_190 = TR_87 ;
	7'h53 :
		TR_190 = TR_87 ;
	7'h54 :
		TR_190 = TR_87 ;
	7'h55 :
		TR_190 = TR_87 ;
	7'h56 :
		TR_190 = TR_87 ;
	7'h57 :
		TR_190 = TR_87 ;
	7'h58 :
		TR_190 = TR_87 ;
	7'h59 :
		TR_190 = TR_87 ;
	7'h5a :
		TR_190 = TR_87 ;
	7'h5b :
		TR_190 = TR_87 ;
	7'h5c :
		TR_190 = TR_87 ;
	7'h5d :
		TR_190 = TR_87 ;
	7'h5e :
		TR_190 = TR_87 ;
	7'h5f :
		TR_190 = TR_87 ;
	7'h60 :
		TR_190 = TR_87 ;
	7'h61 :
		TR_190 = TR_87 ;
	7'h62 :
		TR_190 = TR_87 ;
	7'h63 :
		TR_190 = TR_87 ;
	7'h64 :
		TR_190 = TR_87 ;
	7'h65 :
		TR_190 = TR_87 ;
	7'h66 :
		TR_190 = TR_87 ;
	7'h67 :
		TR_190 = TR_87 ;
	7'h68 :
		TR_190 = TR_87 ;
	7'h69 :
		TR_190 = TR_87 ;
	7'h6a :
		TR_190 = TR_87 ;
	7'h6b :
		TR_190 = TR_87 ;
	7'h6c :
		TR_190 = TR_87 ;
	7'h6d :
		TR_190 = TR_87 ;
	7'h6e :
		TR_190 = TR_87 ;
	7'h6f :
		TR_190 = TR_87 ;
	7'h70 :
		TR_190 = TR_87 ;
	7'h71 :
		TR_190 = TR_87 ;
	7'h72 :
		TR_190 = TR_87 ;
	7'h73 :
		TR_190 = TR_87 ;
	7'h74 :
		TR_190 = TR_87 ;
	7'h75 :
		TR_190 = TR_87 ;
	7'h76 :
		TR_190 = TR_87 ;
	7'h77 :
		TR_190 = TR_87 ;
	7'h78 :
		TR_190 = TR_87 ;
	7'h79 :
		TR_190 = TR_87 ;
	7'h7a :
		TR_190 = TR_87 ;
	7'h7b :
		TR_190 = TR_87 ;
	7'h7c :
		TR_190 = TR_87 ;
	7'h7d :
		TR_190 = TR_87 ;
	7'h7e :
		TR_190 = TR_87 ;
	7'h7f :
		TR_190 = TR_87 ;
	default :
		TR_190 = 9'hx ;
	endcase
always @ ( TR_190 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_35 or 
	U_174 or RG_rl_166 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_75_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h4b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_75_t = ( ( { 9{ ST1_03d } } & RG_rl_166 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_35 )
		| ( { 9{ U_173 } } & TR_190 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_75_en = ( ST1_03d | U_174 | RG_rl_75_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_75_en )
		RG_rl_75 <= RG_rl_75_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_88 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_189 = TR_88 ;
	7'h01 :
		TR_189 = TR_88 ;
	7'h02 :
		TR_189 = TR_88 ;
	7'h03 :
		TR_189 = TR_88 ;
	7'h04 :
		TR_189 = TR_88 ;
	7'h05 :
		TR_189 = TR_88 ;
	7'h06 :
		TR_189 = TR_88 ;
	7'h07 :
		TR_189 = TR_88 ;
	7'h08 :
		TR_189 = TR_88 ;
	7'h09 :
		TR_189 = TR_88 ;
	7'h0a :
		TR_189 = TR_88 ;
	7'h0b :
		TR_189 = TR_88 ;
	7'h0c :
		TR_189 = TR_88 ;
	7'h0d :
		TR_189 = TR_88 ;
	7'h0e :
		TR_189 = TR_88 ;
	7'h0f :
		TR_189 = TR_88 ;
	7'h10 :
		TR_189 = TR_88 ;
	7'h11 :
		TR_189 = TR_88 ;
	7'h12 :
		TR_189 = TR_88 ;
	7'h13 :
		TR_189 = TR_88 ;
	7'h14 :
		TR_189 = TR_88 ;
	7'h15 :
		TR_189 = TR_88 ;
	7'h16 :
		TR_189 = TR_88 ;
	7'h17 :
		TR_189 = TR_88 ;
	7'h18 :
		TR_189 = TR_88 ;
	7'h19 :
		TR_189 = TR_88 ;
	7'h1a :
		TR_189 = TR_88 ;
	7'h1b :
		TR_189 = TR_88 ;
	7'h1c :
		TR_189 = TR_88 ;
	7'h1d :
		TR_189 = TR_88 ;
	7'h1e :
		TR_189 = TR_88 ;
	7'h1f :
		TR_189 = TR_88 ;
	7'h20 :
		TR_189 = TR_88 ;
	7'h21 :
		TR_189 = TR_88 ;
	7'h22 :
		TR_189 = TR_88 ;
	7'h23 :
		TR_189 = TR_88 ;
	7'h24 :
		TR_189 = TR_88 ;
	7'h25 :
		TR_189 = TR_88 ;
	7'h26 :
		TR_189 = TR_88 ;
	7'h27 :
		TR_189 = TR_88 ;
	7'h28 :
		TR_189 = TR_88 ;
	7'h29 :
		TR_189 = TR_88 ;
	7'h2a :
		TR_189 = TR_88 ;
	7'h2b :
		TR_189 = TR_88 ;
	7'h2c :
		TR_189 = TR_88 ;
	7'h2d :
		TR_189 = TR_88 ;
	7'h2e :
		TR_189 = TR_88 ;
	7'h2f :
		TR_189 = TR_88 ;
	7'h30 :
		TR_189 = TR_88 ;
	7'h31 :
		TR_189 = TR_88 ;
	7'h32 :
		TR_189 = TR_88 ;
	7'h33 :
		TR_189 = TR_88 ;
	7'h34 :
		TR_189 = TR_88 ;
	7'h35 :
		TR_189 = TR_88 ;
	7'h36 :
		TR_189 = TR_88 ;
	7'h37 :
		TR_189 = TR_88 ;
	7'h38 :
		TR_189 = TR_88 ;
	7'h39 :
		TR_189 = TR_88 ;
	7'h3a :
		TR_189 = TR_88 ;
	7'h3b :
		TR_189 = TR_88 ;
	7'h3c :
		TR_189 = TR_88 ;
	7'h3d :
		TR_189 = TR_88 ;
	7'h3e :
		TR_189 = TR_88 ;
	7'h3f :
		TR_189 = TR_88 ;
	7'h40 :
		TR_189 = TR_88 ;
	7'h41 :
		TR_189 = TR_88 ;
	7'h42 :
		TR_189 = TR_88 ;
	7'h43 :
		TR_189 = TR_88 ;
	7'h44 :
		TR_189 = TR_88 ;
	7'h45 :
		TR_189 = TR_88 ;
	7'h46 :
		TR_189 = TR_88 ;
	7'h47 :
		TR_189 = TR_88 ;
	7'h48 :
		TR_189 = TR_88 ;
	7'h49 :
		TR_189 = TR_88 ;
	7'h4a :
		TR_189 = TR_88 ;
	7'h4b :
		TR_189 = TR_88 ;
	7'h4c :
		TR_189 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4d :
		TR_189 = TR_88 ;
	7'h4e :
		TR_189 = TR_88 ;
	7'h4f :
		TR_189 = TR_88 ;
	7'h50 :
		TR_189 = TR_88 ;
	7'h51 :
		TR_189 = TR_88 ;
	7'h52 :
		TR_189 = TR_88 ;
	7'h53 :
		TR_189 = TR_88 ;
	7'h54 :
		TR_189 = TR_88 ;
	7'h55 :
		TR_189 = TR_88 ;
	7'h56 :
		TR_189 = TR_88 ;
	7'h57 :
		TR_189 = TR_88 ;
	7'h58 :
		TR_189 = TR_88 ;
	7'h59 :
		TR_189 = TR_88 ;
	7'h5a :
		TR_189 = TR_88 ;
	7'h5b :
		TR_189 = TR_88 ;
	7'h5c :
		TR_189 = TR_88 ;
	7'h5d :
		TR_189 = TR_88 ;
	7'h5e :
		TR_189 = TR_88 ;
	7'h5f :
		TR_189 = TR_88 ;
	7'h60 :
		TR_189 = TR_88 ;
	7'h61 :
		TR_189 = TR_88 ;
	7'h62 :
		TR_189 = TR_88 ;
	7'h63 :
		TR_189 = TR_88 ;
	7'h64 :
		TR_189 = TR_88 ;
	7'h65 :
		TR_189 = TR_88 ;
	7'h66 :
		TR_189 = TR_88 ;
	7'h67 :
		TR_189 = TR_88 ;
	7'h68 :
		TR_189 = TR_88 ;
	7'h69 :
		TR_189 = TR_88 ;
	7'h6a :
		TR_189 = TR_88 ;
	7'h6b :
		TR_189 = TR_88 ;
	7'h6c :
		TR_189 = TR_88 ;
	7'h6d :
		TR_189 = TR_88 ;
	7'h6e :
		TR_189 = TR_88 ;
	7'h6f :
		TR_189 = TR_88 ;
	7'h70 :
		TR_189 = TR_88 ;
	7'h71 :
		TR_189 = TR_88 ;
	7'h72 :
		TR_189 = TR_88 ;
	7'h73 :
		TR_189 = TR_88 ;
	7'h74 :
		TR_189 = TR_88 ;
	7'h75 :
		TR_189 = TR_88 ;
	7'h76 :
		TR_189 = TR_88 ;
	7'h77 :
		TR_189 = TR_88 ;
	7'h78 :
		TR_189 = TR_88 ;
	7'h79 :
		TR_189 = TR_88 ;
	7'h7a :
		TR_189 = TR_88 ;
	7'h7b :
		TR_189 = TR_88 ;
	7'h7c :
		TR_189 = TR_88 ;
	7'h7d :
		TR_189 = TR_88 ;
	7'h7e :
		TR_189 = TR_88 ;
	7'h7f :
		TR_189 = TR_88 ;
	default :
		TR_189 = 9'hx ;
	endcase
always @ ( TR_189 or U_173 or sub8u_71ot or U_183 or RG_rl_167 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_76_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h4c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_76_t = ( ( { 9{ M_180 } } & RG_rl_167 )
		| ( { 9{ U_173 } } & TR_189 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_76_en = ( M_180 | RG_rl_76_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_76_en )
		RG_rl_76 <= RG_rl_76_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_89 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_188 = TR_89 ;
	7'h01 :
		TR_188 = TR_89 ;
	7'h02 :
		TR_188 = TR_89 ;
	7'h03 :
		TR_188 = TR_89 ;
	7'h04 :
		TR_188 = TR_89 ;
	7'h05 :
		TR_188 = TR_89 ;
	7'h06 :
		TR_188 = TR_89 ;
	7'h07 :
		TR_188 = TR_89 ;
	7'h08 :
		TR_188 = TR_89 ;
	7'h09 :
		TR_188 = TR_89 ;
	7'h0a :
		TR_188 = TR_89 ;
	7'h0b :
		TR_188 = TR_89 ;
	7'h0c :
		TR_188 = TR_89 ;
	7'h0d :
		TR_188 = TR_89 ;
	7'h0e :
		TR_188 = TR_89 ;
	7'h0f :
		TR_188 = TR_89 ;
	7'h10 :
		TR_188 = TR_89 ;
	7'h11 :
		TR_188 = TR_89 ;
	7'h12 :
		TR_188 = TR_89 ;
	7'h13 :
		TR_188 = TR_89 ;
	7'h14 :
		TR_188 = TR_89 ;
	7'h15 :
		TR_188 = TR_89 ;
	7'h16 :
		TR_188 = TR_89 ;
	7'h17 :
		TR_188 = TR_89 ;
	7'h18 :
		TR_188 = TR_89 ;
	7'h19 :
		TR_188 = TR_89 ;
	7'h1a :
		TR_188 = TR_89 ;
	7'h1b :
		TR_188 = TR_89 ;
	7'h1c :
		TR_188 = TR_89 ;
	7'h1d :
		TR_188 = TR_89 ;
	7'h1e :
		TR_188 = TR_89 ;
	7'h1f :
		TR_188 = TR_89 ;
	7'h20 :
		TR_188 = TR_89 ;
	7'h21 :
		TR_188 = TR_89 ;
	7'h22 :
		TR_188 = TR_89 ;
	7'h23 :
		TR_188 = TR_89 ;
	7'h24 :
		TR_188 = TR_89 ;
	7'h25 :
		TR_188 = TR_89 ;
	7'h26 :
		TR_188 = TR_89 ;
	7'h27 :
		TR_188 = TR_89 ;
	7'h28 :
		TR_188 = TR_89 ;
	7'h29 :
		TR_188 = TR_89 ;
	7'h2a :
		TR_188 = TR_89 ;
	7'h2b :
		TR_188 = TR_89 ;
	7'h2c :
		TR_188 = TR_89 ;
	7'h2d :
		TR_188 = TR_89 ;
	7'h2e :
		TR_188 = TR_89 ;
	7'h2f :
		TR_188 = TR_89 ;
	7'h30 :
		TR_188 = TR_89 ;
	7'h31 :
		TR_188 = TR_89 ;
	7'h32 :
		TR_188 = TR_89 ;
	7'h33 :
		TR_188 = TR_89 ;
	7'h34 :
		TR_188 = TR_89 ;
	7'h35 :
		TR_188 = TR_89 ;
	7'h36 :
		TR_188 = TR_89 ;
	7'h37 :
		TR_188 = TR_89 ;
	7'h38 :
		TR_188 = TR_89 ;
	7'h39 :
		TR_188 = TR_89 ;
	7'h3a :
		TR_188 = TR_89 ;
	7'h3b :
		TR_188 = TR_89 ;
	7'h3c :
		TR_188 = TR_89 ;
	7'h3d :
		TR_188 = TR_89 ;
	7'h3e :
		TR_188 = TR_89 ;
	7'h3f :
		TR_188 = TR_89 ;
	7'h40 :
		TR_188 = TR_89 ;
	7'h41 :
		TR_188 = TR_89 ;
	7'h42 :
		TR_188 = TR_89 ;
	7'h43 :
		TR_188 = TR_89 ;
	7'h44 :
		TR_188 = TR_89 ;
	7'h45 :
		TR_188 = TR_89 ;
	7'h46 :
		TR_188 = TR_89 ;
	7'h47 :
		TR_188 = TR_89 ;
	7'h48 :
		TR_188 = TR_89 ;
	7'h49 :
		TR_188 = TR_89 ;
	7'h4a :
		TR_188 = TR_89 ;
	7'h4b :
		TR_188 = TR_89 ;
	7'h4c :
		TR_188 = TR_89 ;
	7'h4d :
		TR_188 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4e :
		TR_188 = TR_89 ;
	7'h4f :
		TR_188 = TR_89 ;
	7'h50 :
		TR_188 = TR_89 ;
	7'h51 :
		TR_188 = TR_89 ;
	7'h52 :
		TR_188 = TR_89 ;
	7'h53 :
		TR_188 = TR_89 ;
	7'h54 :
		TR_188 = TR_89 ;
	7'h55 :
		TR_188 = TR_89 ;
	7'h56 :
		TR_188 = TR_89 ;
	7'h57 :
		TR_188 = TR_89 ;
	7'h58 :
		TR_188 = TR_89 ;
	7'h59 :
		TR_188 = TR_89 ;
	7'h5a :
		TR_188 = TR_89 ;
	7'h5b :
		TR_188 = TR_89 ;
	7'h5c :
		TR_188 = TR_89 ;
	7'h5d :
		TR_188 = TR_89 ;
	7'h5e :
		TR_188 = TR_89 ;
	7'h5f :
		TR_188 = TR_89 ;
	7'h60 :
		TR_188 = TR_89 ;
	7'h61 :
		TR_188 = TR_89 ;
	7'h62 :
		TR_188 = TR_89 ;
	7'h63 :
		TR_188 = TR_89 ;
	7'h64 :
		TR_188 = TR_89 ;
	7'h65 :
		TR_188 = TR_89 ;
	7'h66 :
		TR_188 = TR_89 ;
	7'h67 :
		TR_188 = TR_89 ;
	7'h68 :
		TR_188 = TR_89 ;
	7'h69 :
		TR_188 = TR_89 ;
	7'h6a :
		TR_188 = TR_89 ;
	7'h6b :
		TR_188 = TR_89 ;
	7'h6c :
		TR_188 = TR_89 ;
	7'h6d :
		TR_188 = TR_89 ;
	7'h6e :
		TR_188 = TR_89 ;
	7'h6f :
		TR_188 = TR_89 ;
	7'h70 :
		TR_188 = TR_89 ;
	7'h71 :
		TR_188 = TR_89 ;
	7'h72 :
		TR_188 = TR_89 ;
	7'h73 :
		TR_188 = TR_89 ;
	7'h74 :
		TR_188 = TR_89 ;
	7'h75 :
		TR_188 = TR_89 ;
	7'h76 :
		TR_188 = TR_89 ;
	7'h77 :
		TR_188 = TR_89 ;
	7'h78 :
		TR_188 = TR_89 ;
	7'h79 :
		TR_188 = TR_89 ;
	7'h7a :
		TR_188 = TR_89 ;
	7'h7b :
		TR_188 = TR_89 ;
	7'h7c :
		TR_188 = TR_89 ;
	7'h7d :
		TR_188 = TR_89 ;
	7'h7e :
		TR_188 = TR_89 ;
	7'h7f :
		TR_188 = TR_89 ;
	default :
		TR_188 = 9'hx ;
	endcase
always @ ( TR_188 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_36 or 
	U_174 or RG_rl_167 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_77_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h4d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_77_t = ( ( { 9{ ST1_03d } } & RG_rl_167 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_36 )
		| ( { 9{ U_173 } } & TR_188 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_77_en = ( ST1_03d | U_174 | RG_rl_77_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_77_en )
		RG_rl_77 <= RG_rl_77_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_90 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_187 = TR_90 ;
	7'h01 :
		TR_187 = TR_90 ;
	7'h02 :
		TR_187 = TR_90 ;
	7'h03 :
		TR_187 = TR_90 ;
	7'h04 :
		TR_187 = TR_90 ;
	7'h05 :
		TR_187 = TR_90 ;
	7'h06 :
		TR_187 = TR_90 ;
	7'h07 :
		TR_187 = TR_90 ;
	7'h08 :
		TR_187 = TR_90 ;
	7'h09 :
		TR_187 = TR_90 ;
	7'h0a :
		TR_187 = TR_90 ;
	7'h0b :
		TR_187 = TR_90 ;
	7'h0c :
		TR_187 = TR_90 ;
	7'h0d :
		TR_187 = TR_90 ;
	7'h0e :
		TR_187 = TR_90 ;
	7'h0f :
		TR_187 = TR_90 ;
	7'h10 :
		TR_187 = TR_90 ;
	7'h11 :
		TR_187 = TR_90 ;
	7'h12 :
		TR_187 = TR_90 ;
	7'h13 :
		TR_187 = TR_90 ;
	7'h14 :
		TR_187 = TR_90 ;
	7'h15 :
		TR_187 = TR_90 ;
	7'h16 :
		TR_187 = TR_90 ;
	7'h17 :
		TR_187 = TR_90 ;
	7'h18 :
		TR_187 = TR_90 ;
	7'h19 :
		TR_187 = TR_90 ;
	7'h1a :
		TR_187 = TR_90 ;
	7'h1b :
		TR_187 = TR_90 ;
	7'h1c :
		TR_187 = TR_90 ;
	7'h1d :
		TR_187 = TR_90 ;
	7'h1e :
		TR_187 = TR_90 ;
	7'h1f :
		TR_187 = TR_90 ;
	7'h20 :
		TR_187 = TR_90 ;
	7'h21 :
		TR_187 = TR_90 ;
	7'h22 :
		TR_187 = TR_90 ;
	7'h23 :
		TR_187 = TR_90 ;
	7'h24 :
		TR_187 = TR_90 ;
	7'h25 :
		TR_187 = TR_90 ;
	7'h26 :
		TR_187 = TR_90 ;
	7'h27 :
		TR_187 = TR_90 ;
	7'h28 :
		TR_187 = TR_90 ;
	7'h29 :
		TR_187 = TR_90 ;
	7'h2a :
		TR_187 = TR_90 ;
	7'h2b :
		TR_187 = TR_90 ;
	7'h2c :
		TR_187 = TR_90 ;
	7'h2d :
		TR_187 = TR_90 ;
	7'h2e :
		TR_187 = TR_90 ;
	7'h2f :
		TR_187 = TR_90 ;
	7'h30 :
		TR_187 = TR_90 ;
	7'h31 :
		TR_187 = TR_90 ;
	7'h32 :
		TR_187 = TR_90 ;
	7'h33 :
		TR_187 = TR_90 ;
	7'h34 :
		TR_187 = TR_90 ;
	7'h35 :
		TR_187 = TR_90 ;
	7'h36 :
		TR_187 = TR_90 ;
	7'h37 :
		TR_187 = TR_90 ;
	7'h38 :
		TR_187 = TR_90 ;
	7'h39 :
		TR_187 = TR_90 ;
	7'h3a :
		TR_187 = TR_90 ;
	7'h3b :
		TR_187 = TR_90 ;
	7'h3c :
		TR_187 = TR_90 ;
	7'h3d :
		TR_187 = TR_90 ;
	7'h3e :
		TR_187 = TR_90 ;
	7'h3f :
		TR_187 = TR_90 ;
	7'h40 :
		TR_187 = TR_90 ;
	7'h41 :
		TR_187 = TR_90 ;
	7'h42 :
		TR_187 = TR_90 ;
	7'h43 :
		TR_187 = TR_90 ;
	7'h44 :
		TR_187 = TR_90 ;
	7'h45 :
		TR_187 = TR_90 ;
	7'h46 :
		TR_187 = TR_90 ;
	7'h47 :
		TR_187 = TR_90 ;
	7'h48 :
		TR_187 = TR_90 ;
	7'h49 :
		TR_187 = TR_90 ;
	7'h4a :
		TR_187 = TR_90 ;
	7'h4b :
		TR_187 = TR_90 ;
	7'h4c :
		TR_187 = TR_90 ;
	7'h4d :
		TR_187 = TR_90 ;
	7'h4e :
		TR_187 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4f :
		TR_187 = TR_90 ;
	7'h50 :
		TR_187 = TR_90 ;
	7'h51 :
		TR_187 = TR_90 ;
	7'h52 :
		TR_187 = TR_90 ;
	7'h53 :
		TR_187 = TR_90 ;
	7'h54 :
		TR_187 = TR_90 ;
	7'h55 :
		TR_187 = TR_90 ;
	7'h56 :
		TR_187 = TR_90 ;
	7'h57 :
		TR_187 = TR_90 ;
	7'h58 :
		TR_187 = TR_90 ;
	7'h59 :
		TR_187 = TR_90 ;
	7'h5a :
		TR_187 = TR_90 ;
	7'h5b :
		TR_187 = TR_90 ;
	7'h5c :
		TR_187 = TR_90 ;
	7'h5d :
		TR_187 = TR_90 ;
	7'h5e :
		TR_187 = TR_90 ;
	7'h5f :
		TR_187 = TR_90 ;
	7'h60 :
		TR_187 = TR_90 ;
	7'h61 :
		TR_187 = TR_90 ;
	7'h62 :
		TR_187 = TR_90 ;
	7'h63 :
		TR_187 = TR_90 ;
	7'h64 :
		TR_187 = TR_90 ;
	7'h65 :
		TR_187 = TR_90 ;
	7'h66 :
		TR_187 = TR_90 ;
	7'h67 :
		TR_187 = TR_90 ;
	7'h68 :
		TR_187 = TR_90 ;
	7'h69 :
		TR_187 = TR_90 ;
	7'h6a :
		TR_187 = TR_90 ;
	7'h6b :
		TR_187 = TR_90 ;
	7'h6c :
		TR_187 = TR_90 ;
	7'h6d :
		TR_187 = TR_90 ;
	7'h6e :
		TR_187 = TR_90 ;
	7'h6f :
		TR_187 = TR_90 ;
	7'h70 :
		TR_187 = TR_90 ;
	7'h71 :
		TR_187 = TR_90 ;
	7'h72 :
		TR_187 = TR_90 ;
	7'h73 :
		TR_187 = TR_90 ;
	7'h74 :
		TR_187 = TR_90 ;
	7'h75 :
		TR_187 = TR_90 ;
	7'h76 :
		TR_187 = TR_90 ;
	7'h77 :
		TR_187 = TR_90 ;
	7'h78 :
		TR_187 = TR_90 ;
	7'h79 :
		TR_187 = TR_90 ;
	7'h7a :
		TR_187 = TR_90 ;
	7'h7b :
		TR_187 = TR_90 ;
	7'h7c :
		TR_187 = TR_90 ;
	7'h7d :
		TR_187 = TR_90 ;
	7'h7e :
		TR_187 = TR_90 ;
	7'h7f :
		TR_187 = TR_90 ;
	default :
		TR_187 = 9'hx ;
	endcase
always @ ( TR_187 or U_173 or sub8u_71ot or U_183 or RG_rl_168 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_78_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h4e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_78_t = ( ( { 9{ M_180 } } & RG_rl_168 )
		| ( { 9{ U_173 } } & TR_187 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_78_en = ( M_180 | RG_rl_78_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_78_en )
		RG_rl_78 <= RG_rl_78_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_91 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_186 = TR_91 ;
	7'h01 :
		TR_186 = TR_91 ;
	7'h02 :
		TR_186 = TR_91 ;
	7'h03 :
		TR_186 = TR_91 ;
	7'h04 :
		TR_186 = TR_91 ;
	7'h05 :
		TR_186 = TR_91 ;
	7'h06 :
		TR_186 = TR_91 ;
	7'h07 :
		TR_186 = TR_91 ;
	7'h08 :
		TR_186 = TR_91 ;
	7'h09 :
		TR_186 = TR_91 ;
	7'h0a :
		TR_186 = TR_91 ;
	7'h0b :
		TR_186 = TR_91 ;
	7'h0c :
		TR_186 = TR_91 ;
	7'h0d :
		TR_186 = TR_91 ;
	7'h0e :
		TR_186 = TR_91 ;
	7'h0f :
		TR_186 = TR_91 ;
	7'h10 :
		TR_186 = TR_91 ;
	7'h11 :
		TR_186 = TR_91 ;
	7'h12 :
		TR_186 = TR_91 ;
	7'h13 :
		TR_186 = TR_91 ;
	7'h14 :
		TR_186 = TR_91 ;
	7'h15 :
		TR_186 = TR_91 ;
	7'h16 :
		TR_186 = TR_91 ;
	7'h17 :
		TR_186 = TR_91 ;
	7'h18 :
		TR_186 = TR_91 ;
	7'h19 :
		TR_186 = TR_91 ;
	7'h1a :
		TR_186 = TR_91 ;
	7'h1b :
		TR_186 = TR_91 ;
	7'h1c :
		TR_186 = TR_91 ;
	7'h1d :
		TR_186 = TR_91 ;
	7'h1e :
		TR_186 = TR_91 ;
	7'h1f :
		TR_186 = TR_91 ;
	7'h20 :
		TR_186 = TR_91 ;
	7'h21 :
		TR_186 = TR_91 ;
	7'h22 :
		TR_186 = TR_91 ;
	7'h23 :
		TR_186 = TR_91 ;
	7'h24 :
		TR_186 = TR_91 ;
	7'h25 :
		TR_186 = TR_91 ;
	7'h26 :
		TR_186 = TR_91 ;
	7'h27 :
		TR_186 = TR_91 ;
	7'h28 :
		TR_186 = TR_91 ;
	7'h29 :
		TR_186 = TR_91 ;
	7'h2a :
		TR_186 = TR_91 ;
	7'h2b :
		TR_186 = TR_91 ;
	7'h2c :
		TR_186 = TR_91 ;
	7'h2d :
		TR_186 = TR_91 ;
	7'h2e :
		TR_186 = TR_91 ;
	7'h2f :
		TR_186 = TR_91 ;
	7'h30 :
		TR_186 = TR_91 ;
	7'h31 :
		TR_186 = TR_91 ;
	7'h32 :
		TR_186 = TR_91 ;
	7'h33 :
		TR_186 = TR_91 ;
	7'h34 :
		TR_186 = TR_91 ;
	7'h35 :
		TR_186 = TR_91 ;
	7'h36 :
		TR_186 = TR_91 ;
	7'h37 :
		TR_186 = TR_91 ;
	7'h38 :
		TR_186 = TR_91 ;
	7'h39 :
		TR_186 = TR_91 ;
	7'h3a :
		TR_186 = TR_91 ;
	7'h3b :
		TR_186 = TR_91 ;
	7'h3c :
		TR_186 = TR_91 ;
	7'h3d :
		TR_186 = TR_91 ;
	7'h3e :
		TR_186 = TR_91 ;
	7'h3f :
		TR_186 = TR_91 ;
	7'h40 :
		TR_186 = TR_91 ;
	7'h41 :
		TR_186 = TR_91 ;
	7'h42 :
		TR_186 = TR_91 ;
	7'h43 :
		TR_186 = TR_91 ;
	7'h44 :
		TR_186 = TR_91 ;
	7'h45 :
		TR_186 = TR_91 ;
	7'h46 :
		TR_186 = TR_91 ;
	7'h47 :
		TR_186 = TR_91 ;
	7'h48 :
		TR_186 = TR_91 ;
	7'h49 :
		TR_186 = TR_91 ;
	7'h4a :
		TR_186 = TR_91 ;
	7'h4b :
		TR_186 = TR_91 ;
	7'h4c :
		TR_186 = TR_91 ;
	7'h4d :
		TR_186 = TR_91 ;
	7'h4e :
		TR_186 = TR_91 ;
	7'h4f :
		TR_186 = 9'h000 ;	// line#=../rle.cpp:80
	7'h50 :
		TR_186 = TR_91 ;
	7'h51 :
		TR_186 = TR_91 ;
	7'h52 :
		TR_186 = TR_91 ;
	7'h53 :
		TR_186 = TR_91 ;
	7'h54 :
		TR_186 = TR_91 ;
	7'h55 :
		TR_186 = TR_91 ;
	7'h56 :
		TR_186 = TR_91 ;
	7'h57 :
		TR_186 = TR_91 ;
	7'h58 :
		TR_186 = TR_91 ;
	7'h59 :
		TR_186 = TR_91 ;
	7'h5a :
		TR_186 = TR_91 ;
	7'h5b :
		TR_186 = TR_91 ;
	7'h5c :
		TR_186 = TR_91 ;
	7'h5d :
		TR_186 = TR_91 ;
	7'h5e :
		TR_186 = TR_91 ;
	7'h5f :
		TR_186 = TR_91 ;
	7'h60 :
		TR_186 = TR_91 ;
	7'h61 :
		TR_186 = TR_91 ;
	7'h62 :
		TR_186 = TR_91 ;
	7'h63 :
		TR_186 = TR_91 ;
	7'h64 :
		TR_186 = TR_91 ;
	7'h65 :
		TR_186 = TR_91 ;
	7'h66 :
		TR_186 = TR_91 ;
	7'h67 :
		TR_186 = TR_91 ;
	7'h68 :
		TR_186 = TR_91 ;
	7'h69 :
		TR_186 = TR_91 ;
	7'h6a :
		TR_186 = TR_91 ;
	7'h6b :
		TR_186 = TR_91 ;
	7'h6c :
		TR_186 = TR_91 ;
	7'h6d :
		TR_186 = TR_91 ;
	7'h6e :
		TR_186 = TR_91 ;
	7'h6f :
		TR_186 = TR_91 ;
	7'h70 :
		TR_186 = TR_91 ;
	7'h71 :
		TR_186 = TR_91 ;
	7'h72 :
		TR_186 = TR_91 ;
	7'h73 :
		TR_186 = TR_91 ;
	7'h74 :
		TR_186 = TR_91 ;
	7'h75 :
		TR_186 = TR_91 ;
	7'h76 :
		TR_186 = TR_91 ;
	7'h77 :
		TR_186 = TR_91 ;
	7'h78 :
		TR_186 = TR_91 ;
	7'h79 :
		TR_186 = TR_91 ;
	7'h7a :
		TR_186 = TR_91 ;
	7'h7b :
		TR_186 = TR_91 ;
	7'h7c :
		TR_186 = TR_91 ;
	7'h7d :
		TR_186 = TR_91 ;
	7'h7e :
		TR_186 = TR_91 ;
	7'h7f :
		TR_186 = TR_91 ;
	default :
		TR_186 = 9'hx ;
	endcase
always @ ( TR_186 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_37 or 
	U_174 or RG_rl_168 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_79_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h4f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_79_t = ( ( { 9{ ST1_03d } } & RG_rl_168 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_37 )
		| ( { 9{ U_173 } } & TR_186 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_79_en = ( ST1_03d | U_174 | RG_rl_79_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_79_en )
		RG_rl_79 <= RG_rl_79_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_92 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_185 = TR_92 ;
	7'h01 :
		TR_185 = TR_92 ;
	7'h02 :
		TR_185 = TR_92 ;
	7'h03 :
		TR_185 = TR_92 ;
	7'h04 :
		TR_185 = TR_92 ;
	7'h05 :
		TR_185 = TR_92 ;
	7'h06 :
		TR_185 = TR_92 ;
	7'h07 :
		TR_185 = TR_92 ;
	7'h08 :
		TR_185 = TR_92 ;
	7'h09 :
		TR_185 = TR_92 ;
	7'h0a :
		TR_185 = TR_92 ;
	7'h0b :
		TR_185 = TR_92 ;
	7'h0c :
		TR_185 = TR_92 ;
	7'h0d :
		TR_185 = TR_92 ;
	7'h0e :
		TR_185 = TR_92 ;
	7'h0f :
		TR_185 = TR_92 ;
	7'h10 :
		TR_185 = TR_92 ;
	7'h11 :
		TR_185 = TR_92 ;
	7'h12 :
		TR_185 = TR_92 ;
	7'h13 :
		TR_185 = TR_92 ;
	7'h14 :
		TR_185 = TR_92 ;
	7'h15 :
		TR_185 = TR_92 ;
	7'h16 :
		TR_185 = TR_92 ;
	7'h17 :
		TR_185 = TR_92 ;
	7'h18 :
		TR_185 = TR_92 ;
	7'h19 :
		TR_185 = TR_92 ;
	7'h1a :
		TR_185 = TR_92 ;
	7'h1b :
		TR_185 = TR_92 ;
	7'h1c :
		TR_185 = TR_92 ;
	7'h1d :
		TR_185 = TR_92 ;
	7'h1e :
		TR_185 = TR_92 ;
	7'h1f :
		TR_185 = TR_92 ;
	7'h20 :
		TR_185 = TR_92 ;
	7'h21 :
		TR_185 = TR_92 ;
	7'h22 :
		TR_185 = TR_92 ;
	7'h23 :
		TR_185 = TR_92 ;
	7'h24 :
		TR_185 = TR_92 ;
	7'h25 :
		TR_185 = TR_92 ;
	7'h26 :
		TR_185 = TR_92 ;
	7'h27 :
		TR_185 = TR_92 ;
	7'h28 :
		TR_185 = TR_92 ;
	7'h29 :
		TR_185 = TR_92 ;
	7'h2a :
		TR_185 = TR_92 ;
	7'h2b :
		TR_185 = TR_92 ;
	7'h2c :
		TR_185 = TR_92 ;
	7'h2d :
		TR_185 = TR_92 ;
	7'h2e :
		TR_185 = TR_92 ;
	7'h2f :
		TR_185 = TR_92 ;
	7'h30 :
		TR_185 = TR_92 ;
	7'h31 :
		TR_185 = TR_92 ;
	7'h32 :
		TR_185 = TR_92 ;
	7'h33 :
		TR_185 = TR_92 ;
	7'h34 :
		TR_185 = TR_92 ;
	7'h35 :
		TR_185 = TR_92 ;
	7'h36 :
		TR_185 = TR_92 ;
	7'h37 :
		TR_185 = TR_92 ;
	7'h38 :
		TR_185 = TR_92 ;
	7'h39 :
		TR_185 = TR_92 ;
	7'h3a :
		TR_185 = TR_92 ;
	7'h3b :
		TR_185 = TR_92 ;
	7'h3c :
		TR_185 = TR_92 ;
	7'h3d :
		TR_185 = TR_92 ;
	7'h3e :
		TR_185 = TR_92 ;
	7'h3f :
		TR_185 = TR_92 ;
	7'h40 :
		TR_185 = TR_92 ;
	7'h41 :
		TR_185 = TR_92 ;
	7'h42 :
		TR_185 = TR_92 ;
	7'h43 :
		TR_185 = TR_92 ;
	7'h44 :
		TR_185 = TR_92 ;
	7'h45 :
		TR_185 = TR_92 ;
	7'h46 :
		TR_185 = TR_92 ;
	7'h47 :
		TR_185 = TR_92 ;
	7'h48 :
		TR_185 = TR_92 ;
	7'h49 :
		TR_185 = TR_92 ;
	7'h4a :
		TR_185 = TR_92 ;
	7'h4b :
		TR_185 = TR_92 ;
	7'h4c :
		TR_185 = TR_92 ;
	7'h4d :
		TR_185 = TR_92 ;
	7'h4e :
		TR_185 = TR_92 ;
	7'h4f :
		TR_185 = TR_92 ;
	7'h50 :
		TR_185 = 9'h000 ;	// line#=../rle.cpp:80
	7'h51 :
		TR_185 = TR_92 ;
	7'h52 :
		TR_185 = TR_92 ;
	7'h53 :
		TR_185 = TR_92 ;
	7'h54 :
		TR_185 = TR_92 ;
	7'h55 :
		TR_185 = TR_92 ;
	7'h56 :
		TR_185 = TR_92 ;
	7'h57 :
		TR_185 = TR_92 ;
	7'h58 :
		TR_185 = TR_92 ;
	7'h59 :
		TR_185 = TR_92 ;
	7'h5a :
		TR_185 = TR_92 ;
	7'h5b :
		TR_185 = TR_92 ;
	7'h5c :
		TR_185 = TR_92 ;
	7'h5d :
		TR_185 = TR_92 ;
	7'h5e :
		TR_185 = TR_92 ;
	7'h5f :
		TR_185 = TR_92 ;
	7'h60 :
		TR_185 = TR_92 ;
	7'h61 :
		TR_185 = TR_92 ;
	7'h62 :
		TR_185 = TR_92 ;
	7'h63 :
		TR_185 = TR_92 ;
	7'h64 :
		TR_185 = TR_92 ;
	7'h65 :
		TR_185 = TR_92 ;
	7'h66 :
		TR_185 = TR_92 ;
	7'h67 :
		TR_185 = TR_92 ;
	7'h68 :
		TR_185 = TR_92 ;
	7'h69 :
		TR_185 = TR_92 ;
	7'h6a :
		TR_185 = TR_92 ;
	7'h6b :
		TR_185 = TR_92 ;
	7'h6c :
		TR_185 = TR_92 ;
	7'h6d :
		TR_185 = TR_92 ;
	7'h6e :
		TR_185 = TR_92 ;
	7'h6f :
		TR_185 = TR_92 ;
	7'h70 :
		TR_185 = TR_92 ;
	7'h71 :
		TR_185 = TR_92 ;
	7'h72 :
		TR_185 = TR_92 ;
	7'h73 :
		TR_185 = TR_92 ;
	7'h74 :
		TR_185 = TR_92 ;
	7'h75 :
		TR_185 = TR_92 ;
	7'h76 :
		TR_185 = TR_92 ;
	7'h77 :
		TR_185 = TR_92 ;
	7'h78 :
		TR_185 = TR_92 ;
	7'h79 :
		TR_185 = TR_92 ;
	7'h7a :
		TR_185 = TR_92 ;
	7'h7b :
		TR_185 = TR_92 ;
	7'h7c :
		TR_185 = TR_92 ;
	7'h7d :
		TR_185 = TR_92 ;
	7'h7e :
		TR_185 = TR_92 ;
	7'h7f :
		TR_185 = TR_92 ;
	default :
		TR_185 = 9'hx ;
	endcase
always @ ( TR_185 or U_173 or sub8u_71ot or U_183 or RG_rl_169 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_80_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h50 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_80_t = ( ( { 9{ M_180 } } & RG_rl_169 )
		| ( { 9{ U_173 } } & TR_185 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_80_en = ( M_180 | RG_rl_80_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_80_en )
		RG_rl_80 <= RG_rl_80_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_93 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_184 = TR_93 ;
	7'h01 :
		TR_184 = TR_93 ;
	7'h02 :
		TR_184 = TR_93 ;
	7'h03 :
		TR_184 = TR_93 ;
	7'h04 :
		TR_184 = TR_93 ;
	7'h05 :
		TR_184 = TR_93 ;
	7'h06 :
		TR_184 = TR_93 ;
	7'h07 :
		TR_184 = TR_93 ;
	7'h08 :
		TR_184 = TR_93 ;
	7'h09 :
		TR_184 = TR_93 ;
	7'h0a :
		TR_184 = TR_93 ;
	7'h0b :
		TR_184 = TR_93 ;
	7'h0c :
		TR_184 = TR_93 ;
	7'h0d :
		TR_184 = TR_93 ;
	7'h0e :
		TR_184 = TR_93 ;
	7'h0f :
		TR_184 = TR_93 ;
	7'h10 :
		TR_184 = TR_93 ;
	7'h11 :
		TR_184 = TR_93 ;
	7'h12 :
		TR_184 = TR_93 ;
	7'h13 :
		TR_184 = TR_93 ;
	7'h14 :
		TR_184 = TR_93 ;
	7'h15 :
		TR_184 = TR_93 ;
	7'h16 :
		TR_184 = TR_93 ;
	7'h17 :
		TR_184 = TR_93 ;
	7'h18 :
		TR_184 = TR_93 ;
	7'h19 :
		TR_184 = TR_93 ;
	7'h1a :
		TR_184 = TR_93 ;
	7'h1b :
		TR_184 = TR_93 ;
	7'h1c :
		TR_184 = TR_93 ;
	7'h1d :
		TR_184 = TR_93 ;
	7'h1e :
		TR_184 = TR_93 ;
	7'h1f :
		TR_184 = TR_93 ;
	7'h20 :
		TR_184 = TR_93 ;
	7'h21 :
		TR_184 = TR_93 ;
	7'h22 :
		TR_184 = TR_93 ;
	7'h23 :
		TR_184 = TR_93 ;
	7'h24 :
		TR_184 = TR_93 ;
	7'h25 :
		TR_184 = TR_93 ;
	7'h26 :
		TR_184 = TR_93 ;
	7'h27 :
		TR_184 = TR_93 ;
	7'h28 :
		TR_184 = TR_93 ;
	7'h29 :
		TR_184 = TR_93 ;
	7'h2a :
		TR_184 = TR_93 ;
	7'h2b :
		TR_184 = TR_93 ;
	7'h2c :
		TR_184 = TR_93 ;
	7'h2d :
		TR_184 = TR_93 ;
	7'h2e :
		TR_184 = TR_93 ;
	7'h2f :
		TR_184 = TR_93 ;
	7'h30 :
		TR_184 = TR_93 ;
	7'h31 :
		TR_184 = TR_93 ;
	7'h32 :
		TR_184 = TR_93 ;
	7'h33 :
		TR_184 = TR_93 ;
	7'h34 :
		TR_184 = TR_93 ;
	7'h35 :
		TR_184 = TR_93 ;
	7'h36 :
		TR_184 = TR_93 ;
	7'h37 :
		TR_184 = TR_93 ;
	7'h38 :
		TR_184 = TR_93 ;
	7'h39 :
		TR_184 = TR_93 ;
	7'h3a :
		TR_184 = TR_93 ;
	7'h3b :
		TR_184 = TR_93 ;
	7'h3c :
		TR_184 = TR_93 ;
	7'h3d :
		TR_184 = TR_93 ;
	7'h3e :
		TR_184 = TR_93 ;
	7'h3f :
		TR_184 = TR_93 ;
	7'h40 :
		TR_184 = TR_93 ;
	7'h41 :
		TR_184 = TR_93 ;
	7'h42 :
		TR_184 = TR_93 ;
	7'h43 :
		TR_184 = TR_93 ;
	7'h44 :
		TR_184 = TR_93 ;
	7'h45 :
		TR_184 = TR_93 ;
	7'h46 :
		TR_184 = TR_93 ;
	7'h47 :
		TR_184 = TR_93 ;
	7'h48 :
		TR_184 = TR_93 ;
	7'h49 :
		TR_184 = TR_93 ;
	7'h4a :
		TR_184 = TR_93 ;
	7'h4b :
		TR_184 = TR_93 ;
	7'h4c :
		TR_184 = TR_93 ;
	7'h4d :
		TR_184 = TR_93 ;
	7'h4e :
		TR_184 = TR_93 ;
	7'h4f :
		TR_184 = TR_93 ;
	7'h50 :
		TR_184 = TR_93 ;
	7'h51 :
		TR_184 = 9'h000 ;	// line#=../rle.cpp:80
	7'h52 :
		TR_184 = TR_93 ;
	7'h53 :
		TR_184 = TR_93 ;
	7'h54 :
		TR_184 = TR_93 ;
	7'h55 :
		TR_184 = TR_93 ;
	7'h56 :
		TR_184 = TR_93 ;
	7'h57 :
		TR_184 = TR_93 ;
	7'h58 :
		TR_184 = TR_93 ;
	7'h59 :
		TR_184 = TR_93 ;
	7'h5a :
		TR_184 = TR_93 ;
	7'h5b :
		TR_184 = TR_93 ;
	7'h5c :
		TR_184 = TR_93 ;
	7'h5d :
		TR_184 = TR_93 ;
	7'h5e :
		TR_184 = TR_93 ;
	7'h5f :
		TR_184 = TR_93 ;
	7'h60 :
		TR_184 = TR_93 ;
	7'h61 :
		TR_184 = TR_93 ;
	7'h62 :
		TR_184 = TR_93 ;
	7'h63 :
		TR_184 = TR_93 ;
	7'h64 :
		TR_184 = TR_93 ;
	7'h65 :
		TR_184 = TR_93 ;
	7'h66 :
		TR_184 = TR_93 ;
	7'h67 :
		TR_184 = TR_93 ;
	7'h68 :
		TR_184 = TR_93 ;
	7'h69 :
		TR_184 = TR_93 ;
	7'h6a :
		TR_184 = TR_93 ;
	7'h6b :
		TR_184 = TR_93 ;
	7'h6c :
		TR_184 = TR_93 ;
	7'h6d :
		TR_184 = TR_93 ;
	7'h6e :
		TR_184 = TR_93 ;
	7'h6f :
		TR_184 = TR_93 ;
	7'h70 :
		TR_184 = TR_93 ;
	7'h71 :
		TR_184 = TR_93 ;
	7'h72 :
		TR_184 = TR_93 ;
	7'h73 :
		TR_184 = TR_93 ;
	7'h74 :
		TR_184 = TR_93 ;
	7'h75 :
		TR_184 = TR_93 ;
	7'h76 :
		TR_184 = TR_93 ;
	7'h77 :
		TR_184 = TR_93 ;
	7'h78 :
		TR_184 = TR_93 ;
	7'h79 :
		TR_184 = TR_93 ;
	7'h7a :
		TR_184 = TR_93 ;
	7'h7b :
		TR_184 = TR_93 ;
	7'h7c :
		TR_184 = TR_93 ;
	7'h7d :
		TR_184 = TR_93 ;
	7'h7e :
		TR_184 = TR_93 ;
	7'h7f :
		TR_184 = TR_93 ;
	default :
		TR_184 = 9'hx ;
	endcase
always @ ( TR_184 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_38 or 
	U_174 or RG_rl_169 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_81_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h51 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_81_t = ( ( { 9{ ST1_03d } } & RG_rl_169 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_38 )
		| ( { 9{ U_173 } } & TR_184 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_81_en = ( ST1_03d | U_174 | RG_rl_81_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_81_en )
		RG_rl_81 <= RG_rl_81_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_94 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_183 = TR_94 ;
	7'h01 :
		TR_183 = TR_94 ;
	7'h02 :
		TR_183 = TR_94 ;
	7'h03 :
		TR_183 = TR_94 ;
	7'h04 :
		TR_183 = TR_94 ;
	7'h05 :
		TR_183 = TR_94 ;
	7'h06 :
		TR_183 = TR_94 ;
	7'h07 :
		TR_183 = TR_94 ;
	7'h08 :
		TR_183 = TR_94 ;
	7'h09 :
		TR_183 = TR_94 ;
	7'h0a :
		TR_183 = TR_94 ;
	7'h0b :
		TR_183 = TR_94 ;
	7'h0c :
		TR_183 = TR_94 ;
	7'h0d :
		TR_183 = TR_94 ;
	7'h0e :
		TR_183 = TR_94 ;
	7'h0f :
		TR_183 = TR_94 ;
	7'h10 :
		TR_183 = TR_94 ;
	7'h11 :
		TR_183 = TR_94 ;
	7'h12 :
		TR_183 = TR_94 ;
	7'h13 :
		TR_183 = TR_94 ;
	7'h14 :
		TR_183 = TR_94 ;
	7'h15 :
		TR_183 = TR_94 ;
	7'h16 :
		TR_183 = TR_94 ;
	7'h17 :
		TR_183 = TR_94 ;
	7'h18 :
		TR_183 = TR_94 ;
	7'h19 :
		TR_183 = TR_94 ;
	7'h1a :
		TR_183 = TR_94 ;
	7'h1b :
		TR_183 = TR_94 ;
	7'h1c :
		TR_183 = TR_94 ;
	7'h1d :
		TR_183 = TR_94 ;
	7'h1e :
		TR_183 = TR_94 ;
	7'h1f :
		TR_183 = TR_94 ;
	7'h20 :
		TR_183 = TR_94 ;
	7'h21 :
		TR_183 = TR_94 ;
	7'h22 :
		TR_183 = TR_94 ;
	7'h23 :
		TR_183 = TR_94 ;
	7'h24 :
		TR_183 = TR_94 ;
	7'h25 :
		TR_183 = TR_94 ;
	7'h26 :
		TR_183 = TR_94 ;
	7'h27 :
		TR_183 = TR_94 ;
	7'h28 :
		TR_183 = TR_94 ;
	7'h29 :
		TR_183 = TR_94 ;
	7'h2a :
		TR_183 = TR_94 ;
	7'h2b :
		TR_183 = TR_94 ;
	7'h2c :
		TR_183 = TR_94 ;
	7'h2d :
		TR_183 = TR_94 ;
	7'h2e :
		TR_183 = TR_94 ;
	7'h2f :
		TR_183 = TR_94 ;
	7'h30 :
		TR_183 = TR_94 ;
	7'h31 :
		TR_183 = TR_94 ;
	7'h32 :
		TR_183 = TR_94 ;
	7'h33 :
		TR_183 = TR_94 ;
	7'h34 :
		TR_183 = TR_94 ;
	7'h35 :
		TR_183 = TR_94 ;
	7'h36 :
		TR_183 = TR_94 ;
	7'h37 :
		TR_183 = TR_94 ;
	7'h38 :
		TR_183 = TR_94 ;
	7'h39 :
		TR_183 = TR_94 ;
	7'h3a :
		TR_183 = TR_94 ;
	7'h3b :
		TR_183 = TR_94 ;
	7'h3c :
		TR_183 = TR_94 ;
	7'h3d :
		TR_183 = TR_94 ;
	7'h3e :
		TR_183 = TR_94 ;
	7'h3f :
		TR_183 = TR_94 ;
	7'h40 :
		TR_183 = TR_94 ;
	7'h41 :
		TR_183 = TR_94 ;
	7'h42 :
		TR_183 = TR_94 ;
	7'h43 :
		TR_183 = TR_94 ;
	7'h44 :
		TR_183 = TR_94 ;
	7'h45 :
		TR_183 = TR_94 ;
	7'h46 :
		TR_183 = TR_94 ;
	7'h47 :
		TR_183 = TR_94 ;
	7'h48 :
		TR_183 = TR_94 ;
	7'h49 :
		TR_183 = TR_94 ;
	7'h4a :
		TR_183 = TR_94 ;
	7'h4b :
		TR_183 = TR_94 ;
	7'h4c :
		TR_183 = TR_94 ;
	7'h4d :
		TR_183 = TR_94 ;
	7'h4e :
		TR_183 = TR_94 ;
	7'h4f :
		TR_183 = TR_94 ;
	7'h50 :
		TR_183 = TR_94 ;
	7'h51 :
		TR_183 = TR_94 ;
	7'h52 :
		TR_183 = 9'h000 ;	// line#=../rle.cpp:80
	7'h53 :
		TR_183 = TR_94 ;
	7'h54 :
		TR_183 = TR_94 ;
	7'h55 :
		TR_183 = TR_94 ;
	7'h56 :
		TR_183 = TR_94 ;
	7'h57 :
		TR_183 = TR_94 ;
	7'h58 :
		TR_183 = TR_94 ;
	7'h59 :
		TR_183 = TR_94 ;
	7'h5a :
		TR_183 = TR_94 ;
	7'h5b :
		TR_183 = TR_94 ;
	7'h5c :
		TR_183 = TR_94 ;
	7'h5d :
		TR_183 = TR_94 ;
	7'h5e :
		TR_183 = TR_94 ;
	7'h5f :
		TR_183 = TR_94 ;
	7'h60 :
		TR_183 = TR_94 ;
	7'h61 :
		TR_183 = TR_94 ;
	7'h62 :
		TR_183 = TR_94 ;
	7'h63 :
		TR_183 = TR_94 ;
	7'h64 :
		TR_183 = TR_94 ;
	7'h65 :
		TR_183 = TR_94 ;
	7'h66 :
		TR_183 = TR_94 ;
	7'h67 :
		TR_183 = TR_94 ;
	7'h68 :
		TR_183 = TR_94 ;
	7'h69 :
		TR_183 = TR_94 ;
	7'h6a :
		TR_183 = TR_94 ;
	7'h6b :
		TR_183 = TR_94 ;
	7'h6c :
		TR_183 = TR_94 ;
	7'h6d :
		TR_183 = TR_94 ;
	7'h6e :
		TR_183 = TR_94 ;
	7'h6f :
		TR_183 = TR_94 ;
	7'h70 :
		TR_183 = TR_94 ;
	7'h71 :
		TR_183 = TR_94 ;
	7'h72 :
		TR_183 = TR_94 ;
	7'h73 :
		TR_183 = TR_94 ;
	7'h74 :
		TR_183 = TR_94 ;
	7'h75 :
		TR_183 = TR_94 ;
	7'h76 :
		TR_183 = TR_94 ;
	7'h77 :
		TR_183 = TR_94 ;
	7'h78 :
		TR_183 = TR_94 ;
	7'h79 :
		TR_183 = TR_94 ;
	7'h7a :
		TR_183 = TR_94 ;
	7'h7b :
		TR_183 = TR_94 ;
	7'h7c :
		TR_183 = TR_94 ;
	7'h7d :
		TR_183 = TR_94 ;
	7'h7e :
		TR_183 = TR_94 ;
	7'h7f :
		TR_183 = TR_94 ;
	default :
		TR_183 = 9'hx ;
	endcase
always @ ( TR_183 or U_173 or sub8u_71ot or U_183 or RG_rl_170 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_82_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h52 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_82_t = ( ( { 9{ M_180 } } & RG_rl_170 )
		| ( { 9{ U_173 } } & TR_183 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_82_en = ( M_180 | RG_rl_82_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_82_en )
		RG_rl_82 <= RG_rl_82_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_95 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_182 = TR_95 ;
	7'h01 :
		TR_182 = TR_95 ;
	7'h02 :
		TR_182 = TR_95 ;
	7'h03 :
		TR_182 = TR_95 ;
	7'h04 :
		TR_182 = TR_95 ;
	7'h05 :
		TR_182 = TR_95 ;
	7'h06 :
		TR_182 = TR_95 ;
	7'h07 :
		TR_182 = TR_95 ;
	7'h08 :
		TR_182 = TR_95 ;
	7'h09 :
		TR_182 = TR_95 ;
	7'h0a :
		TR_182 = TR_95 ;
	7'h0b :
		TR_182 = TR_95 ;
	7'h0c :
		TR_182 = TR_95 ;
	7'h0d :
		TR_182 = TR_95 ;
	7'h0e :
		TR_182 = TR_95 ;
	7'h0f :
		TR_182 = TR_95 ;
	7'h10 :
		TR_182 = TR_95 ;
	7'h11 :
		TR_182 = TR_95 ;
	7'h12 :
		TR_182 = TR_95 ;
	7'h13 :
		TR_182 = TR_95 ;
	7'h14 :
		TR_182 = TR_95 ;
	7'h15 :
		TR_182 = TR_95 ;
	7'h16 :
		TR_182 = TR_95 ;
	7'h17 :
		TR_182 = TR_95 ;
	7'h18 :
		TR_182 = TR_95 ;
	7'h19 :
		TR_182 = TR_95 ;
	7'h1a :
		TR_182 = TR_95 ;
	7'h1b :
		TR_182 = TR_95 ;
	7'h1c :
		TR_182 = TR_95 ;
	7'h1d :
		TR_182 = TR_95 ;
	7'h1e :
		TR_182 = TR_95 ;
	7'h1f :
		TR_182 = TR_95 ;
	7'h20 :
		TR_182 = TR_95 ;
	7'h21 :
		TR_182 = TR_95 ;
	7'h22 :
		TR_182 = TR_95 ;
	7'h23 :
		TR_182 = TR_95 ;
	7'h24 :
		TR_182 = TR_95 ;
	7'h25 :
		TR_182 = TR_95 ;
	7'h26 :
		TR_182 = TR_95 ;
	7'h27 :
		TR_182 = TR_95 ;
	7'h28 :
		TR_182 = TR_95 ;
	7'h29 :
		TR_182 = TR_95 ;
	7'h2a :
		TR_182 = TR_95 ;
	7'h2b :
		TR_182 = TR_95 ;
	7'h2c :
		TR_182 = TR_95 ;
	7'h2d :
		TR_182 = TR_95 ;
	7'h2e :
		TR_182 = TR_95 ;
	7'h2f :
		TR_182 = TR_95 ;
	7'h30 :
		TR_182 = TR_95 ;
	7'h31 :
		TR_182 = TR_95 ;
	7'h32 :
		TR_182 = TR_95 ;
	7'h33 :
		TR_182 = TR_95 ;
	7'h34 :
		TR_182 = TR_95 ;
	7'h35 :
		TR_182 = TR_95 ;
	7'h36 :
		TR_182 = TR_95 ;
	7'h37 :
		TR_182 = TR_95 ;
	7'h38 :
		TR_182 = TR_95 ;
	7'h39 :
		TR_182 = TR_95 ;
	7'h3a :
		TR_182 = TR_95 ;
	7'h3b :
		TR_182 = TR_95 ;
	7'h3c :
		TR_182 = TR_95 ;
	7'h3d :
		TR_182 = TR_95 ;
	7'h3e :
		TR_182 = TR_95 ;
	7'h3f :
		TR_182 = TR_95 ;
	7'h40 :
		TR_182 = TR_95 ;
	7'h41 :
		TR_182 = TR_95 ;
	7'h42 :
		TR_182 = TR_95 ;
	7'h43 :
		TR_182 = TR_95 ;
	7'h44 :
		TR_182 = TR_95 ;
	7'h45 :
		TR_182 = TR_95 ;
	7'h46 :
		TR_182 = TR_95 ;
	7'h47 :
		TR_182 = TR_95 ;
	7'h48 :
		TR_182 = TR_95 ;
	7'h49 :
		TR_182 = TR_95 ;
	7'h4a :
		TR_182 = TR_95 ;
	7'h4b :
		TR_182 = TR_95 ;
	7'h4c :
		TR_182 = TR_95 ;
	7'h4d :
		TR_182 = TR_95 ;
	7'h4e :
		TR_182 = TR_95 ;
	7'h4f :
		TR_182 = TR_95 ;
	7'h50 :
		TR_182 = TR_95 ;
	7'h51 :
		TR_182 = TR_95 ;
	7'h52 :
		TR_182 = TR_95 ;
	7'h53 :
		TR_182 = 9'h000 ;	// line#=../rle.cpp:80
	7'h54 :
		TR_182 = TR_95 ;
	7'h55 :
		TR_182 = TR_95 ;
	7'h56 :
		TR_182 = TR_95 ;
	7'h57 :
		TR_182 = TR_95 ;
	7'h58 :
		TR_182 = TR_95 ;
	7'h59 :
		TR_182 = TR_95 ;
	7'h5a :
		TR_182 = TR_95 ;
	7'h5b :
		TR_182 = TR_95 ;
	7'h5c :
		TR_182 = TR_95 ;
	7'h5d :
		TR_182 = TR_95 ;
	7'h5e :
		TR_182 = TR_95 ;
	7'h5f :
		TR_182 = TR_95 ;
	7'h60 :
		TR_182 = TR_95 ;
	7'h61 :
		TR_182 = TR_95 ;
	7'h62 :
		TR_182 = TR_95 ;
	7'h63 :
		TR_182 = TR_95 ;
	7'h64 :
		TR_182 = TR_95 ;
	7'h65 :
		TR_182 = TR_95 ;
	7'h66 :
		TR_182 = TR_95 ;
	7'h67 :
		TR_182 = TR_95 ;
	7'h68 :
		TR_182 = TR_95 ;
	7'h69 :
		TR_182 = TR_95 ;
	7'h6a :
		TR_182 = TR_95 ;
	7'h6b :
		TR_182 = TR_95 ;
	7'h6c :
		TR_182 = TR_95 ;
	7'h6d :
		TR_182 = TR_95 ;
	7'h6e :
		TR_182 = TR_95 ;
	7'h6f :
		TR_182 = TR_95 ;
	7'h70 :
		TR_182 = TR_95 ;
	7'h71 :
		TR_182 = TR_95 ;
	7'h72 :
		TR_182 = TR_95 ;
	7'h73 :
		TR_182 = TR_95 ;
	7'h74 :
		TR_182 = TR_95 ;
	7'h75 :
		TR_182 = TR_95 ;
	7'h76 :
		TR_182 = TR_95 ;
	7'h77 :
		TR_182 = TR_95 ;
	7'h78 :
		TR_182 = TR_95 ;
	7'h79 :
		TR_182 = TR_95 ;
	7'h7a :
		TR_182 = TR_95 ;
	7'h7b :
		TR_182 = TR_95 ;
	7'h7c :
		TR_182 = TR_95 ;
	7'h7d :
		TR_182 = TR_95 ;
	7'h7e :
		TR_182 = TR_95 ;
	7'h7f :
		TR_182 = TR_95 ;
	default :
		TR_182 = 9'hx ;
	endcase
always @ ( TR_182 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_39 or 
	U_174 or RG_rl_170 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_83_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h53 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_83_t = ( ( { 9{ ST1_03d } } & RG_rl_170 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_39 )
		| ( { 9{ U_173 } } & TR_182 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_83_en = ( ST1_03d | U_174 | RG_rl_83_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_83_en )
		RG_rl_83 <= RG_rl_83_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_96 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_181 = TR_96 ;
	7'h01 :
		TR_181 = TR_96 ;
	7'h02 :
		TR_181 = TR_96 ;
	7'h03 :
		TR_181 = TR_96 ;
	7'h04 :
		TR_181 = TR_96 ;
	7'h05 :
		TR_181 = TR_96 ;
	7'h06 :
		TR_181 = TR_96 ;
	7'h07 :
		TR_181 = TR_96 ;
	7'h08 :
		TR_181 = TR_96 ;
	7'h09 :
		TR_181 = TR_96 ;
	7'h0a :
		TR_181 = TR_96 ;
	7'h0b :
		TR_181 = TR_96 ;
	7'h0c :
		TR_181 = TR_96 ;
	7'h0d :
		TR_181 = TR_96 ;
	7'h0e :
		TR_181 = TR_96 ;
	7'h0f :
		TR_181 = TR_96 ;
	7'h10 :
		TR_181 = TR_96 ;
	7'h11 :
		TR_181 = TR_96 ;
	7'h12 :
		TR_181 = TR_96 ;
	7'h13 :
		TR_181 = TR_96 ;
	7'h14 :
		TR_181 = TR_96 ;
	7'h15 :
		TR_181 = TR_96 ;
	7'h16 :
		TR_181 = TR_96 ;
	7'h17 :
		TR_181 = TR_96 ;
	7'h18 :
		TR_181 = TR_96 ;
	7'h19 :
		TR_181 = TR_96 ;
	7'h1a :
		TR_181 = TR_96 ;
	7'h1b :
		TR_181 = TR_96 ;
	7'h1c :
		TR_181 = TR_96 ;
	7'h1d :
		TR_181 = TR_96 ;
	7'h1e :
		TR_181 = TR_96 ;
	7'h1f :
		TR_181 = TR_96 ;
	7'h20 :
		TR_181 = TR_96 ;
	7'h21 :
		TR_181 = TR_96 ;
	7'h22 :
		TR_181 = TR_96 ;
	7'h23 :
		TR_181 = TR_96 ;
	7'h24 :
		TR_181 = TR_96 ;
	7'h25 :
		TR_181 = TR_96 ;
	7'h26 :
		TR_181 = TR_96 ;
	7'h27 :
		TR_181 = TR_96 ;
	7'h28 :
		TR_181 = TR_96 ;
	7'h29 :
		TR_181 = TR_96 ;
	7'h2a :
		TR_181 = TR_96 ;
	7'h2b :
		TR_181 = TR_96 ;
	7'h2c :
		TR_181 = TR_96 ;
	7'h2d :
		TR_181 = TR_96 ;
	7'h2e :
		TR_181 = TR_96 ;
	7'h2f :
		TR_181 = TR_96 ;
	7'h30 :
		TR_181 = TR_96 ;
	7'h31 :
		TR_181 = TR_96 ;
	7'h32 :
		TR_181 = TR_96 ;
	7'h33 :
		TR_181 = TR_96 ;
	7'h34 :
		TR_181 = TR_96 ;
	7'h35 :
		TR_181 = TR_96 ;
	7'h36 :
		TR_181 = TR_96 ;
	7'h37 :
		TR_181 = TR_96 ;
	7'h38 :
		TR_181 = TR_96 ;
	7'h39 :
		TR_181 = TR_96 ;
	7'h3a :
		TR_181 = TR_96 ;
	7'h3b :
		TR_181 = TR_96 ;
	7'h3c :
		TR_181 = TR_96 ;
	7'h3d :
		TR_181 = TR_96 ;
	7'h3e :
		TR_181 = TR_96 ;
	7'h3f :
		TR_181 = TR_96 ;
	7'h40 :
		TR_181 = TR_96 ;
	7'h41 :
		TR_181 = TR_96 ;
	7'h42 :
		TR_181 = TR_96 ;
	7'h43 :
		TR_181 = TR_96 ;
	7'h44 :
		TR_181 = TR_96 ;
	7'h45 :
		TR_181 = TR_96 ;
	7'h46 :
		TR_181 = TR_96 ;
	7'h47 :
		TR_181 = TR_96 ;
	7'h48 :
		TR_181 = TR_96 ;
	7'h49 :
		TR_181 = TR_96 ;
	7'h4a :
		TR_181 = TR_96 ;
	7'h4b :
		TR_181 = TR_96 ;
	7'h4c :
		TR_181 = TR_96 ;
	7'h4d :
		TR_181 = TR_96 ;
	7'h4e :
		TR_181 = TR_96 ;
	7'h4f :
		TR_181 = TR_96 ;
	7'h50 :
		TR_181 = TR_96 ;
	7'h51 :
		TR_181 = TR_96 ;
	7'h52 :
		TR_181 = TR_96 ;
	7'h53 :
		TR_181 = TR_96 ;
	7'h54 :
		TR_181 = 9'h000 ;	// line#=../rle.cpp:80
	7'h55 :
		TR_181 = TR_96 ;
	7'h56 :
		TR_181 = TR_96 ;
	7'h57 :
		TR_181 = TR_96 ;
	7'h58 :
		TR_181 = TR_96 ;
	7'h59 :
		TR_181 = TR_96 ;
	7'h5a :
		TR_181 = TR_96 ;
	7'h5b :
		TR_181 = TR_96 ;
	7'h5c :
		TR_181 = TR_96 ;
	7'h5d :
		TR_181 = TR_96 ;
	7'h5e :
		TR_181 = TR_96 ;
	7'h5f :
		TR_181 = TR_96 ;
	7'h60 :
		TR_181 = TR_96 ;
	7'h61 :
		TR_181 = TR_96 ;
	7'h62 :
		TR_181 = TR_96 ;
	7'h63 :
		TR_181 = TR_96 ;
	7'h64 :
		TR_181 = TR_96 ;
	7'h65 :
		TR_181 = TR_96 ;
	7'h66 :
		TR_181 = TR_96 ;
	7'h67 :
		TR_181 = TR_96 ;
	7'h68 :
		TR_181 = TR_96 ;
	7'h69 :
		TR_181 = TR_96 ;
	7'h6a :
		TR_181 = TR_96 ;
	7'h6b :
		TR_181 = TR_96 ;
	7'h6c :
		TR_181 = TR_96 ;
	7'h6d :
		TR_181 = TR_96 ;
	7'h6e :
		TR_181 = TR_96 ;
	7'h6f :
		TR_181 = TR_96 ;
	7'h70 :
		TR_181 = TR_96 ;
	7'h71 :
		TR_181 = TR_96 ;
	7'h72 :
		TR_181 = TR_96 ;
	7'h73 :
		TR_181 = TR_96 ;
	7'h74 :
		TR_181 = TR_96 ;
	7'h75 :
		TR_181 = TR_96 ;
	7'h76 :
		TR_181 = TR_96 ;
	7'h77 :
		TR_181 = TR_96 ;
	7'h78 :
		TR_181 = TR_96 ;
	7'h79 :
		TR_181 = TR_96 ;
	7'h7a :
		TR_181 = TR_96 ;
	7'h7b :
		TR_181 = TR_96 ;
	7'h7c :
		TR_181 = TR_96 ;
	7'h7d :
		TR_181 = TR_96 ;
	7'h7e :
		TR_181 = TR_96 ;
	7'h7f :
		TR_181 = TR_96 ;
	default :
		TR_181 = 9'hx ;
	endcase
always @ ( TR_181 or U_173 or sub8u_71ot or U_183 or RG_rl_171 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_84_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h54 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_84_t = ( ( { 9{ M_180 } } & RG_rl_171 )
		| ( { 9{ U_173 } } & TR_181 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_84_en = ( M_180 | RG_rl_84_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_84_en )
		RG_rl_84 <= RG_rl_84_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_97 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_180 = TR_97 ;
	7'h01 :
		TR_180 = TR_97 ;
	7'h02 :
		TR_180 = TR_97 ;
	7'h03 :
		TR_180 = TR_97 ;
	7'h04 :
		TR_180 = TR_97 ;
	7'h05 :
		TR_180 = TR_97 ;
	7'h06 :
		TR_180 = TR_97 ;
	7'h07 :
		TR_180 = TR_97 ;
	7'h08 :
		TR_180 = TR_97 ;
	7'h09 :
		TR_180 = TR_97 ;
	7'h0a :
		TR_180 = TR_97 ;
	7'h0b :
		TR_180 = TR_97 ;
	7'h0c :
		TR_180 = TR_97 ;
	7'h0d :
		TR_180 = TR_97 ;
	7'h0e :
		TR_180 = TR_97 ;
	7'h0f :
		TR_180 = TR_97 ;
	7'h10 :
		TR_180 = TR_97 ;
	7'h11 :
		TR_180 = TR_97 ;
	7'h12 :
		TR_180 = TR_97 ;
	7'h13 :
		TR_180 = TR_97 ;
	7'h14 :
		TR_180 = TR_97 ;
	7'h15 :
		TR_180 = TR_97 ;
	7'h16 :
		TR_180 = TR_97 ;
	7'h17 :
		TR_180 = TR_97 ;
	7'h18 :
		TR_180 = TR_97 ;
	7'h19 :
		TR_180 = TR_97 ;
	7'h1a :
		TR_180 = TR_97 ;
	7'h1b :
		TR_180 = TR_97 ;
	7'h1c :
		TR_180 = TR_97 ;
	7'h1d :
		TR_180 = TR_97 ;
	7'h1e :
		TR_180 = TR_97 ;
	7'h1f :
		TR_180 = TR_97 ;
	7'h20 :
		TR_180 = TR_97 ;
	7'h21 :
		TR_180 = TR_97 ;
	7'h22 :
		TR_180 = TR_97 ;
	7'h23 :
		TR_180 = TR_97 ;
	7'h24 :
		TR_180 = TR_97 ;
	7'h25 :
		TR_180 = TR_97 ;
	7'h26 :
		TR_180 = TR_97 ;
	7'h27 :
		TR_180 = TR_97 ;
	7'h28 :
		TR_180 = TR_97 ;
	7'h29 :
		TR_180 = TR_97 ;
	7'h2a :
		TR_180 = TR_97 ;
	7'h2b :
		TR_180 = TR_97 ;
	7'h2c :
		TR_180 = TR_97 ;
	7'h2d :
		TR_180 = TR_97 ;
	7'h2e :
		TR_180 = TR_97 ;
	7'h2f :
		TR_180 = TR_97 ;
	7'h30 :
		TR_180 = TR_97 ;
	7'h31 :
		TR_180 = TR_97 ;
	7'h32 :
		TR_180 = TR_97 ;
	7'h33 :
		TR_180 = TR_97 ;
	7'h34 :
		TR_180 = TR_97 ;
	7'h35 :
		TR_180 = TR_97 ;
	7'h36 :
		TR_180 = TR_97 ;
	7'h37 :
		TR_180 = TR_97 ;
	7'h38 :
		TR_180 = TR_97 ;
	7'h39 :
		TR_180 = TR_97 ;
	7'h3a :
		TR_180 = TR_97 ;
	7'h3b :
		TR_180 = TR_97 ;
	7'h3c :
		TR_180 = TR_97 ;
	7'h3d :
		TR_180 = TR_97 ;
	7'h3e :
		TR_180 = TR_97 ;
	7'h3f :
		TR_180 = TR_97 ;
	7'h40 :
		TR_180 = TR_97 ;
	7'h41 :
		TR_180 = TR_97 ;
	7'h42 :
		TR_180 = TR_97 ;
	7'h43 :
		TR_180 = TR_97 ;
	7'h44 :
		TR_180 = TR_97 ;
	7'h45 :
		TR_180 = TR_97 ;
	7'h46 :
		TR_180 = TR_97 ;
	7'h47 :
		TR_180 = TR_97 ;
	7'h48 :
		TR_180 = TR_97 ;
	7'h49 :
		TR_180 = TR_97 ;
	7'h4a :
		TR_180 = TR_97 ;
	7'h4b :
		TR_180 = TR_97 ;
	7'h4c :
		TR_180 = TR_97 ;
	7'h4d :
		TR_180 = TR_97 ;
	7'h4e :
		TR_180 = TR_97 ;
	7'h4f :
		TR_180 = TR_97 ;
	7'h50 :
		TR_180 = TR_97 ;
	7'h51 :
		TR_180 = TR_97 ;
	7'h52 :
		TR_180 = TR_97 ;
	7'h53 :
		TR_180 = TR_97 ;
	7'h54 :
		TR_180 = TR_97 ;
	7'h55 :
		TR_180 = 9'h000 ;	// line#=../rle.cpp:80
	7'h56 :
		TR_180 = TR_97 ;
	7'h57 :
		TR_180 = TR_97 ;
	7'h58 :
		TR_180 = TR_97 ;
	7'h59 :
		TR_180 = TR_97 ;
	7'h5a :
		TR_180 = TR_97 ;
	7'h5b :
		TR_180 = TR_97 ;
	7'h5c :
		TR_180 = TR_97 ;
	7'h5d :
		TR_180 = TR_97 ;
	7'h5e :
		TR_180 = TR_97 ;
	7'h5f :
		TR_180 = TR_97 ;
	7'h60 :
		TR_180 = TR_97 ;
	7'h61 :
		TR_180 = TR_97 ;
	7'h62 :
		TR_180 = TR_97 ;
	7'h63 :
		TR_180 = TR_97 ;
	7'h64 :
		TR_180 = TR_97 ;
	7'h65 :
		TR_180 = TR_97 ;
	7'h66 :
		TR_180 = TR_97 ;
	7'h67 :
		TR_180 = TR_97 ;
	7'h68 :
		TR_180 = TR_97 ;
	7'h69 :
		TR_180 = TR_97 ;
	7'h6a :
		TR_180 = TR_97 ;
	7'h6b :
		TR_180 = TR_97 ;
	7'h6c :
		TR_180 = TR_97 ;
	7'h6d :
		TR_180 = TR_97 ;
	7'h6e :
		TR_180 = TR_97 ;
	7'h6f :
		TR_180 = TR_97 ;
	7'h70 :
		TR_180 = TR_97 ;
	7'h71 :
		TR_180 = TR_97 ;
	7'h72 :
		TR_180 = TR_97 ;
	7'h73 :
		TR_180 = TR_97 ;
	7'h74 :
		TR_180 = TR_97 ;
	7'h75 :
		TR_180 = TR_97 ;
	7'h76 :
		TR_180 = TR_97 ;
	7'h77 :
		TR_180 = TR_97 ;
	7'h78 :
		TR_180 = TR_97 ;
	7'h79 :
		TR_180 = TR_97 ;
	7'h7a :
		TR_180 = TR_97 ;
	7'h7b :
		TR_180 = TR_97 ;
	7'h7c :
		TR_180 = TR_97 ;
	7'h7d :
		TR_180 = TR_97 ;
	7'h7e :
		TR_180 = TR_97 ;
	7'h7f :
		TR_180 = TR_97 ;
	default :
		TR_180 = 9'hx ;
	endcase
always @ ( TR_180 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_40 or 
	U_174 or RG_rl_171 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_85_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h55 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_85_t = ( ( { 9{ ST1_03d } } & RG_rl_171 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_40 )
		| ( { 9{ U_173 } } & TR_180 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_85_en = ( ST1_03d | U_174 | RG_rl_85_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_85_en )
		RG_rl_85 <= RG_rl_85_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_98 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_179 = TR_98 ;
	7'h01 :
		TR_179 = TR_98 ;
	7'h02 :
		TR_179 = TR_98 ;
	7'h03 :
		TR_179 = TR_98 ;
	7'h04 :
		TR_179 = TR_98 ;
	7'h05 :
		TR_179 = TR_98 ;
	7'h06 :
		TR_179 = TR_98 ;
	7'h07 :
		TR_179 = TR_98 ;
	7'h08 :
		TR_179 = TR_98 ;
	7'h09 :
		TR_179 = TR_98 ;
	7'h0a :
		TR_179 = TR_98 ;
	7'h0b :
		TR_179 = TR_98 ;
	7'h0c :
		TR_179 = TR_98 ;
	7'h0d :
		TR_179 = TR_98 ;
	7'h0e :
		TR_179 = TR_98 ;
	7'h0f :
		TR_179 = TR_98 ;
	7'h10 :
		TR_179 = TR_98 ;
	7'h11 :
		TR_179 = TR_98 ;
	7'h12 :
		TR_179 = TR_98 ;
	7'h13 :
		TR_179 = TR_98 ;
	7'h14 :
		TR_179 = TR_98 ;
	7'h15 :
		TR_179 = TR_98 ;
	7'h16 :
		TR_179 = TR_98 ;
	7'h17 :
		TR_179 = TR_98 ;
	7'h18 :
		TR_179 = TR_98 ;
	7'h19 :
		TR_179 = TR_98 ;
	7'h1a :
		TR_179 = TR_98 ;
	7'h1b :
		TR_179 = TR_98 ;
	7'h1c :
		TR_179 = TR_98 ;
	7'h1d :
		TR_179 = TR_98 ;
	7'h1e :
		TR_179 = TR_98 ;
	7'h1f :
		TR_179 = TR_98 ;
	7'h20 :
		TR_179 = TR_98 ;
	7'h21 :
		TR_179 = TR_98 ;
	7'h22 :
		TR_179 = TR_98 ;
	7'h23 :
		TR_179 = TR_98 ;
	7'h24 :
		TR_179 = TR_98 ;
	7'h25 :
		TR_179 = TR_98 ;
	7'h26 :
		TR_179 = TR_98 ;
	7'h27 :
		TR_179 = TR_98 ;
	7'h28 :
		TR_179 = TR_98 ;
	7'h29 :
		TR_179 = TR_98 ;
	7'h2a :
		TR_179 = TR_98 ;
	7'h2b :
		TR_179 = TR_98 ;
	7'h2c :
		TR_179 = TR_98 ;
	7'h2d :
		TR_179 = TR_98 ;
	7'h2e :
		TR_179 = TR_98 ;
	7'h2f :
		TR_179 = TR_98 ;
	7'h30 :
		TR_179 = TR_98 ;
	7'h31 :
		TR_179 = TR_98 ;
	7'h32 :
		TR_179 = TR_98 ;
	7'h33 :
		TR_179 = TR_98 ;
	7'h34 :
		TR_179 = TR_98 ;
	7'h35 :
		TR_179 = TR_98 ;
	7'h36 :
		TR_179 = TR_98 ;
	7'h37 :
		TR_179 = TR_98 ;
	7'h38 :
		TR_179 = TR_98 ;
	7'h39 :
		TR_179 = TR_98 ;
	7'h3a :
		TR_179 = TR_98 ;
	7'h3b :
		TR_179 = TR_98 ;
	7'h3c :
		TR_179 = TR_98 ;
	7'h3d :
		TR_179 = TR_98 ;
	7'h3e :
		TR_179 = TR_98 ;
	7'h3f :
		TR_179 = TR_98 ;
	7'h40 :
		TR_179 = TR_98 ;
	7'h41 :
		TR_179 = TR_98 ;
	7'h42 :
		TR_179 = TR_98 ;
	7'h43 :
		TR_179 = TR_98 ;
	7'h44 :
		TR_179 = TR_98 ;
	7'h45 :
		TR_179 = TR_98 ;
	7'h46 :
		TR_179 = TR_98 ;
	7'h47 :
		TR_179 = TR_98 ;
	7'h48 :
		TR_179 = TR_98 ;
	7'h49 :
		TR_179 = TR_98 ;
	7'h4a :
		TR_179 = TR_98 ;
	7'h4b :
		TR_179 = TR_98 ;
	7'h4c :
		TR_179 = TR_98 ;
	7'h4d :
		TR_179 = TR_98 ;
	7'h4e :
		TR_179 = TR_98 ;
	7'h4f :
		TR_179 = TR_98 ;
	7'h50 :
		TR_179 = TR_98 ;
	7'h51 :
		TR_179 = TR_98 ;
	7'h52 :
		TR_179 = TR_98 ;
	7'h53 :
		TR_179 = TR_98 ;
	7'h54 :
		TR_179 = TR_98 ;
	7'h55 :
		TR_179 = TR_98 ;
	7'h56 :
		TR_179 = 9'h000 ;	// line#=../rle.cpp:80
	7'h57 :
		TR_179 = TR_98 ;
	7'h58 :
		TR_179 = TR_98 ;
	7'h59 :
		TR_179 = TR_98 ;
	7'h5a :
		TR_179 = TR_98 ;
	7'h5b :
		TR_179 = TR_98 ;
	7'h5c :
		TR_179 = TR_98 ;
	7'h5d :
		TR_179 = TR_98 ;
	7'h5e :
		TR_179 = TR_98 ;
	7'h5f :
		TR_179 = TR_98 ;
	7'h60 :
		TR_179 = TR_98 ;
	7'h61 :
		TR_179 = TR_98 ;
	7'h62 :
		TR_179 = TR_98 ;
	7'h63 :
		TR_179 = TR_98 ;
	7'h64 :
		TR_179 = TR_98 ;
	7'h65 :
		TR_179 = TR_98 ;
	7'h66 :
		TR_179 = TR_98 ;
	7'h67 :
		TR_179 = TR_98 ;
	7'h68 :
		TR_179 = TR_98 ;
	7'h69 :
		TR_179 = TR_98 ;
	7'h6a :
		TR_179 = TR_98 ;
	7'h6b :
		TR_179 = TR_98 ;
	7'h6c :
		TR_179 = TR_98 ;
	7'h6d :
		TR_179 = TR_98 ;
	7'h6e :
		TR_179 = TR_98 ;
	7'h6f :
		TR_179 = TR_98 ;
	7'h70 :
		TR_179 = TR_98 ;
	7'h71 :
		TR_179 = TR_98 ;
	7'h72 :
		TR_179 = TR_98 ;
	7'h73 :
		TR_179 = TR_98 ;
	7'h74 :
		TR_179 = TR_98 ;
	7'h75 :
		TR_179 = TR_98 ;
	7'h76 :
		TR_179 = TR_98 ;
	7'h77 :
		TR_179 = TR_98 ;
	7'h78 :
		TR_179 = TR_98 ;
	7'h79 :
		TR_179 = TR_98 ;
	7'h7a :
		TR_179 = TR_98 ;
	7'h7b :
		TR_179 = TR_98 ;
	7'h7c :
		TR_179 = TR_98 ;
	7'h7d :
		TR_179 = TR_98 ;
	7'h7e :
		TR_179 = TR_98 ;
	7'h7f :
		TR_179 = TR_98 ;
	default :
		TR_179 = 9'hx ;
	endcase
always @ ( TR_179 or U_173 or sub8u_71ot or U_183 or RG_rl_172 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_86_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h56 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_86_t = ( ( { 9{ M_180 } } & RG_rl_172 )
		| ( { 9{ U_173 } } & TR_179 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_86_en = ( M_180 | RG_rl_86_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_86_en )
		RG_rl_86 <= RG_rl_86_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_99 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_178 = TR_99 ;
	7'h01 :
		TR_178 = TR_99 ;
	7'h02 :
		TR_178 = TR_99 ;
	7'h03 :
		TR_178 = TR_99 ;
	7'h04 :
		TR_178 = TR_99 ;
	7'h05 :
		TR_178 = TR_99 ;
	7'h06 :
		TR_178 = TR_99 ;
	7'h07 :
		TR_178 = TR_99 ;
	7'h08 :
		TR_178 = TR_99 ;
	7'h09 :
		TR_178 = TR_99 ;
	7'h0a :
		TR_178 = TR_99 ;
	7'h0b :
		TR_178 = TR_99 ;
	7'h0c :
		TR_178 = TR_99 ;
	7'h0d :
		TR_178 = TR_99 ;
	7'h0e :
		TR_178 = TR_99 ;
	7'h0f :
		TR_178 = TR_99 ;
	7'h10 :
		TR_178 = TR_99 ;
	7'h11 :
		TR_178 = TR_99 ;
	7'h12 :
		TR_178 = TR_99 ;
	7'h13 :
		TR_178 = TR_99 ;
	7'h14 :
		TR_178 = TR_99 ;
	7'h15 :
		TR_178 = TR_99 ;
	7'h16 :
		TR_178 = TR_99 ;
	7'h17 :
		TR_178 = TR_99 ;
	7'h18 :
		TR_178 = TR_99 ;
	7'h19 :
		TR_178 = TR_99 ;
	7'h1a :
		TR_178 = TR_99 ;
	7'h1b :
		TR_178 = TR_99 ;
	7'h1c :
		TR_178 = TR_99 ;
	7'h1d :
		TR_178 = TR_99 ;
	7'h1e :
		TR_178 = TR_99 ;
	7'h1f :
		TR_178 = TR_99 ;
	7'h20 :
		TR_178 = TR_99 ;
	7'h21 :
		TR_178 = TR_99 ;
	7'h22 :
		TR_178 = TR_99 ;
	7'h23 :
		TR_178 = TR_99 ;
	7'h24 :
		TR_178 = TR_99 ;
	7'h25 :
		TR_178 = TR_99 ;
	7'h26 :
		TR_178 = TR_99 ;
	7'h27 :
		TR_178 = TR_99 ;
	7'h28 :
		TR_178 = TR_99 ;
	7'h29 :
		TR_178 = TR_99 ;
	7'h2a :
		TR_178 = TR_99 ;
	7'h2b :
		TR_178 = TR_99 ;
	7'h2c :
		TR_178 = TR_99 ;
	7'h2d :
		TR_178 = TR_99 ;
	7'h2e :
		TR_178 = TR_99 ;
	7'h2f :
		TR_178 = TR_99 ;
	7'h30 :
		TR_178 = TR_99 ;
	7'h31 :
		TR_178 = TR_99 ;
	7'h32 :
		TR_178 = TR_99 ;
	7'h33 :
		TR_178 = TR_99 ;
	7'h34 :
		TR_178 = TR_99 ;
	7'h35 :
		TR_178 = TR_99 ;
	7'h36 :
		TR_178 = TR_99 ;
	7'h37 :
		TR_178 = TR_99 ;
	7'h38 :
		TR_178 = TR_99 ;
	7'h39 :
		TR_178 = TR_99 ;
	7'h3a :
		TR_178 = TR_99 ;
	7'h3b :
		TR_178 = TR_99 ;
	7'h3c :
		TR_178 = TR_99 ;
	7'h3d :
		TR_178 = TR_99 ;
	7'h3e :
		TR_178 = TR_99 ;
	7'h3f :
		TR_178 = TR_99 ;
	7'h40 :
		TR_178 = TR_99 ;
	7'h41 :
		TR_178 = TR_99 ;
	7'h42 :
		TR_178 = TR_99 ;
	7'h43 :
		TR_178 = TR_99 ;
	7'h44 :
		TR_178 = TR_99 ;
	7'h45 :
		TR_178 = TR_99 ;
	7'h46 :
		TR_178 = TR_99 ;
	7'h47 :
		TR_178 = TR_99 ;
	7'h48 :
		TR_178 = TR_99 ;
	7'h49 :
		TR_178 = TR_99 ;
	7'h4a :
		TR_178 = TR_99 ;
	7'h4b :
		TR_178 = TR_99 ;
	7'h4c :
		TR_178 = TR_99 ;
	7'h4d :
		TR_178 = TR_99 ;
	7'h4e :
		TR_178 = TR_99 ;
	7'h4f :
		TR_178 = TR_99 ;
	7'h50 :
		TR_178 = TR_99 ;
	7'h51 :
		TR_178 = TR_99 ;
	7'h52 :
		TR_178 = TR_99 ;
	7'h53 :
		TR_178 = TR_99 ;
	7'h54 :
		TR_178 = TR_99 ;
	7'h55 :
		TR_178 = TR_99 ;
	7'h56 :
		TR_178 = TR_99 ;
	7'h57 :
		TR_178 = 9'h000 ;	// line#=../rle.cpp:80
	7'h58 :
		TR_178 = TR_99 ;
	7'h59 :
		TR_178 = TR_99 ;
	7'h5a :
		TR_178 = TR_99 ;
	7'h5b :
		TR_178 = TR_99 ;
	7'h5c :
		TR_178 = TR_99 ;
	7'h5d :
		TR_178 = TR_99 ;
	7'h5e :
		TR_178 = TR_99 ;
	7'h5f :
		TR_178 = TR_99 ;
	7'h60 :
		TR_178 = TR_99 ;
	7'h61 :
		TR_178 = TR_99 ;
	7'h62 :
		TR_178 = TR_99 ;
	7'h63 :
		TR_178 = TR_99 ;
	7'h64 :
		TR_178 = TR_99 ;
	7'h65 :
		TR_178 = TR_99 ;
	7'h66 :
		TR_178 = TR_99 ;
	7'h67 :
		TR_178 = TR_99 ;
	7'h68 :
		TR_178 = TR_99 ;
	7'h69 :
		TR_178 = TR_99 ;
	7'h6a :
		TR_178 = TR_99 ;
	7'h6b :
		TR_178 = TR_99 ;
	7'h6c :
		TR_178 = TR_99 ;
	7'h6d :
		TR_178 = TR_99 ;
	7'h6e :
		TR_178 = TR_99 ;
	7'h6f :
		TR_178 = TR_99 ;
	7'h70 :
		TR_178 = TR_99 ;
	7'h71 :
		TR_178 = TR_99 ;
	7'h72 :
		TR_178 = TR_99 ;
	7'h73 :
		TR_178 = TR_99 ;
	7'h74 :
		TR_178 = TR_99 ;
	7'h75 :
		TR_178 = TR_99 ;
	7'h76 :
		TR_178 = TR_99 ;
	7'h77 :
		TR_178 = TR_99 ;
	7'h78 :
		TR_178 = TR_99 ;
	7'h79 :
		TR_178 = TR_99 ;
	7'h7a :
		TR_178 = TR_99 ;
	7'h7b :
		TR_178 = TR_99 ;
	7'h7c :
		TR_178 = TR_99 ;
	7'h7d :
		TR_178 = TR_99 ;
	7'h7e :
		TR_178 = TR_99 ;
	7'h7f :
		TR_178 = TR_99 ;
	default :
		TR_178 = 9'hx ;
	endcase
always @ ( TR_178 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_41 or 
	U_174 or RG_rl_172 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_87_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h57 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_87_t = ( ( { 9{ ST1_03d } } & RG_rl_172 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_41 )
		| ( { 9{ U_173 } } & TR_178 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_87_en = ( ST1_03d | U_174 | RG_rl_87_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_87_en )
		RG_rl_87 <= RG_rl_87_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_100 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_177 = TR_100 ;
	7'h01 :
		TR_177 = TR_100 ;
	7'h02 :
		TR_177 = TR_100 ;
	7'h03 :
		TR_177 = TR_100 ;
	7'h04 :
		TR_177 = TR_100 ;
	7'h05 :
		TR_177 = TR_100 ;
	7'h06 :
		TR_177 = TR_100 ;
	7'h07 :
		TR_177 = TR_100 ;
	7'h08 :
		TR_177 = TR_100 ;
	7'h09 :
		TR_177 = TR_100 ;
	7'h0a :
		TR_177 = TR_100 ;
	7'h0b :
		TR_177 = TR_100 ;
	7'h0c :
		TR_177 = TR_100 ;
	7'h0d :
		TR_177 = TR_100 ;
	7'h0e :
		TR_177 = TR_100 ;
	7'h0f :
		TR_177 = TR_100 ;
	7'h10 :
		TR_177 = TR_100 ;
	7'h11 :
		TR_177 = TR_100 ;
	7'h12 :
		TR_177 = TR_100 ;
	7'h13 :
		TR_177 = TR_100 ;
	7'h14 :
		TR_177 = TR_100 ;
	7'h15 :
		TR_177 = TR_100 ;
	7'h16 :
		TR_177 = TR_100 ;
	7'h17 :
		TR_177 = TR_100 ;
	7'h18 :
		TR_177 = TR_100 ;
	7'h19 :
		TR_177 = TR_100 ;
	7'h1a :
		TR_177 = TR_100 ;
	7'h1b :
		TR_177 = TR_100 ;
	7'h1c :
		TR_177 = TR_100 ;
	7'h1d :
		TR_177 = TR_100 ;
	7'h1e :
		TR_177 = TR_100 ;
	7'h1f :
		TR_177 = TR_100 ;
	7'h20 :
		TR_177 = TR_100 ;
	7'h21 :
		TR_177 = TR_100 ;
	7'h22 :
		TR_177 = TR_100 ;
	7'h23 :
		TR_177 = TR_100 ;
	7'h24 :
		TR_177 = TR_100 ;
	7'h25 :
		TR_177 = TR_100 ;
	7'h26 :
		TR_177 = TR_100 ;
	7'h27 :
		TR_177 = TR_100 ;
	7'h28 :
		TR_177 = TR_100 ;
	7'h29 :
		TR_177 = TR_100 ;
	7'h2a :
		TR_177 = TR_100 ;
	7'h2b :
		TR_177 = TR_100 ;
	7'h2c :
		TR_177 = TR_100 ;
	7'h2d :
		TR_177 = TR_100 ;
	7'h2e :
		TR_177 = TR_100 ;
	7'h2f :
		TR_177 = TR_100 ;
	7'h30 :
		TR_177 = TR_100 ;
	7'h31 :
		TR_177 = TR_100 ;
	7'h32 :
		TR_177 = TR_100 ;
	7'h33 :
		TR_177 = TR_100 ;
	7'h34 :
		TR_177 = TR_100 ;
	7'h35 :
		TR_177 = TR_100 ;
	7'h36 :
		TR_177 = TR_100 ;
	7'h37 :
		TR_177 = TR_100 ;
	7'h38 :
		TR_177 = TR_100 ;
	7'h39 :
		TR_177 = TR_100 ;
	7'h3a :
		TR_177 = TR_100 ;
	7'h3b :
		TR_177 = TR_100 ;
	7'h3c :
		TR_177 = TR_100 ;
	7'h3d :
		TR_177 = TR_100 ;
	7'h3e :
		TR_177 = TR_100 ;
	7'h3f :
		TR_177 = TR_100 ;
	7'h40 :
		TR_177 = TR_100 ;
	7'h41 :
		TR_177 = TR_100 ;
	7'h42 :
		TR_177 = TR_100 ;
	7'h43 :
		TR_177 = TR_100 ;
	7'h44 :
		TR_177 = TR_100 ;
	7'h45 :
		TR_177 = TR_100 ;
	7'h46 :
		TR_177 = TR_100 ;
	7'h47 :
		TR_177 = TR_100 ;
	7'h48 :
		TR_177 = TR_100 ;
	7'h49 :
		TR_177 = TR_100 ;
	7'h4a :
		TR_177 = TR_100 ;
	7'h4b :
		TR_177 = TR_100 ;
	7'h4c :
		TR_177 = TR_100 ;
	7'h4d :
		TR_177 = TR_100 ;
	7'h4e :
		TR_177 = TR_100 ;
	7'h4f :
		TR_177 = TR_100 ;
	7'h50 :
		TR_177 = TR_100 ;
	7'h51 :
		TR_177 = TR_100 ;
	7'h52 :
		TR_177 = TR_100 ;
	7'h53 :
		TR_177 = TR_100 ;
	7'h54 :
		TR_177 = TR_100 ;
	7'h55 :
		TR_177 = TR_100 ;
	7'h56 :
		TR_177 = TR_100 ;
	7'h57 :
		TR_177 = TR_100 ;
	7'h58 :
		TR_177 = 9'h000 ;	// line#=../rle.cpp:80
	7'h59 :
		TR_177 = TR_100 ;
	7'h5a :
		TR_177 = TR_100 ;
	7'h5b :
		TR_177 = TR_100 ;
	7'h5c :
		TR_177 = TR_100 ;
	7'h5d :
		TR_177 = TR_100 ;
	7'h5e :
		TR_177 = TR_100 ;
	7'h5f :
		TR_177 = TR_100 ;
	7'h60 :
		TR_177 = TR_100 ;
	7'h61 :
		TR_177 = TR_100 ;
	7'h62 :
		TR_177 = TR_100 ;
	7'h63 :
		TR_177 = TR_100 ;
	7'h64 :
		TR_177 = TR_100 ;
	7'h65 :
		TR_177 = TR_100 ;
	7'h66 :
		TR_177 = TR_100 ;
	7'h67 :
		TR_177 = TR_100 ;
	7'h68 :
		TR_177 = TR_100 ;
	7'h69 :
		TR_177 = TR_100 ;
	7'h6a :
		TR_177 = TR_100 ;
	7'h6b :
		TR_177 = TR_100 ;
	7'h6c :
		TR_177 = TR_100 ;
	7'h6d :
		TR_177 = TR_100 ;
	7'h6e :
		TR_177 = TR_100 ;
	7'h6f :
		TR_177 = TR_100 ;
	7'h70 :
		TR_177 = TR_100 ;
	7'h71 :
		TR_177 = TR_100 ;
	7'h72 :
		TR_177 = TR_100 ;
	7'h73 :
		TR_177 = TR_100 ;
	7'h74 :
		TR_177 = TR_100 ;
	7'h75 :
		TR_177 = TR_100 ;
	7'h76 :
		TR_177 = TR_100 ;
	7'h77 :
		TR_177 = TR_100 ;
	7'h78 :
		TR_177 = TR_100 ;
	7'h79 :
		TR_177 = TR_100 ;
	7'h7a :
		TR_177 = TR_100 ;
	7'h7b :
		TR_177 = TR_100 ;
	7'h7c :
		TR_177 = TR_100 ;
	7'h7d :
		TR_177 = TR_100 ;
	7'h7e :
		TR_177 = TR_100 ;
	7'h7f :
		TR_177 = TR_100 ;
	default :
		TR_177 = 9'hx ;
	endcase
always @ ( TR_177 or U_173 or sub8u_71ot or U_183 or RG_rl_173 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_88_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h58 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_88_t = ( ( { 9{ M_180 } } & RG_rl_173 )
		| ( { 9{ U_173 } } & TR_177 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_88_en = ( M_180 | RG_rl_88_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_88_en )
		RG_rl_88 <= RG_rl_88_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_101 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_176 = TR_101 ;
	7'h01 :
		TR_176 = TR_101 ;
	7'h02 :
		TR_176 = TR_101 ;
	7'h03 :
		TR_176 = TR_101 ;
	7'h04 :
		TR_176 = TR_101 ;
	7'h05 :
		TR_176 = TR_101 ;
	7'h06 :
		TR_176 = TR_101 ;
	7'h07 :
		TR_176 = TR_101 ;
	7'h08 :
		TR_176 = TR_101 ;
	7'h09 :
		TR_176 = TR_101 ;
	7'h0a :
		TR_176 = TR_101 ;
	7'h0b :
		TR_176 = TR_101 ;
	7'h0c :
		TR_176 = TR_101 ;
	7'h0d :
		TR_176 = TR_101 ;
	7'h0e :
		TR_176 = TR_101 ;
	7'h0f :
		TR_176 = TR_101 ;
	7'h10 :
		TR_176 = TR_101 ;
	7'h11 :
		TR_176 = TR_101 ;
	7'h12 :
		TR_176 = TR_101 ;
	7'h13 :
		TR_176 = TR_101 ;
	7'h14 :
		TR_176 = TR_101 ;
	7'h15 :
		TR_176 = TR_101 ;
	7'h16 :
		TR_176 = TR_101 ;
	7'h17 :
		TR_176 = TR_101 ;
	7'h18 :
		TR_176 = TR_101 ;
	7'h19 :
		TR_176 = TR_101 ;
	7'h1a :
		TR_176 = TR_101 ;
	7'h1b :
		TR_176 = TR_101 ;
	7'h1c :
		TR_176 = TR_101 ;
	7'h1d :
		TR_176 = TR_101 ;
	7'h1e :
		TR_176 = TR_101 ;
	7'h1f :
		TR_176 = TR_101 ;
	7'h20 :
		TR_176 = TR_101 ;
	7'h21 :
		TR_176 = TR_101 ;
	7'h22 :
		TR_176 = TR_101 ;
	7'h23 :
		TR_176 = TR_101 ;
	7'h24 :
		TR_176 = TR_101 ;
	7'h25 :
		TR_176 = TR_101 ;
	7'h26 :
		TR_176 = TR_101 ;
	7'h27 :
		TR_176 = TR_101 ;
	7'h28 :
		TR_176 = TR_101 ;
	7'h29 :
		TR_176 = TR_101 ;
	7'h2a :
		TR_176 = TR_101 ;
	7'h2b :
		TR_176 = TR_101 ;
	7'h2c :
		TR_176 = TR_101 ;
	7'h2d :
		TR_176 = TR_101 ;
	7'h2e :
		TR_176 = TR_101 ;
	7'h2f :
		TR_176 = TR_101 ;
	7'h30 :
		TR_176 = TR_101 ;
	7'h31 :
		TR_176 = TR_101 ;
	7'h32 :
		TR_176 = TR_101 ;
	7'h33 :
		TR_176 = TR_101 ;
	7'h34 :
		TR_176 = TR_101 ;
	7'h35 :
		TR_176 = TR_101 ;
	7'h36 :
		TR_176 = TR_101 ;
	7'h37 :
		TR_176 = TR_101 ;
	7'h38 :
		TR_176 = TR_101 ;
	7'h39 :
		TR_176 = TR_101 ;
	7'h3a :
		TR_176 = TR_101 ;
	7'h3b :
		TR_176 = TR_101 ;
	7'h3c :
		TR_176 = TR_101 ;
	7'h3d :
		TR_176 = TR_101 ;
	7'h3e :
		TR_176 = TR_101 ;
	7'h3f :
		TR_176 = TR_101 ;
	7'h40 :
		TR_176 = TR_101 ;
	7'h41 :
		TR_176 = TR_101 ;
	7'h42 :
		TR_176 = TR_101 ;
	7'h43 :
		TR_176 = TR_101 ;
	7'h44 :
		TR_176 = TR_101 ;
	7'h45 :
		TR_176 = TR_101 ;
	7'h46 :
		TR_176 = TR_101 ;
	7'h47 :
		TR_176 = TR_101 ;
	7'h48 :
		TR_176 = TR_101 ;
	7'h49 :
		TR_176 = TR_101 ;
	7'h4a :
		TR_176 = TR_101 ;
	7'h4b :
		TR_176 = TR_101 ;
	7'h4c :
		TR_176 = TR_101 ;
	7'h4d :
		TR_176 = TR_101 ;
	7'h4e :
		TR_176 = TR_101 ;
	7'h4f :
		TR_176 = TR_101 ;
	7'h50 :
		TR_176 = TR_101 ;
	7'h51 :
		TR_176 = TR_101 ;
	7'h52 :
		TR_176 = TR_101 ;
	7'h53 :
		TR_176 = TR_101 ;
	7'h54 :
		TR_176 = TR_101 ;
	7'h55 :
		TR_176 = TR_101 ;
	7'h56 :
		TR_176 = TR_101 ;
	7'h57 :
		TR_176 = TR_101 ;
	7'h58 :
		TR_176 = TR_101 ;
	7'h59 :
		TR_176 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5a :
		TR_176 = TR_101 ;
	7'h5b :
		TR_176 = TR_101 ;
	7'h5c :
		TR_176 = TR_101 ;
	7'h5d :
		TR_176 = TR_101 ;
	7'h5e :
		TR_176 = TR_101 ;
	7'h5f :
		TR_176 = TR_101 ;
	7'h60 :
		TR_176 = TR_101 ;
	7'h61 :
		TR_176 = TR_101 ;
	7'h62 :
		TR_176 = TR_101 ;
	7'h63 :
		TR_176 = TR_101 ;
	7'h64 :
		TR_176 = TR_101 ;
	7'h65 :
		TR_176 = TR_101 ;
	7'h66 :
		TR_176 = TR_101 ;
	7'h67 :
		TR_176 = TR_101 ;
	7'h68 :
		TR_176 = TR_101 ;
	7'h69 :
		TR_176 = TR_101 ;
	7'h6a :
		TR_176 = TR_101 ;
	7'h6b :
		TR_176 = TR_101 ;
	7'h6c :
		TR_176 = TR_101 ;
	7'h6d :
		TR_176 = TR_101 ;
	7'h6e :
		TR_176 = TR_101 ;
	7'h6f :
		TR_176 = TR_101 ;
	7'h70 :
		TR_176 = TR_101 ;
	7'h71 :
		TR_176 = TR_101 ;
	7'h72 :
		TR_176 = TR_101 ;
	7'h73 :
		TR_176 = TR_101 ;
	7'h74 :
		TR_176 = TR_101 ;
	7'h75 :
		TR_176 = TR_101 ;
	7'h76 :
		TR_176 = TR_101 ;
	7'h77 :
		TR_176 = TR_101 ;
	7'h78 :
		TR_176 = TR_101 ;
	7'h79 :
		TR_176 = TR_101 ;
	7'h7a :
		TR_176 = TR_101 ;
	7'h7b :
		TR_176 = TR_101 ;
	7'h7c :
		TR_176 = TR_101 ;
	7'h7d :
		TR_176 = TR_101 ;
	7'h7e :
		TR_176 = TR_101 ;
	7'h7f :
		TR_176 = TR_101 ;
	default :
		TR_176 = 9'hx ;
	endcase
always @ ( TR_176 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_42 or 
	U_174 or RG_rl_173 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_89_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h59 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_89_t = ( ( { 9{ ST1_03d } } & RG_rl_173 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_42 )
		| ( { 9{ U_173 } } & TR_176 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_89_en = ( ST1_03d | U_174 | RG_rl_89_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_89_en )
		RG_rl_89 <= RG_rl_89_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_102 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_175 = TR_102 ;
	7'h01 :
		TR_175 = TR_102 ;
	7'h02 :
		TR_175 = TR_102 ;
	7'h03 :
		TR_175 = TR_102 ;
	7'h04 :
		TR_175 = TR_102 ;
	7'h05 :
		TR_175 = TR_102 ;
	7'h06 :
		TR_175 = TR_102 ;
	7'h07 :
		TR_175 = TR_102 ;
	7'h08 :
		TR_175 = TR_102 ;
	7'h09 :
		TR_175 = TR_102 ;
	7'h0a :
		TR_175 = TR_102 ;
	7'h0b :
		TR_175 = TR_102 ;
	7'h0c :
		TR_175 = TR_102 ;
	7'h0d :
		TR_175 = TR_102 ;
	7'h0e :
		TR_175 = TR_102 ;
	7'h0f :
		TR_175 = TR_102 ;
	7'h10 :
		TR_175 = TR_102 ;
	7'h11 :
		TR_175 = TR_102 ;
	7'h12 :
		TR_175 = TR_102 ;
	7'h13 :
		TR_175 = TR_102 ;
	7'h14 :
		TR_175 = TR_102 ;
	7'h15 :
		TR_175 = TR_102 ;
	7'h16 :
		TR_175 = TR_102 ;
	7'h17 :
		TR_175 = TR_102 ;
	7'h18 :
		TR_175 = TR_102 ;
	7'h19 :
		TR_175 = TR_102 ;
	7'h1a :
		TR_175 = TR_102 ;
	7'h1b :
		TR_175 = TR_102 ;
	7'h1c :
		TR_175 = TR_102 ;
	7'h1d :
		TR_175 = TR_102 ;
	7'h1e :
		TR_175 = TR_102 ;
	7'h1f :
		TR_175 = TR_102 ;
	7'h20 :
		TR_175 = TR_102 ;
	7'h21 :
		TR_175 = TR_102 ;
	7'h22 :
		TR_175 = TR_102 ;
	7'h23 :
		TR_175 = TR_102 ;
	7'h24 :
		TR_175 = TR_102 ;
	7'h25 :
		TR_175 = TR_102 ;
	7'h26 :
		TR_175 = TR_102 ;
	7'h27 :
		TR_175 = TR_102 ;
	7'h28 :
		TR_175 = TR_102 ;
	7'h29 :
		TR_175 = TR_102 ;
	7'h2a :
		TR_175 = TR_102 ;
	7'h2b :
		TR_175 = TR_102 ;
	7'h2c :
		TR_175 = TR_102 ;
	7'h2d :
		TR_175 = TR_102 ;
	7'h2e :
		TR_175 = TR_102 ;
	7'h2f :
		TR_175 = TR_102 ;
	7'h30 :
		TR_175 = TR_102 ;
	7'h31 :
		TR_175 = TR_102 ;
	7'h32 :
		TR_175 = TR_102 ;
	7'h33 :
		TR_175 = TR_102 ;
	7'h34 :
		TR_175 = TR_102 ;
	7'h35 :
		TR_175 = TR_102 ;
	7'h36 :
		TR_175 = TR_102 ;
	7'h37 :
		TR_175 = TR_102 ;
	7'h38 :
		TR_175 = TR_102 ;
	7'h39 :
		TR_175 = TR_102 ;
	7'h3a :
		TR_175 = TR_102 ;
	7'h3b :
		TR_175 = TR_102 ;
	7'h3c :
		TR_175 = TR_102 ;
	7'h3d :
		TR_175 = TR_102 ;
	7'h3e :
		TR_175 = TR_102 ;
	7'h3f :
		TR_175 = TR_102 ;
	7'h40 :
		TR_175 = TR_102 ;
	7'h41 :
		TR_175 = TR_102 ;
	7'h42 :
		TR_175 = TR_102 ;
	7'h43 :
		TR_175 = TR_102 ;
	7'h44 :
		TR_175 = TR_102 ;
	7'h45 :
		TR_175 = TR_102 ;
	7'h46 :
		TR_175 = TR_102 ;
	7'h47 :
		TR_175 = TR_102 ;
	7'h48 :
		TR_175 = TR_102 ;
	7'h49 :
		TR_175 = TR_102 ;
	7'h4a :
		TR_175 = TR_102 ;
	7'h4b :
		TR_175 = TR_102 ;
	7'h4c :
		TR_175 = TR_102 ;
	7'h4d :
		TR_175 = TR_102 ;
	7'h4e :
		TR_175 = TR_102 ;
	7'h4f :
		TR_175 = TR_102 ;
	7'h50 :
		TR_175 = TR_102 ;
	7'h51 :
		TR_175 = TR_102 ;
	7'h52 :
		TR_175 = TR_102 ;
	7'h53 :
		TR_175 = TR_102 ;
	7'h54 :
		TR_175 = TR_102 ;
	7'h55 :
		TR_175 = TR_102 ;
	7'h56 :
		TR_175 = TR_102 ;
	7'h57 :
		TR_175 = TR_102 ;
	7'h58 :
		TR_175 = TR_102 ;
	7'h59 :
		TR_175 = TR_102 ;
	7'h5a :
		TR_175 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5b :
		TR_175 = TR_102 ;
	7'h5c :
		TR_175 = TR_102 ;
	7'h5d :
		TR_175 = TR_102 ;
	7'h5e :
		TR_175 = TR_102 ;
	7'h5f :
		TR_175 = TR_102 ;
	7'h60 :
		TR_175 = TR_102 ;
	7'h61 :
		TR_175 = TR_102 ;
	7'h62 :
		TR_175 = TR_102 ;
	7'h63 :
		TR_175 = TR_102 ;
	7'h64 :
		TR_175 = TR_102 ;
	7'h65 :
		TR_175 = TR_102 ;
	7'h66 :
		TR_175 = TR_102 ;
	7'h67 :
		TR_175 = TR_102 ;
	7'h68 :
		TR_175 = TR_102 ;
	7'h69 :
		TR_175 = TR_102 ;
	7'h6a :
		TR_175 = TR_102 ;
	7'h6b :
		TR_175 = TR_102 ;
	7'h6c :
		TR_175 = TR_102 ;
	7'h6d :
		TR_175 = TR_102 ;
	7'h6e :
		TR_175 = TR_102 ;
	7'h6f :
		TR_175 = TR_102 ;
	7'h70 :
		TR_175 = TR_102 ;
	7'h71 :
		TR_175 = TR_102 ;
	7'h72 :
		TR_175 = TR_102 ;
	7'h73 :
		TR_175 = TR_102 ;
	7'h74 :
		TR_175 = TR_102 ;
	7'h75 :
		TR_175 = TR_102 ;
	7'h76 :
		TR_175 = TR_102 ;
	7'h77 :
		TR_175 = TR_102 ;
	7'h78 :
		TR_175 = TR_102 ;
	7'h79 :
		TR_175 = TR_102 ;
	7'h7a :
		TR_175 = TR_102 ;
	7'h7b :
		TR_175 = TR_102 ;
	7'h7c :
		TR_175 = TR_102 ;
	7'h7d :
		TR_175 = TR_102 ;
	7'h7e :
		TR_175 = TR_102 ;
	7'h7f :
		TR_175 = TR_102 ;
	default :
		TR_175 = 9'hx ;
	endcase
always @ ( TR_175 or U_173 or sub8u_71ot or U_183 or RG_rl_174 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_90_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h5a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_90_t = ( ( { 9{ M_180 } } & RG_rl_174 )
		| ( { 9{ U_173 } } & TR_175 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_90_en = ( M_180 | RG_rl_90_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_90_en )
		RG_rl_90 <= RG_rl_90_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_103 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_174 = TR_103 ;
	7'h01 :
		TR_174 = TR_103 ;
	7'h02 :
		TR_174 = TR_103 ;
	7'h03 :
		TR_174 = TR_103 ;
	7'h04 :
		TR_174 = TR_103 ;
	7'h05 :
		TR_174 = TR_103 ;
	7'h06 :
		TR_174 = TR_103 ;
	7'h07 :
		TR_174 = TR_103 ;
	7'h08 :
		TR_174 = TR_103 ;
	7'h09 :
		TR_174 = TR_103 ;
	7'h0a :
		TR_174 = TR_103 ;
	7'h0b :
		TR_174 = TR_103 ;
	7'h0c :
		TR_174 = TR_103 ;
	7'h0d :
		TR_174 = TR_103 ;
	7'h0e :
		TR_174 = TR_103 ;
	7'h0f :
		TR_174 = TR_103 ;
	7'h10 :
		TR_174 = TR_103 ;
	7'h11 :
		TR_174 = TR_103 ;
	7'h12 :
		TR_174 = TR_103 ;
	7'h13 :
		TR_174 = TR_103 ;
	7'h14 :
		TR_174 = TR_103 ;
	7'h15 :
		TR_174 = TR_103 ;
	7'h16 :
		TR_174 = TR_103 ;
	7'h17 :
		TR_174 = TR_103 ;
	7'h18 :
		TR_174 = TR_103 ;
	7'h19 :
		TR_174 = TR_103 ;
	7'h1a :
		TR_174 = TR_103 ;
	7'h1b :
		TR_174 = TR_103 ;
	7'h1c :
		TR_174 = TR_103 ;
	7'h1d :
		TR_174 = TR_103 ;
	7'h1e :
		TR_174 = TR_103 ;
	7'h1f :
		TR_174 = TR_103 ;
	7'h20 :
		TR_174 = TR_103 ;
	7'h21 :
		TR_174 = TR_103 ;
	7'h22 :
		TR_174 = TR_103 ;
	7'h23 :
		TR_174 = TR_103 ;
	7'h24 :
		TR_174 = TR_103 ;
	7'h25 :
		TR_174 = TR_103 ;
	7'h26 :
		TR_174 = TR_103 ;
	7'h27 :
		TR_174 = TR_103 ;
	7'h28 :
		TR_174 = TR_103 ;
	7'h29 :
		TR_174 = TR_103 ;
	7'h2a :
		TR_174 = TR_103 ;
	7'h2b :
		TR_174 = TR_103 ;
	7'h2c :
		TR_174 = TR_103 ;
	7'h2d :
		TR_174 = TR_103 ;
	7'h2e :
		TR_174 = TR_103 ;
	7'h2f :
		TR_174 = TR_103 ;
	7'h30 :
		TR_174 = TR_103 ;
	7'h31 :
		TR_174 = TR_103 ;
	7'h32 :
		TR_174 = TR_103 ;
	7'h33 :
		TR_174 = TR_103 ;
	7'h34 :
		TR_174 = TR_103 ;
	7'h35 :
		TR_174 = TR_103 ;
	7'h36 :
		TR_174 = TR_103 ;
	7'h37 :
		TR_174 = TR_103 ;
	7'h38 :
		TR_174 = TR_103 ;
	7'h39 :
		TR_174 = TR_103 ;
	7'h3a :
		TR_174 = TR_103 ;
	7'h3b :
		TR_174 = TR_103 ;
	7'h3c :
		TR_174 = TR_103 ;
	7'h3d :
		TR_174 = TR_103 ;
	7'h3e :
		TR_174 = TR_103 ;
	7'h3f :
		TR_174 = TR_103 ;
	7'h40 :
		TR_174 = TR_103 ;
	7'h41 :
		TR_174 = TR_103 ;
	7'h42 :
		TR_174 = TR_103 ;
	7'h43 :
		TR_174 = TR_103 ;
	7'h44 :
		TR_174 = TR_103 ;
	7'h45 :
		TR_174 = TR_103 ;
	7'h46 :
		TR_174 = TR_103 ;
	7'h47 :
		TR_174 = TR_103 ;
	7'h48 :
		TR_174 = TR_103 ;
	7'h49 :
		TR_174 = TR_103 ;
	7'h4a :
		TR_174 = TR_103 ;
	7'h4b :
		TR_174 = TR_103 ;
	7'h4c :
		TR_174 = TR_103 ;
	7'h4d :
		TR_174 = TR_103 ;
	7'h4e :
		TR_174 = TR_103 ;
	7'h4f :
		TR_174 = TR_103 ;
	7'h50 :
		TR_174 = TR_103 ;
	7'h51 :
		TR_174 = TR_103 ;
	7'h52 :
		TR_174 = TR_103 ;
	7'h53 :
		TR_174 = TR_103 ;
	7'h54 :
		TR_174 = TR_103 ;
	7'h55 :
		TR_174 = TR_103 ;
	7'h56 :
		TR_174 = TR_103 ;
	7'h57 :
		TR_174 = TR_103 ;
	7'h58 :
		TR_174 = TR_103 ;
	7'h59 :
		TR_174 = TR_103 ;
	7'h5a :
		TR_174 = TR_103 ;
	7'h5b :
		TR_174 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5c :
		TR_174 = TR_103 ;
	7'h5d :
		TR_174 = TR_103 ;
	7'h5e :
		TR_174 = TR_103 ;
	7'h5f :
		TR_174 = TR_103 ;
	7'h60 :
		TR_174 = TR_103 ;
	7'h61 :
		TR_174 = TR_103 ;
	7'h62 :
		TR_174 = TR_103 ;
	7'h63 :
		TR_174 = TR_103 ;
	7'h64 :
		TR_174 = TR_103 ;
	7'h65 :
		TR_174 = TR_103 ;
	7'h66 :
		TR_174 = TR_103 ;
	7'h67 :
		TR_174 = TR_103 ;
	7'h68 :
		TR_174 = TR_103 ;
	7'h69 :
		TR_174 = TR_103 ;
	7'h6a :
		TR_174 = TR_103 ;
	7'h6b :
		TR_174 = TR_103 ;
	7'h6c :
		TR_174 = TR_103 ;
	7'h6d :
		TR_174 = TR_103 ;
	7'h6e :
		TR_174 = TR_103 ;
	7'h6f :
		TR_174 = TR_103 ;
	7'h70 :
		TR_174 = TR_103 ;
	7'h71 :
		TR_174 = TR_103 ;
	7'h72 :
		TR_174 = TR_103 ;
	7'h73 :
		TR_174 = TR_103 ;
	7'h74 :
		TR_174 = TR_103 ;
	7'h75 :
		TR_174 = TR_103 ;
	7'h76 :
		TR_174 = TR_103 ;
	7'h77 :
		TR_174 = TR_103 ;
	7'h78 :
		TR_174 = TR_103 ;
	7'h79 :
		TR_174 = TR_103 ;
	7'h7a :
		TR_174 = TR_103 ;
	7'h7b :
		TR_174 = TR_103 ;
	7'h7c :
		TR_174 = TR_103 ;
	7'h7d :
		TR_174 = TR_103 ;
	7'h7e :
		TR_174 = TR_103 ;
	7'h7f :
		TR_174 = TR_103 ;
	default :
		TR_174 = 9'hx ;
	endcase
always @ ( TR_174 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_43 or 
	U_174 or RG_rl_174 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_91_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h5b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_91_t = ( ( { 9{ ST1_03d } } & RG_rl_174 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_43 )
		| ( { 9{ U_173 } } & TR_174 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_91_en = ( ST1_03d | U_174 | RG_rl_91_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_91_en )
		RG_rl_91 <= RG_rl_91_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_104 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_173 = TR_104 ;
	7'h01 :
		TR_173 = TR_104 ;
	7'h02 :
		TR_173 = TR_104 ;
	7'h03 :
		TR_173 = TR_104 ;
	7'h04 :
		TR_173 = TR_104 ;
	7'h05 :
		TR_173 = TR_104 ;
	7'h06 :
		TR_173 = TR_104 ;
	7'h07 :
		TR_173 = TR_104 ;
	7'h08 :
		TR_173 = TR_104 ;
	7'h09 :
		TR_173 = TR_104 ;
	7'h0a :
		TR_173 = TR_104 ;
	7'h0b :
		TR_173 = TR_104 ;
	7'h0c :
		TR_173 = TR_104 ;
	7'h0d :
		TR_173 = TR_104 ;
	7'h0e :
		TR_173 = TR_104 ;
	7'h0f :
		TR_173 = TR_104 ;
	7'h10 :
		TR_173 = TR_104 ;
	7'h11 :
		TR_173 = TR_104 ;
	7'h12 :
		TR_173 = TR_104 ;
	7'h13 :
		TR_173 = TR_104 ;
	7'h14 :
		TR_173 = TR_104 ;
	7'h15 :
		TR_173 = TR_104 ;
	7'h16 :
		TR_173 = TR_104 ;
	7'h17 :
		TR_173 = TR_104 ;
	7'h18 :
		TR_173 = TR_104 ;
	7'h19 :
		TR_173 = TR_104 ;
	7'h1a :
		TR_173 = TR_104 ;
	7'h1b :
		TR_173 = TR_104 ;
	7'h1c :
		TR_173 = TR_104 ;
	7'h1d :
		TR_173 = TR_104 ;
	7'h1e :
		TR_173 = TR_104 ;
	7'h1f :
		TR_173 = TR_104 ;
	7'h20 :
		TR_173 = TR_104 ;
	7'h21 :
		TR_173 = TR_104 ;
	7'h22 :
		TR_173 = TR_104 ;
	7'h23 :
		TR_173 = TR_104 ;
	7'h24 :
		TR_173 = TR_104 ;
	7'h25 :
		TR_173 = TR_104 ;
	7'h26 :
		TR_173 = TR_104 ;
	7'h27 :
		TR_173 = TR_104 ;
	7'h28 :
		TR_173 = TR_104 ;
	7'h29 :
		TR_173 = TR_104 ;
	7'h2a :
		TR_173 = TR_104 ;
	7'h2b :
		TR_173 = TR_104 ;
	7'h2c :
		TR_173 = TR_104 ;
	7'h2d :
		TR_173 = TR_104 ;
	7'h2e :
		TR_173 = TR_104 ;
	7'h2f :
		TR_173 = TR_104 ;
	7'h30 :
		TR_173 = TR_104 ;
	7'h31 :
		TR_173 = TR_104 ;
	7'h32 :
		TR_173 = TR_104 ;
	7'h33 :
		TR_173 = TR_104 ;
	7'h34 :
		TR_173 = TR_104 ;
	7'h35 :
		TR_173 = TR_104 ;
	7'h36 :
		TR_173 = TR_104 ;
	7'h37 :
		TR_173 = TR_104 ;
	7'h38 :
		TR_173 = TR_104 ;
	7'h39 :
		TR_173 = TR_104 ;
	7'h3a :
		TR_173 = TR_104 ;
	7'h3b :
		TR_173 = TR_104 ;
	7'h3c :
		TR_173 = TR_104 ;
	7'h3d :
		TR_173 = TR_104 ;
	7'h3e :
		TR_173 = TR_104 ;
	7'h3f :
		TR_173 = TR_104 ;
	7'h40 :
		TR_173 = TR_104 ;
	7'h41 :
		TR_173 = TR_104 ;
	7'h42 :
		TR_173 = TR_104 ;
	7'h43 :
		TR_173 = TR_104 ;
	7'h44 :
		TR_173 = TR_104 ;
	7'h45 :
		TR_173 = TR_104 ;
	7'h46 :
		TR_173 = TR_104 ;
	7'h47 :
		TR_173 = TR_104 ;
	7'h48 :
		TR_173 = TR_104 ;
	7'h49 :
		TR_173 = TR_104 ;
	7'h4a :
		TR_173 = TR_104 ;
	7'h4b :
		TR_173 = TR_104 ;
	7'h4c :
		TR_173 = TR_104 ;
	7'h4d :
		TR_173 = TR_104 ;
	7'h4e :
		TR_173 = TR_104 ;
	7'h4f :
		TR_173 = TR_104 ;
	7'h50 :
		TR_173 = TR_104 ;
	7'h51 :
		TR_173 = TR_104 ;
	7'h52 :
		TR_173 = TR_104 ;
	7'h53 :
		TR_173 = TR_104 ;
	7'h54 :
		TR_173 = TR_104 ;
	7'h55 :
		TR_173 = TR_104 ;
	7'h56 :
		TR_173 = TR_104 ;
	7'h57 :
		TR_173 = TR_104 ;
	7'h58 :
		TR_173 = TR_104 ;
	7'h59 :
		TR_173 = TR_104 ;
	7'h5a :
		TR_173 = TR_104 ;
	7'h5b :
		TR_173 = TR_104 ;
	7'h5c :
		TR_173 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5d :
		TR_173 = TR_104 ;
	7'h5e :
		TR_173 = TR_104 ;
	7'h5f :
		TR_173 = TR_104 ;
	7'h60 :
		TR_173 = TR_104 ;
	7'h61 :
		TR_173 = TR_104 ;
	7'h62 :
		TR_173 = TR_104 ;
	7'h63 :
		TR_173 = TR_104 ;
	7'h64 :
		TR_173 = TR_104 ;
	7'h65 :
		TR_173 = TR_104 ;
	7'h66 :
		TR_173 = TR_104 ;
	7'h67 :
		TR_173 = TR_104 ;
	7'h68 :
		TR_173 = TR_104 ;
	7'h69 :
		TR_173 = TR_104 ;
	7'h6a :
		TR_173 = TR_104 ;
	7'h6b :
		TR_173 = TR_104 ;
	7'h6c :
		TR_173 = TR_104 ;
	7'h6d :
		TR_173 = TR_104 ;
	7'h6e :
		TR_173 = TR_104 ;
	7'h6f :
		TR_173 = TR_104 ;
	7'h70 :
		TR_173 = TR_104 ;
	7'h71 :
		TR_173 = TR_104 ;
	7'h72 :
		TR_173 = TR_104 ;
	7'h73 :
		TR_173 = TR_104 ;
	7'h74 :
		TR_173 = TR_104 ;
	7'h75 :
		TR_173 = TR_104 ;
	7'h76 :
		TR_173 = TR_104 ;
	7'h77 :
		TR_173 = TR_104 ;
	7'h78 :
		TR_173 = TR_104 ;
	7'h79 :
		TR_173 = TR_104 ;
	7'h7a :
		TR_173 = TR_104 ;
	7'h7b :
		TR_173 = TR_104 ;
	7'h7c :
		TR_173 = TR_104 ;
	7'h7d :
		TR_173 = TR_104 ;
	7'h7e :
		TR_173 = TR_104 ;
	7'h7f :
		TR_173 = TR_104 ;
	default :
		TR_173 = 9'hx ;
	endcase
always @ ( TR_173 or U_173 or sub8u_71ot or U_183 or RG_rl_175 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_92_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h5c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_92_t = ( ( { 9{ M_180 } } & RG_rl_175 )
		| ( { 9{ U_173 } } & TR_173 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_92_en = ( M_180 | RG_rl_92_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_92_en )
		RG_rl_92 <= RG_rl_92_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_105 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_172 = TR_105 ;
	7'h01 :
		TR_172 = TR_105 ;
	7'h02 :
		TR_172 = TR_105 ;
	7'h03 :
		TR_172 = TR_105 ;
	7'h04 :
		TR_172 = TR_105 ;
	7'h05 :
		TR_172 = TR_105 ;
	7'h06 :
		TR_172 = TR_105 ;
	7'h07 :
		TR_172 = TR_105 ;
	7'h08 :
		TR_172 = TR_105 ;
	7'h09 :
		TR_172 = TR_105 ;
	7'h0a :
		TR_172 = TR_105 ;
	7'h0b :
		TR_172 = TR_105 ;
	7'h0c :
		TR_172 = TR_105 ;
	7'h0d :
		TR_172 = TR_105 ;
	7'h0e :
		TR_172 = TR_105 ;
	7'h0f :
		TR_172 = TR_105 ;
	7'h10 :
		TR_172 = TR_105 ;
	7'h11 :
		TR_172 = TR_105 ;
	7'h12 :
		TR_172 = TR_105 ;
	7'h13 :
		TR_172 = TR_105 ;
	7'h14 :
		TR_172 = TR_105 ;
	7'h15 :
		TR_172 = TR_105 ;
	7'h16 :
		TR_172 = TR_105 ;
	7'h17 :
		TR_172 = TR_105 ;
	7'h18 :
		TR_172 = TR_105 ;
	7'h19 :
		TR_172 = TR_105 ;
	7'h1a :
		TR_172 = TR_105 ;
	7'h1b :
		TR_172 = TR_105 ;
	7'h1c :
		TR_172 = TR_105 ;
	7'h1d :
		TR_172 = TR_105 ;
	7'h1e :
		TR_172 = TR_105 ;
	7'h1f :
		TR_172 = TR_105 ;
	7'h20 :
		TR_172 = TR_105 ;
	7'h21 :
		TR_172 = TR_105 ;
	7'h22 :
		TR_172 = TR_105 ;
	7'h23 :
		TR_172 = TR_105 ;
	7'h24 :
		TR_172 = TR_105 ;
	7'h25 :
		TR_172 = TR_105 ;
	7'h26 :
		TR_172 = TR_105 ;
	7'h27 :
		TR_172 = TR_105 ;
	7'h28 :
		TR_172 = TR_105 ;
	7'h29 :
		TR_172 = TR_105 ;
	7'h2a :
		TR_172 = TR_105 ;
	7'h2b :
		TR_172 = TR_105 ;
	7'h2c :
		TR_172 = TR_105 ;
	7'h2d :
		TR_172 = TR_105 ;
	7'h2e :
		TR_172 = TR_105 ;
	7'h2f :
		TR_172 = TR_105 ;
	7'h30 :
		TR_172 = TR_105 ;
	7'h31 :
		TR_172 = TR_105 ;
	7'h32 :
		TR_172 = TR_105 ;
	7'h33 :
		TR_172 = TR_105 ;
	7'h34 :
		TR_172 = TR_105 ;
	7'h35 :
		TR_172 = TR_105 ;
	7'h36 :
		TR_172 = TR_105 ;
	7'h37 :
		TR_172 = TR_105 ;
	7'h38 :
		TR_172 = TR_105 ;
	7'h39 :
		TR_172 = TR_105 ;
	7'h3a :
		TR_172 = TR_105 ;
	7'h3b :
		TR_172 = TR_105 ;
	7'h3c :
		TR_172 = TR_105 ;
	7'h3d :
		TR_172 = TR_105 ;
	7'h3e :
		TR_172 = TR_105 ;
	7'h3f :
		TR_172 = TR_105 ;
	7'h40 :
		TR_172 = TR_105 ;
	7'h41 :
		TR_172 = TR_105 ;
	7'h42 :
		TR_172 = TR_105 ;
	7'h43 :
		TR_172 = TR_105 ;
	7'h44 :
		TR_172 = TR_105 ;
	7'h45 :
		TR_172 = TR_105 ;
	7'h46 :
		TR_172 = TR_105 ;
	7'h47 :
		TR_172 = TR_105 ;
	7'h48 :
		TR_172 = TR_105 ;
	7'h49 :
		TR_172 = TR_105 ;
	7'h4a :
		TR_172 = TR_105 ;
	7'h4b :
		TR_172 = TR_105 ;
	7'h4c :
		TR_172 = TR_105 ;
	7'h4d :
		TR_172 = TR_105 ;
	7'h4e :
		TR_172 = TR_105 ;
	7'h4f :
		TR_172 = TR_105 ;
	7'h50 :
		TR_172 = TR_105 ;
	7'h51 :
		TR_172 = TR_105 ;
	7'h52 :
		TR_172 = TR_105 ;
	7'h53 :
		TR_172 = TR_105 ;
	7'h54 :
		TR_172 = TR_105 ;
	7'h55 :
		TR_172 = TR_105 ;
	7'h56 :
		TR_172 = TR_105 ;
	7'h57 :
		TR_172 = TR_105 ;
	7'h58 :
		TR_172 = TR_105 ;
	7'h59 :
		TR_172 = TR_105 ;
	7'h5a :
		TR_172 = TR_105 ;
	7'h5b :
		TR_172 = TR_105 ;
	7'h5c :
		TR_172 = TR_105 ;
	7'h5d :
		TR_172 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5e :
		TR_172 = TR_105 ;
	7'h5f :
		TR_172 = TR_105 ;
	7'h60 :
		TR_172 = TR_105 ;
	7'h61 :
		TR_172 = TR_105 ;
	7'h62 :
		TR_172 = TR_105 ;
	7'h63 :
		TR_172 = TR_105 ;
	7'h64 :
		TR_172 = TR_105 ;
	7'h65 :
		TR_172 = TR_105 ;
	7'h66 :
		TR_172 = TR_105 ;
	7'h67 :
		TR_172 = TR_105 ;
	7'h68 :
		TR_172 = TR_105 ;
	7'h69 :
		TR_172 = TR_105 ;
	7'h6a :
		TR_172 = TR_105 ;
	7'h6b :
		TR_172 = TR_105 ;
	7'h6c :
		TR_172 = TR_105 ;
	7'h6d :
		TR_172 = TR_105 ;
	7'h6e :
		TR_172 = TR_105 ;
	7'h6f :
		TR_172 = TR_105 ;
	7'h70 :
		TR_172 = TR_105 ;
	7'h71 :
		TR_172 = TR_105 ;
	7'h72 :
		TR_172 = TR_105 ;
	7'h73 :
		TR_172 = TR_105 ;
	7'h74 :
		TR_172 = TR_105 ;
	7'h75 :
		TR_172 = TR_105 ;
	7'h76 :
		TR_172 = TR_105 ;
	7'h77 :
		TR_172 = TR_105 ;
	7'h78 :
		TR_172 = TR_105 ;
	7'h79 :
		TR_172 = TR_105 ;
	7'h7a :
		TR_172 = TR_105 ;
	7'h7b :
		TR_172 = TR_105 ;
	7'h7c :
		TR_172 = TR_105 ;
	7'h7d :
		TR_172 = TR_105 ;
	7'h7e :
		TR_172 = TR_105 ;
	7'h7f :
		TR_172 = TR_105 ;
	default :
		TR_172 = 9'hx ;
	endcase
always @ ( TR_172 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_44 or 
	U_174 or RG_rl_175 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_93_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h5d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_93_t = ( ( { 9{ ST1_03d } } & RG_rl_175 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_44 )
		| ( { 9{ U_173 } } & TR_172 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_93_en = ( ST1_03d | U_174 | RG_rl_93_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_93_en )
		RG_rl_93 <= RG_rl_93_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_106 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_171 = TR_106 ;
	7'h01 :
		TR_171 = TR_106 ;
	7'h02 :
		TR_171 = TR_106 ;
	7'h03 :
		TR_171 = TR_106 ;
	7'h04 :
		TR_171 = TR_106 ;
	7'h05 :
		TR_171 = TR_106 ;
	7'h06 :
		TR_171 = TR_106 ;
	7'h07 :
		TR_171 = TR_106 ;
	7'h08 :
		TR_171 = TR_106 ;
	7'h09 :
		TR_171 = TR_106 ;
	7'h0a :
		TR_171 = TR_106 ;
	7'h0b :
		TR_171 = TR_106 ;
	7'h0c :
		TR_171 = TR_106 ;
	7'h0d :
		TR_171 = TR_106 ;
	7'h0e :
		TR_171 = TR_106 ;
	7'h0f :
		TR_171 = TR_106 ;
	7'h10 :
		TR_171 = TR_106 ;
	7'h11 :
		TR_171 = TR_106 ;
	7'h12 :
		TR_171 = TR_106 ;
	7'h13 :
		TR_171 = TR_106 ;
	7'h14 :
		TR_171 = TR_106 ;
	7'h15 :
		TR_171 = TR_106 ;
	7'h16 :
		TR_171 = TR_106 ;
	7'h17 :
		TR_171 = TR_106 ;
	7'h18 :
		TR_171 = TR_106 ;
	7'h19 :
		TR_171 = TR_106 ;
	7'h1a :
		TR_171 = TR_106 ;
	7'h1b :
		TR_171 = TR_106 ;
	7'h1c :
		TR_171 = TR_106 ;
	7'h1d :
		TR_171 = TR_106 ;
	7'h1e :
		TR_171 = TR_106 ;
	7'h1f :
		TR_171 = TR_106 ;
	7'h20 :
		TR_171 = TR_106 ;
	7'h21 :
		TR_171 = TR_106 ;
	7'h22 :
		TR_171 = TR_106 ;
	7'h23 :
		TR_171 = TR_106 ;
	7'h24 :
		TR_171 = TR_106 ;
	7'h25 :
		TR_171 = TR_106 ;
	7'h26 :
		TR_171 = TR_106 ;
	7'h27 :
		TR_171 = TR_106 ;
	7'h28 :
		TR_171 = TR_106 ;
	7'h29 :
		TR_171 = TR_106 ;
	7'h2a :
		TR_171 = TR_106 ;
	7'h2b :
		TR_171 = TR_106 ;
	7'h2c :
		TR_171 = TR_106 ;
	7'h2d :
		TR_171 = TR_106 ;
	7'h2e :
		TR_171 = TR_106 ;
	7'h2f :
		TR_171 = TR_106 ;
	7'h30 :
		TR_171 = TR_106 ;
	7'h31 :
		TR_171 = TR_106 ;
	7'h32 :
		TR_171 = TR_106 ;
	7'h33 :
		TR_171 = TR_106 ;
	7'h34 :
		TR_171 = TR_106 ;
	7'h35 :
		TR_171 = TR_106 ;
	7'h36 :
		TR_171 = TR_106 ;
	7'h37 :
		TR_171 = TR_106 ;
	7'h38 :
		TR_171 = TR_106 ;
	7'h39 :
		TR_171 = TR_106 ;
	7'h3a :
		TR_171 = TR_106 ;
	7'h3b :
		TR_171 = TR_106 ;
	7'h3c :
		TR_171 = TR_106 ;
	7'h3d :
		TR_171 = TR_106 ;
	7'h3e :
		TR_171 = TR_106 ;
	7'h3f :
		TR_171 = TR_106 ;
	7'h40 :
		TR_171 = TR_106 ;
	7'h41 :
		TR_171 = TR_106 ;
	7'h42 :
		TR_171 = TR_106 ;
	7'h43 :
		TR_171 = TR_106 ;
	7'h44 :
		TR_171 = TR_106 ;
	7'h45 :
		TR_171 = TR_106 ;
	7'h46 :
		TR_171 = TR_106 ;
	7'h47 :
		TR_171 = TR_106 ;
	7'h48 :
		TR_171 = TR_106 ;
	7'h49 :
		TR_171 = TR_106 ;
	7'h4a :
		TR_171 = TR_106 ;
	7'h4b :
		TR_171 = TR_106 ;
	7'h4c :
		TR_171 = TR_106 ;
	7'h4d :
		TR_171 = TR_106 ;
	7'h4e :
		TR_171 = TR_106 ;
	7'h4f :
		TR_171 = TR_106 ;
	7'h50 :
		TR_171 = TR_106 ;
	7'h51 :
		TR_171 = TR_106 ;
	7'h52 :
		TR_171 = TR_106 ;
	7'h53 :
		TR_171 = TR_106 ;
	7'h54 :
		TR_171 = TR_106 ;
	7'h55 :
		TR_171 = TR_106 ;
	7'h56 :
		TR_171 = TR_106 ;
	7'h57 :
		TR_171 = TR_106 ;
	7'h58 :
		TR_171 = TR_106 ;
	7'h59 :
		TR_171 = TR_106 ;
	7'h5a :
		TR_171 = TR_106 ;
	7'h5b :
		TR_171 = TR_106 ;
	7'h5c :
		TR_171 = TR_106 ;
	7'h5d :
		TR_171 = TR_106 ;
	7'h5e :
		TR_171 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5f :
		TR_171 = TR_106 ;
	7'h60 :
		TR_171 = TR_106 ;
	7'h61 :
		TR_171 = TR_106 ;
	7'h62 :
		TR_171 = TR_106 ;
	7'h63 :
		TR_171 = TR_106 ;
	7'h64 :
		TR_171 = TR_106 ;
	7'h65 :
		TR_171 = TR_106 ;
	7'h66 :
		TR_171 = TR_106 ;
	7'h67 :
		TR_171 = TR_106 ;
	7'h68 :
		TR_171 = TR_106 ;
	7'h69 :
		TR_171 = TR_106 ;
	7'h6a :
		TR_171 = TR_106 ;
	7'h6b :
		TR_171 = TR_106 ;
	7'h6c :
		TR_171 = TR_106 ;
	7'h6d :
		TR_171 = TR_106 ;
	7'h6e :
		TR_171 = TR_106 ;
	7'h6f :
		TR_171 = TR_106 ;
	7'h70 :
		TR_171 = TR_106 ;
	7'h71 :
		TR_171 = TR_106 ;
	7'h72 :
		TR_171 = TR_106 ;
	7'h73 :
		TR_171 = TR_106 ;
	7'h74 :
		TR_171 = TR_106 ;
	7'h75 :
		TR_171 = TR_106 ;
	7'h76 :
		TR_171 = TR_106 ;
	7'h77 :
		TR_171 = TR_106 ;
	7'h78 :
		TR_171 = TR_106 ;
	7'h79 :
		TR_171 = TR_106 ;
	7'h7a :
		TR_171 = TR_106 ;
	7'h7b :
		TR_171 = TR_106 ;
	7'h7c :
		TR_171 = TR_106 ;
	7'h7d :
		TR_171 = TR_106 ;
	7'h7e :
		TR_171 = TR_106 ;
	7'h7f :
		TR_171 = TR_106 ;
	default :
		TR_171 = 9'hx ;
	endcase
always @ ( TR_171 or U_173 or sub8u_71ot or U_183 or RG_rl_176 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_94_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h5e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_94_t = ( ( { 9{ M_180 } } & RG_rl_176 )
		| ( { 9{ U_173 } } & TR_171 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_94_en = ( M_180 | RG_rl_94_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_94_en )
		RG_rl_94 <= RG_rl_94_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_107 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_170 = TR_107 ;
	7'h01 :
		TR_170 = TR_107 ;
	7'h02 :
		TR_170 = TR_107 ;
	7'h03 :
		TR_170 = TR_107 ;
	7'h04 :
		TR_170 = TR_107 ;
	7'h05 :
		TR_170 = TR_107 ;
	7'h06 :
		TR_170 = TR_107 ;
	7'h07 :
		TR_170 = TR_107 ;
	7'h08 :
		TR_170 = TR_107 ;
	7'h09 :
		TR_170 = TR_107 ;
	7'h0a :
		TR_170 = TR_107 ;
	7'h0b :
		TR_170 = TR_107 ;
	7'h0c :
		TR_170 = TR_107 ;
	7'h0d :
		TR_170 = TR_107 ;
	7'h0e :
		TR_170 = TR_107 ;
	7'h0f :
		TR_170 = TR_107 ;
	7'h10 :
		TR_170 = TR_107 ;
	7'h11 :
		TR_170 = TR_107 ;
	7'h12 :
		TR_170 = TR_107 ;
	7'h13 :
		TR_170 = TR_107 ;
	7'h14 :
		TR_170 = TR_107 ;
	7'h15 :
		TR_170 = TR_107 ;
	7'h16 :
		TR_170 = TR_107 ;
	7'h17 :
		TR_170 = TR_107 ;
	7'h18 :
		TR_170 = TR_107 ;
	7'h19 :
		TR_170 = TR_107 ;
	7'h1a :
		TR_170 = TR_107 ;
	7'h1b :
		TR_170 = TR_107 ;
	7'h1c :
		TR_170 = TR_107 ;
	7'h1d :
		TR_170 = TR_107 ;
	7'h1e :
		TR_170 = TR_107 ;
	7'h1f :
		TR_170 = TR_107 ;
	7'h20 :
		TR_170 = TR_107 ;
	7'h21 :
		TR_170 = TR_107 ;
	7'h22 :
		TR_170 = TR_107 ;
	7'h23 :
		TR_170 = TR_107 ;
	7'h24 :
		TR_170 = TR_107 ;
	7'h25 :
		TR_170 = TR_107 ;
	7'h26 :
		TR_170 = TR_107 ;
	7'h27 :
		TR_170 = TR_107 ;
	7'h28 :
		TR_170 = TR_107 ;
	7'h29 :
		TR_170 = TR_107 ;
	7'h2a :
		TR_170 = TR_107 ;
	7'h2b :
		TR_170 = TR_107 ;
	7'h2c :
		TR_170 = TR_107 ;
	7'h2d :
		TR_170 = TR_107 ;
	7'h2e :
		TR_170 = TR_107 ;
	7'h2f :
		TR_170 = TR_107 ;
	7'h30 :
		TR_170 = TR_107 ;
	7'h31 :
		TR_170 = TR_107 ;
	7'h32 :
		TR_170 = TR_107 ;
	7'h33 :
		TR_170 = TR_107 ;
	7'h34 :
		TR_170 = TR_107 ;
	7'h35 :
		TR_170 = TR_107 ;
	7'h36 :
		TR_170 = TR_107 ;
	7'h37 :
		TR_170 = TR_107 ;
	7'h38 :
		TR_170 = TR_107 ;
	7'h39 :
		TR_170 = TR_107 ;
	7'h3a :
		TR_170 = TR_107 ;
	7'h3b :
		TR_170 = TR_107 ;
	7'h3c :
		TR_170 = TR_107 ;
	7'h3d :
		TR_170 = TR_107 ;
	7'h3e :
		TR_170 = TR_107 ;
	7'h3f :
		TR_170 = TR_107 ;
	7'h40 :
		TR_170 = TR_107 ;
	7'h41 :
		TR_170 = TR_107 ;
	7'h42 :
		TR_170 = TR_107 ;
	7'h43 :
		TR_170 = TR_107 ;
	7'h44 :
		TR_170 = TR_107 ;
	7'h45 :
		TR_170 = TR_107 ;
	7'h46 :
		TR_170 = TR_107 ;
	7'h47 :
		TR_170 = TR_107 ;
	7'h48 :
		TR_170 = TR_107 ;
	7'h49 :
		TR_170 = TR_107 ;
	7'h4a :
		TR_170 = TR_107 ;
	7'h4b :
		TR_170 = TR_107 ;
	7'h4c :
		TR_170 = TR_107 ;
	7'h4d :
		TR_170 = TR_107 ;
	7'h4e :
		TR_170 = TR_107 ;
	7'h4f :
		TR_170 = TR_107 ;
	7'h50 :
		TR_170 = TR_107 ;
	7'h51 :
		TR_170 = TR_107 ;
	7'h52 :
		TR_170 = TR_107 ;
	7'h53 :
		TR_170 = TR_107 ;
	7'h54 :
		TR_170 = TR_107 ;
	7'h55 :
		TR_170 = TR_107 ;
	7'h56 :
		TR_170 = TR_107 ;
	7'h57 :
		TR_170 = TR_107 ;
	7'h58 :
		TR_170 = TR_107 ;
	7'h59 :
		TR_170 = TR_107 ;
	7'h5a :
		TR_170 = TR_107 ;
	7'h5b :
		TR_170 = TR_107 ;
	7'h5c :
		TR_170 = TR_107 ;
	7'h5d :
		TR_170 = TR_107 ;
	7'h5e :
		TR_170 = TR_107 ;
	7'h5f :
		TR_170 = 9'h000 ;	// line#=../rle.cpp:80
	7'h60 :
		TR_170 = TR_107 ;
	7'h61 :
		TR_170 = TR_107 ;
	7'h62 :
		TR_170 = TR_107 ;
	7'h63 :
		TR_170 = TR_107 ;
	7'h64 :
		TR_170 = TR_107 ;
	7'h65 :
		TR_170 = TR_107 ;
	7'h66 :
		TR_170 = TR_107 ;
	7'h67 :
		TR_170 = TR_107 ;
	7'h68 :
		TR_170 = TR_107 ;
	7'h69 :
		TR_170 = TR_107 ;
	7'h6a :
		TR_170 = TR_107 ;
	7'h6b :
		TR_170 = TR_107 ;
	7'h6c :
		TR_170 = TR_107 ;
	7'h6d :
		TR_170 = TR_107 ;
	7'h6e :
		TR_170 = TR_107 ;
	7'h6f :
		TR_170 = TR_107 ;
	7'h70 :
		TR_170 = TR_107 ;
	7'h71 :
		TR_170 = TR_107 ;
	7'h72 :
		TR_170 = TR_107 ;
	7'h73 :
		TR_170 = TR_107 ;
	7'h74 :
		TR_170 = TR_107 ;
	7'h75 :
		TR_170 = TR_107 ;
	7'h76 :
		TR_170 = TR_107 ;
	7'h77 :
		TR_170 = TR_107 ;
	7'h78 :
		TR_170 = TR_107 ;
	7'h79 :
		TR_170 = TR_107 ;
	7'h7a :
		TR_170 = TR_107 ;
	7'h7b :
		TR_170 = TR_107 ;
	7'h7c :
		TR_170 = TR_107 ;
	7'h7d :
		TR_170 = TR_107 ;
	7'h7e :
		TR_170 = TR_107 ;
	7'h7f :
		TR_170 = TR_107 ;
	default :
		TR_170 = 9'hx ;
	endcase
always @ ( TR_170 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_45 or 
	U_174 or RG_rl_176 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_95_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h5f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_95_t = ( ( { 9{ ST1_03d } } & RG_rl_176 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_45 )
		| ( { 9{ U_173 } } & TR_170 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_95_en = ( ST1_03d | U_174 | RG_rl_95_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_95_en )
		RG_rl_95 <= RG_rl_95_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_108 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_169 = TR_108 ;
	7'h01 :
		TR_169 = TR_108 ;
	7'h02 :
		TR_169 = TR_108 ;
	7'h03 :
		TR_169 = TR_108 ;
	7'h04 :
		TR_169 = TR_108 ;
	7'h05 :
		TR_169 = TR_108 ;
	7'h06 :
		TR_169 = TR_108 ;
	7'h07 :
		TR_169 = TR_108 ;
	7'h08 :
		TR_169 = TR_108 ;
	7'h09 :
		TR_169 = TR_108 ;
	7'h0a :
		TR_169 = TR_108 ;
	7'h0b :
		TR_169 = TR_108 ;
	7'h0c :
		TR_169 = TR_108 ;
	7'h0d :
		TR_169 = TR_108 ;
	7'h0e :
		TR_169 = TR_108 ;
	7'h0f :
		TR_169 = TR_108 ;
	7'h10 :
		TR_169 = TR_108 ;
	7'h11 :
		TR_169 = TR_108 ;
	7'h12 :
		TR_169 = TR_108 ;
	7'h13 :
		TR_169 = TR_108 ;
	7'h14 :
		TR_169 = TR_108 ;
	7'h15 :
		TR_169 = TR_108 ;
	7'h16 :
		TR_169 = TR_108 ;
	7'h17 :
		TR_169 = TR_108 ;
	7'h18 :
		TR_169 = TR_108 ;
	7'h19 :
		TR_169 = TR_108 ;
	7'h1a :
		TR_169 = TR_108 ;
	7'h1b :
		TR_169 = TR_108 ;
	7'h1c :
		TR_169 = TR_108 ;
	7'h1d :
		TR_169 = TR_108 ;
	7'h1e :
		TR_169 = TR_108 ;
	7'h1f :
		TR_169 = TR_108 ;
	7'h20 :
		TR_169 = TR_108 ;
	7'h21 :
		TR_169 = TR_108 ;
	7'h22 :
		TR_169 = TR_108 ;
	7'h23 :
		TR_169 = TR_108 ;
	7'h24 :
		TR_169 = TR_108 ;
	7'h25 :
		TR_169 = TR_108 ;
	7'h26 :
		TR_169 = TR_108 ;
	7'h27 :
		TR_169 = TR_108 ;
	7'h28 :
		TR_169 = TR_108 ;
	7'h29 :
		TR_169 = TR_108 ;
	7'h2a :
		TR_169 = TR_108 ;
	7'h2b :
		TR_169 = TR_108 ;
	7'h2c :
		TR_169 = TR_108 ;
	7'h2d :
		TR_169 = TR_108 ;
	7'h2e :
		TR_169 = TR_108 ;
	7'h2f :
		TR_169 = TR_108 ;
	7'h30 :
		TR_169 = TR_108 ;
	7'h31 :
		TR_169 = TR_108 ;
	7'h32 :
		TR_169 = TR_108 ;
	7'h33 :
		TR_169 = TR_108 ;
	7'h34 :
		TR_169 = TR_108 ;
	7'h35 :
		TR_169 = TR_108 ;
	7'h36 :
		TR_169 = TR_108 ;
	7'h37 :
		TR_169 = TR_108 ;
	7'h38 :
		TR_169 = TR_108 ;
	7'h39 :
		TR_169 = TR_108 ;
	7'h3a :
		TR_169 = TR_108 ;
	7'h3b :
		TR_169 = TR_108 ;
	7'h3c :
		TR_169 = TR_108 ;
	7'h3d :
		TR_169 = TR_108 ;
	7'h3e :
		TR_169 = TR_108 ;
	7'h3f :
		TR_169 = TR_108 ;
	7'h40 :
		TR_169 = TR_108 ;
	7'h41 :
		TR_169 = TR_108 ;
	7'h42 :
		TR_169 = TR_108 ;
	7'h43 :
		TR_169 = TR_108 ;
	7'h44 :
		TR_169 = TR_108 ;
	7'h45 :
		TR_169 = TR_108 ;
	7'h46 :
		TR_169 = TR_108 ;
	7'h47 :
		TR_169 = TR_108 ;
	7'h48 :
		TR_169 = TR_108 ;
	7'h49 :
		TR_169 = TR_108 ;
	7'h4a :
		TR_169 = TR_108 ;
	7'h4b :
		TR_169 = TR_108 ;
	7'h4c :
		TR_169 = TR_108 ;
	7'h4d :
		TR_169 = TR_108 ;
	7'h4e :
		TR_169 = TR_108 ;
	7'h4f :
		TR_169 = TR_108 ;
	7'h50 :
		TR_169 = TR_108 ;
	7'h51 :
		TR_169 = TR_108 ;
	7'h52 :
		TR_169 = TR_108 ;
	7'h53 :
		TR_169 = TR_108 ;
	7'h54 :
		TR_169 = TR_108 ;
	7'h55 :
		TR_169 = TR_108 ;
	7'h56 :
		TR_169 = TR_108 ;
	7'h57 :
		TR_169 = TR_108 ;
	7'h58 :
		TR_169 = TR_108 ;
	7'h59 :
		TR_169 = TR_108 ;
	7'h5a :
		TR_169 = TR_108 ;
	7'h5b :
		TR_169 = TR_108 ;
	7'h5c :
		TR_169 = TR_108 ;
	7'h5d :
		TR_169 = TR_108 ;
	7'h5e :
		TR_169 = TR_108 ;
	7'h5f :
		TR_169 = TR_108 ;
	7'h60 :
		TR_169 = 9'h000 ;	// line#=../rle.cpp:80
	7'h61 :
		TR_169 = TR_108 ;
	7'h62 :
		TR_169 = TR_108 ;
	7'h63 :
		TR_169 = TR_108 ;
	7'h64 :
		TR_169 = TR_108 ;
	7'h65 :
		TR_169 = TR_108 ;
	7'h66 :
		TR_169 = TR_108 ;
	7'h67 :
		TR_169 = TR_108 ;
	7'h68 :
		TR_169 = TR_108 ;
	7'h69 :
		TR_169 = TR_108 ;
	7'h6a :
		TR_169 = TR_108 ;
	7'h6b :
		TR_169 = TR_108 ;
	7'h6c :
		TR_169 = TR_108 ;
	7'h6d :
		TR_169 = TR_108 ;
	7'h6e :
		TR_169 = TR_108 ;
	7'h6f :
		TR_169 = TR_108 ;
	7'h70 :
		TR_169 = TR_108 ;
	7'h71 :
		TR_169 = TR_108 ;
	7'h72 :
		TR_169 = TR_108 ;
	7'h73 :
		TR_169 = TR_108 ;
	7'h74 :
		TR_169 = TR_108 ;
	7'h75 :
		TR_169 = TR_108 ;
	7'h76 :
		TR_169 = TR_108 ;
	7'h77 :
		TR_169 = TR_108 ;
	7'h78 :
		TR_169 = TR_108 ;
	7'h79 :
		TR_169 = TR_108 ;
	7'h7a :
		TR_169 = TR_108 ;
	7'h7b :
		TR_169 = TR_108 ;
	7'h7c :
		TR_169 = TR_108 ;
	7'h7d :
		TR_169 = TR_108 ;
	7'h7e :
		TR_169 = TR_108 ;
	7'h7f :
		TR_169 = TR_108 ;
	default :
		TR_169 = 9'hx ;
	endcase
always @ ( TR_169 or U_173 or sub8u_71ot or U_183 or RG_rl_177 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_96_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h60 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_96_t = ( ( { 9{ M_180 } } & RG_rl_177 )
		| ( { 9{ U_173 } } & TR_169 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_96_en = ( M_180 | RG_rl_96_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_96_en )
		RG_rl_96 <= RG_rl_96_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_109 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_168 = TR_109 ;
	7'h01 :
		TR_168 = TR_109 ;
	7'h02 :
		TR_168 = TR_109 ;
	7'h03 :
		TR_168 = TR_109 ;
	7'h04 :
		TR_168 = TR_109 ;
	7'h05 :
		TR_168 = TR_109 ;
	7'h06 :
		TR_168 = TR_109 ;
	7'h07 :
		TR_168 = TR_109 ;
	7'h08 :
		TR_168 = TR_109 ;
	7'h09 :
		TR_168 = TR_109 ;
	7'h0a :
		TR_168 = TR_109 ;
	7'h0b :
		TR_168 = TR_109 ;
	7'h0c :
		TR_168 = TR_109 ;
	7'h0d :
		TR_168 = TR_109 ;
	7'h0e :
		TR_168 = TR_109 ;
	7'h0f :
		TR_168 = TR_109 ;
	7'h10 :
		TR_168 = TR_109 ;
	7'h11 :
		TR_168 = TR_109 ;
	7'h12 :
		TR_168 = TR_109 ;
	7'h13 :
		TR_168 = TR_109 ;
	7'h14 :
		TR_168 = TR_109 ;
	7'h15 :
		TR_168 = TR_109 ;
	7'h16 :
		TR_168 = TR_109 ;
	7'h17 :
		TR_168 = TR_109 ;
	7'h18 :
		TR_168 = TR_109 ;
	7'h19 :
		TR_168 = TR_109 ;
	7'h1a :
		TR_168 = TR_109 ;
	7'h1b :
		TR_168 = TR_109 ;
	7'h1c :
		TR_168 = TR_109 ;
	7'h1d :
		TR_168 = TR_109 ;
	7'h1e :
		TR_168 = TR_109 ;
	7'h1f :
		TR_168 = TR_109 ;
	7'h20 :
		TR_168 = TR_109 ;
	7'h21 :
		TR_168 = TR_109 ;
	7'h22 :
		TR_168 = TR_109 ;
	7'h23 :
		TR_168 = TR_109 ;
	7'h24 :
		TR_168 = TR_109 ;
	7'h25 :
		TR_168 = TR_109 ;
	7'h26 :
		TR_168 = TR_109 ;
	7'h27 :
		TR_168 = TR_109 ;
	7'h28 :
		TR_168 = TR_109 ;
	7'h29 :
		TR_168 = TR_109 ;
	7'h2a :
		TR_168 = TR_109 ;
	7'h2b :
		TR_168 = TR_109 ;
	7'h2c :
		TR_168 = TR_109 ;
	7'h2d :
		TR_168 = TR_109 ;
	7'h2e :
		TR_168 = TR_109 ;
	7'h2f :
		TR_168 = TR_109 ;
	7'h30 :
		TR_168 = TR_109 ;
	7'h31 :
		TR_168 = TR_109 ;
	7'h32 :
		TR_168 = TR_109 ;
	7'h33 :
		TR_168 = TR_109 ;
	7'h34 :
		TR_168 = TR_109 ;
	7'h35 :
		TR_168 = TR_109 ;
	7'h36 :
		TR_168 = TR_109 ;
	7'h37 :
		TR_168 = TR_109 ;
	7'h38 :
		TR_168 = TR_109 ;
	7'h39 :
		TR_168 = TR_109 ;
	7'h3a :
		TR_168 = TR_109 ;
	7'h3b :
		TR_168 = TR_109 ;
	7'h3c :
		TR_168 = TR_109 ;
	7'h3d :
		TR_168 = TR_109 ;
	7'h3e :
		TR_168 = TR_109 ;
	7'h3f :
		TR_168 = TR_109 ;
	7'h40 :
		TR_168 = TR_109 ;
	7'h41 :
		TR_168 = TR_109 ;
	7'h42 :
		TR_168 = TR_109 ;
	7'h43 :
		TR_168 = TR_109 ;
	7'h44 :
		TR_168 = TR_109 ;
	7'h45 :
		TR_168 = TR_109 ;
	7'h46 :
		TR_168 = TR_109 ;
	7'h47 :
		TR_168 = TR_109 ;
	7'h48 :
		TR_168 = TR_109 ;
	7'h49 :
		TR_168 = TR_109 ;
	7'h4a :
		TR_168 = TR_109 ;
	7'h4b :
		TR_168 = TR_109 ;
	7'h4c :
		TR_168 = TR_109 ;
	7'h4d :
		TR_168 = TR_109 ;
	7'h4e :
		TR_168 = TR_109 ;
	7'h4f :
		TR_168 = TR_109 ;
	7'h50 :
		TR_168 = TR_109 ;
	7'h51 :
		TR_168 = TR_109 ;
	7'h52 :
		TR_168 = TR_109 ;
	7'h53 :
		TR_168 = TR_109 ;
	7'h54 :
		TR_168 = TR_109 ;
	7'h55 :
		TR_168 = TR_109 ;
	7'h56 :
		TR_168 = TR_109 ;
	7'h57 :
		TR_168 = TR_109 ;
	7'h58 :
		TR_168 = TR_109 ;
	7'h59 :
		TR_168 = TR_109 ;
	7'h5a :
		TR_168 = TR_109 ;
	7'h5b :
		TR_168 = TR_109 ;
	7'h5c :
		TR_168 = TR_109 ;
	7'h5d :
		TR_168 = TR_109 ;
	7'h5e :
		TR_168 = TR_109 ;
	7'h5f :
		TR_168 = TR_109 ;
	7'h60 :
		TR_168 = TR_109 ;
	7'h61 :
		TR_168 = 9'h000 ;	// line#=../rle.cpp:80
	7'h62 :
		TR_168 = TR_109 ;
	7'h63 :
		TR_168 = TR_109 ;
	7'h64 :
		TR_168 = TR_109 ;
	7'h65 :
		TR_168 = TR_109 ;
	7'h66 :
		TR_168 = TR_109 ;
	7'h67 :
		TR_168 = TR_109 ;
	7'h68 :
		TR_168 = TR_109 ;
	7'h69 :
		TR_168 = TR_109 ;
	7'h6a :
		TR_168 = TR_109 ;
	7'h6b :
		TR_168 = TR_109 ;
	7'h6c :
		TR_168 = TR_109 ;
	7'h6d :
		TR_168 = TR_109 ;
	7'h6e :
		TR_168 = TR_109 ;
	7'h6f :
		TR_168 = TR_109 ;
	7'h70 :
		TR_168 = TR_109 ;
	7'h71 :
		TR_168 = TR_109 ;
	7'h72 :
		TR_168 = TR_109 ;
	7'h73 :
		TR_168 = TR_109 ;
	7'h74 :
		TR_168 = TR_109 ;
	7'h75 :
		TR_168 = TR_109 ;
	7'h76 :
		TR_168 = TR_109 ;
	7'h77 :
		TR_168 = TR_109 ;
	7'h78 :
		TR_168 = TR_109 ;
	7'h79 :
		TR_168 = TR_109 ;
	7'h7a :
		TR_168 = TR_109 ;
	7'h7b :
		TR_168 = TR_109 ;
	7'h7c :
		TR_168 = TR_109 ;
	7'h7d :
		TR_168 = TR_109 ;
	7'h7e :
		TR_168 = TR_109 ;
	7'h7f :
		TR_168 = TR_109 ;
	default :
		TR_168 = 9'hx ;
	endcase
always @ ( TR_168 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_46 or 
	U_174 or RG_rl_177 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_97_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h61 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_97_t = ( ( { 9{ ST1_03d } } & RG_rl_177 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_46 )
		| ( { 9{ U_173 } } & TR_168 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_97_en = ( ST1_03d | U_174 | RG_rl_97_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_97_en )
		RG_rl_97 <= RG_rl_97_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_110 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_167 = TR_110 ;
	7'h01 :
		TR_167 = TR_110 ;
	7'h02 :
		TR_167 = TR_110 ;
	7'h03 :
		TR_167 = TR_110 ;
	7'h04 :
		TR_167 = TR_110 ;
	7'h05 :
		TR_167 = TR_110 ;
	7'h06 :
		TR_167 = TR_110 ;
	7'h07 :
		TR_167 = TR_110 ;
	7'h08 :
		TR_167 = TR_110 ;
	7'h09 :
		TR_167 = TR_110 ;
	7'h0a :
		TR_167 = TR_110 ;
	7'h0b :
		TR_167 = TR_110 ;
	7'h0c :
		TR_167 = TR_110 ;
	7'h0d :
		TR_167 = TR_110 ;
	7'h0e :
		TR_167 = TR_110 ;
	7'h0f :
		TR_167 = TR_110 ;
	7'h10 :
		TR_167 = TR_110 ;
	7'h11 :
		TR_167 = TR_110 ;
	7'h12 :
		TR_167 = TR_110 ;
	7'h13 :
		TR_167 = TR_110 ;
	7'h14 :
		TR_167 = TR_110 ;
	7'h15 :
		TR_167 = TR_110 ;
	7'h16 :
		TR_167 = TR_110 ;
	7'h17 :
		TR_167 = TR_110 ;
	7'h18 :
		TR_167 = TR_110 ;
	7'h19 :
		TR_167 = TR_110 ;
	7'h1a :
		TR_167 = TR_110 ;
	7'h1b :
		TR_167 = TR_110 ;
	7'h1c :
		TR_167 = TR_110 ;
	7'h1d :
		TR_167 = TR_110 ;
	7'h1e :
		TR_167 = TR_110 ;
	7'h1f :
		TR_167 = TR_110 ;
	7'h20 :
		TR_167 = TR_110 ;
	7'h21 :
		TR_167 = TR_110 ;
	7'h22 :
		TR_167 = TR_110 ;
	7'h23 :
		TR_167 = TR_110 ;
	7'h24 :
		TR_167 = TR_110 ;
	7'h25 :
		TR_167 = TR_110 ;
	7'h26 :
		TR_167 = TR_110 ;
	7'h27 :
		TR_167 = TR_110 ;
	7'h28 :
		TR_167 = TR_110 ;
	7'h29 :
		TR_167 = TR_110 ;
	7'h2a :
		TR_167 = TR_110 ;
	7'h2b :
		TR_167 = TR_110 ;
	7'h2c :
		TR_167 = TR_110 ;
	7'h2d :
		TR_167 = TR_110 ;
	7'h2e :
		TR_167 = TR_110 ;
	7'h2f :
		TR_167 = TR_110 ;
	7'h30 :
		TR_167 = TR_110 ;
	7'h31 :
		TR_167 = TR_110 ;
	7'h32 :
		TR_167 = TR_110 ;
	7'h33 :
		TR_167 = TR_110 ;
	7'h34 :
		TR_167 = TR_110 ;
	7'h35 :
		TR_167 = TR_110 ;
	7'h36 :
		TR_167 = TR_110 ;
	7'h37 :
		TR_167 = TR_110 ;
	7'h38 :
		TR_167 = TR_110 ;
	7'h39 :
		TR_167 = TR_110 ;
	7'h3a :
		TR_167 = TR_110 ;
	7'h3b :
		TR_167 = TR_110 ;
	7'h3c :
		TR_167 = TR_110 ;
	7'h3d :
		TR_167 = TR_110 ;
	7'h3e :
		TR_167 = TR_110 ;
	7'h3f :
		TR_167 = TR_110 ;
	7'h40 :
		TR_167 = TR_110 ;
	7'h41 :
		TR_167 = TR_110 ;
	7'h42 :
		TR_167 = TR_110 ;
	7'h43 :
		TR_167 = TR_110 ;
	7'h44 :
		TR_167 = TR_110 ;
	7'h45 :
		TR_167 = TR_110 ;
	7'h46 :
		TR_167 = TR_110 ;
	7'h47 :
		TR_167 = TR_110 ;
	7'h48 :
		TR_167 = TR_110 ;
	7'h49 :
		TR_167 = TR_110 ;
	7'h4a :
		TR_167 = TR_110 ;
	7'h4b :
		TR_167 = TR_110 ;
	7'h4c :
		TR_167 = TR_110 ;
	7'h4d :
		TR_167 = TR_110 ;
	7'h4e :
		TR_167 = TR_110 ;
	7'h4f :
		TR_167 = TR_110 ;
	7'h50 :
		TR_167 = TR_110 ;
	7'h51 :
		TR_167 = TR_110 ;
	7'h52 :
		TR_167 = TR_110 ;
	7'h53 :
		TR_167 = TR_110 ;
	7'h54 :
		TR_167 = TR_110 ;
	7'h55 :
		TR_167 = TR_110 ;
	7'h56 :
		TR_167 = TR_110 ;
	7'h57 :
		TR_167 = TR_110 ;
	7'h58 :
		TR_167 = TR_110 ;
	7'h59 :
		TR_167 = TR_110 ;
	7'h5a :
		TR_167 = TR_110 ;
	7'h5b :
		TR_167 = TR_110 ;
	7'h5c :
		TR_167 = TR_110 ;
	7'h5d :
		TR_167 = TR_110 ;
	7'h5e :
		TR_167 = TR_110 ;
	7'h5f :
		TR_167 = TR_110 ;
	7'h60 :
		TR_167 = TR_110 ;
	7'h61 :
		TR_167 = TR_110 ;
	7'h62 :
		TR_167 = 9'h000 ;	// line#=../rle.cpp:80
	7'h63 :
		TR_167 = TR_110 ;
	7'h64 :
		TR_167 = TR_110 ;
	7'h65 :
		TR_167 = TR_110 ;
	7'h66 :
		TR_167 = TR_110 ;
	7'h67 :
		TR_167 = TR_110 ;
	7'h68 :
		TR_167 = TR_110 ;
	7'h69 :
		TR_167 = TR_110 ;
	7'h6a :
		TR_167 = TR_110 ;
	7'h6b :
		TR_167 = TR_110 ;
	7'h6c :
		TR_167 = TR_110 ;
	7'h6d :
		TR_167 = TR_110 ;
	7'h6e :
		TR_167 = TR_110 ;
	7'h6f :
		TR_167 = TR_110 ;
	7'h70 :
		TR_167 = TR_110 ;
	7'h71 :
		TR_167 = TR_110 ;
	7'h72 :
		TR_167 = TR_110 ;
	7'h73 :
		TR_167 = TR_110 ;
	7'h74 :
		TR_167 = TR_110 ;
	7'h75 :
		TR_167 = TR_110 ;
	7'h76 :
		TR_167 = TR_110 ;
	7'h77 :
		TR_167 = TR_110 ;
	7'h78 :
		TR_167 = TR_110 ;
	7'h79 :
		TR_167 = TR_110 ;
	7'h7a :
		TR_167 = TR_110 ;
	7'h7b :
		TR_167 = TR_110 ;
	7'h7c :
		TR_167 = TR_110 ;
	7'h7d :
		TR_167 = TR_110 ;
	7'h7e :
		TR_167 = TR_110 ;
	7'h7f :
		TR_167 = TR_110 ;
	default :
		TR_167 = 9'hx ;
	endcase
always @ ( TR_167 or U_173 or sub8u_71ot or U_183 or RG_rl_178 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_98_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h62 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_98_t = ( ( { 9{ M_180 } } & RG_rl_178 )
		| ( { 9{ U_173 } } & TR_167 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_98_en = ( M_180 | RG_rl_98_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_98_en )
		RG_rl_98 <= RG_rl_98_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_111 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_166 = TR_111 ;
	7'h01 :
		TR_166 = TR_111 ;
	7'h02 :
		TR_166 = TR_111 ;
	7'h03 :
		TR_166 = TR_111 ;
	7'h04 :
		TR_166 = TR_111 ;
	7'h05 :
		TR_166 = TR_111 ;
	7'h06 :
		TR_166 = TR_111 ;
	7'h07 :
		TR_166 = TR_111 ;
	7'h08 :
		TR_166 = TR_111 ;
	7'h09 :
		TR_166 = TR_111 ;
	7'h0a :
		TR_166 = TR_111 ;
	7'h0b :
		TR_166 = TR_111 ;
	7'h0c :
		TR_166 = TR_111 ;
	7'h0d :
		TR_166 = TR_111 ;
	7'h0e :
		TR_166 = TR_111 ;
	7'h0f :
		TR_166 = TR_111 ;
	7'h10 :
		TR_166 = TR_111 ;
	7'h11 :
		TR_166 = TR_111 ;
	7'h12 :
		TR_166 = TR_111 ;
	7'h13 :
		TR_166 = TR_111 ;
	7'h14 :
		TR_166 = TR_111 ;
	7'h15 :
		TR_166 = TR_111 ;
	7'h16 :
		TR_166 = TR_111 ;
	7'h17 :
		TR_166 = TR_111 ;
	7'h18 :
		TR_166 = TR_111 ;
	7'h19 :
		TR_166 = TR_111 ;
	7'h1a :
		TR_166 = TR_111 ;
	7'h1b :
		TR_166 = TR_111 ;
	7'h1c :
		TR_166 = TR_111 ;
	7'h1d :
		TR_166 = TR_111 ;
	7'h1e :
		TR_166 = TR_111 ;
	7'h1f :
		TR_166 = TR_111 ;
	7'h20 :
		TR_166 = TR_111 ;
	7'h21 :
		TR_166 = TR_111 ;
	7'h22 :
		TR_166 = TR_111 ;
	7'h23 :
		TR_166 = TR_111 ;
	7'h24 :
		TR_166 = TR_111 ;
	7'h25 :
		TR_166 = TR_111 ;
	7'h26 :
		TR_166 = TR_111 ;
	7'h27 :
		TR_166 = TR_111 ;
	7'h28 :
		TR_166 = TR_111 ;
	7'h29 :
		TR_166 = TR_111 ;
	7'h2a :
		TR_166 = TR_111 ;
	7'h2b :
		TR_166 = TR_111 ;
	7'h2c :
		TR_166 = TR_111 ;
	7'h2d :
		TR_166 = TR_111 ;
	7'h2e :
		TR_166 = TR_111 ;
	7'h2f :
		TR_166 = TR_111 ;
	7'h30 :
		TR_166 = TR_111 ;
	7'h31 :
		TR_166 = TR_111 ;
	7'h32 :
		TR_166 = TR_111 ;
	7'h33 :
		TR_166 = TR_111 ;
	7'h34 :
		TR_166 = TR_111 ;
	7'h35 :
		TR_166 = TR_111 ;
	7'h36 :
		TR_166 = TR_111 ;
	7'h37 :
		TR_166 = TR_111 ;
	7'h38 :
		TR_166 = TR_111 ;
	7'h39 :
		TR_166 = TR_111 ;
	7'h3a :
		TR_166 = TR_111 ;
	7'h3b :
		TR_166 = TR_111 ;
	7'h3c :
		TR_166 = TR_111 ;
	7'h3d :
		TR_166 = TR_111 ;
	7'h3e :
		TR_166 = TR_111 ;
	7'h3f :
		TR_166 = TR_111 ;
	7'h40 :
		TR_166 = TR_111 ;
	7'h41 :
		TR_166 = TR_111 ;
	7'h42 :
		TR_166 = TR_111 ;
	7'h43 :
		TR_166 = TR_111 ;
	7'h44 :
		TR_166 = TR_111 ;
	7'h45 :
		TR_166 = TR_111 ;
	7'h46 :
		TR_166 = TR_111 ;
	7'h47 :
		TR_166 = TR_111 ;
	7'h48 :
		TR_166 = TR_111 ;
	7'h49 :
		TR_166 = TR_111 ;
	7'h4a :
		TR_166 = TR_111 ;
	7'h4b :
		TR_166 = TR_111 ;
	7'h4c :
		TR_166 = TR_111 ;
	7'h4d :
		TR_166 = TR_111 ;
	7'h4e :
		TR_166 = TR_111 ;
	7'h4f :
		TR_166 = TR_111 ;
	7'h50 :
		TR_166 = TR_111 ;
	7'h51 :
		TR_166 = TR_111 ;
	7'h52 :
		TR_166 = TR_111 ;
	7'h53 :
		TR_166 = TR_111 ;
	7'h54 :
		TR_166 = TR_111 ;
	7'h55 :
		TR_166 = TR_111 ;
	7'h56 :
		TR_166 = TR_111 ;
	7'h57 :
		TR_166 = TR_111 ;
	7'h58 :
		TR_166 = TR_111 ;
	7'h59 :
		TR_166 = TR_111 ;
	7'h5a :
		TR_166 = TR_111 ;
	7'h5b :
		TR_166 = TR_111 ;
	7'h5c :
		TR_166 = TR_111 ;
	7'h5d :
		TR_166 = TR_111 ;
	7'h5e :
		TR_166 = TR_111 ;
	7'h5f :
		TR_166 = TR_111 ;
	7'h60 :
		TR_166 = TR_111 ;
	7'h61 :
		TR_166 = TR_111 ;
	7'h62 :
		TR_166 = TR_111 ;
	7'h63 :
		TR_166 = 9'h000 ;	// line#=../rle.cpp:80
	7'h64 :
		TR_166 = TR_111 ;
	7'h65 :
		TR_166 = TR_111 ;
	7'h66 :
		TR_166 = TR_111 ;
	7'h67 :
		TR_166 = TR_111 ;
	7'h68 :
		TR_166 = TR_111 ;
	7'h69 :
		TR_166 = TR_111 ;
	7'h6a :
		TR_166 = TR_111 ;
	7'h6b :
		TR_166 = TR_111 ;
	7'h6c :
		TR_166 = TR_111 ;
	7'h6d :
		TR_166 = TR_111 ;
	7'h6e :
		TR_166 = TR_111 ;
	7'h6f :
		TR_166 = TR_111 ;
	7'h70 :
		TR_166 = TR_111 ;
	7'h71 :
		TR_166 = TR_111 ;
	7'h72 :
		TR_166 = TR_111 ;
	7'h73 :
		TR_166 = TR_111 ;
	7'h74 :
		TR_166 = TR_111 ;
	7'h75 :
		TR_166 = TR_111 ;
	7'h76 :
		TR_166 = TR_111 ;
	7'h77 :
		TR_166 = TR_111 ;
	7'h78 :
		TR_166 = TR_111 ;
	7'h79 :
		TR_166 = TR_111 ;
	7'h7a :
		TR_166 = TR_111 ;
	7'h7b :
		TR_166 = TR_111 ;
	7'h7c :
		TR_166 = TR_111 ;
	7'h7d :
		TR_166 = TR_111 ;
	7'h7e :
		TR_166 = TR_111 ;
	7'h7f :
		TR_166 = TR_111 ;
	default :
		TR_166 = 9'hx ;
	endcase
always @ ( TR_166 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_47 or 
	U_174 or RG_rl_178 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_99_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h63 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_99_t = ( ( { 9{ ST1_03d } } & RG_rl_178 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_47 )
		| ( { 9{ U_173 } } & TR_166 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_99_en = ( ST1_03d | U_174 | RG_rl_99_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_99_en )
		RG_rl_99 <= RG_rl_99_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_112 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_165 = TR_112 ;
	7'h01 :
		TR_165 = TR_112 ;
	7'h02 :
		TR_165 = TR_112 ;
	7'h03 :
		TR_165 = TR_112 ;
	7'h04 :
		TR_165 = TR_112 ;
	7'h05 :
		TR_165 = TR_112 ;
	7'h06 :
		TR_165 = TR_112 ;
	7'h07 :
		TR_165 = TR_112 ;
	7'h08 :
		TR_165 = TR_112 ;
	7'h09 :
		TR_165 = TR_112 ;
	7'h0a :
		TR_165 = TR_112 ;
	7'h0b :
		TR_165 = TR_112 ;
	7'h0c :
		TR_165 = TR_112 ;
	7'h0d :
		TR_165 = TR_112 ;
	7'h0e :
		TR_165 = TR_112 ;
	7'h0f :
		TR_165 = TR_112 ;
	7'h10 :
		TR_165 = TR_112 ;
	7'h11 :
		TR_165 = TR_112 ;
	7'h12 :
		TR_165 = TR_112 ;
	7'h13 :
		TR_165 = TR_112 ;
	7'h14 :
		TR_165 = TR_112 ;
	7'h15 :
		TR_165 = TR_112 ;
	7'h16 :
		TR_165 = TR_112 ;
	7'h17 :
		TR_165 = TR_112 ;
	7'h18 :
		TR_165 = TR_112 ;
	7'h19 :
		TR_165 = TR_112 ;
	7'h1a :
		TR_165 = TR_112 ;
	7'h1b :
		TR_165 = TR_112 ;
	7'h1c :
		TR_165 = TR_112 ;
	7'h1d :
		TR_165 = TR_112 ;
	7'h1e :
		TR_165 = TR_112 ;
	7'h1f :
		TR_165 = TR_112 ;
	7'h20 :
		TR_165 = TR_112 ;
	7'h21 :
		TR_165 = TR_112 ;
	7'h22 :
		TR_165 = TR_112 ;
	7'h23 :
		TR_165 = TR_112 ;
	7'h24 :
		TR_165 = TR_112 ;
	7'h25 :
		TR_165 = TR_112 ;
	7'h26 :
		TR_165 = TR_112 ;
	7'h27 :
		TR_165 = TR_112 ;
	7'h28 :
		TR_165 = TR_112 ;
	7'h29 :
		TR_165 = TR_112 ;
	7'h2a :
		TR_165 = TR_112 ;
	7'h2b :
		TR_165 = TR_112 ;
	7'h2c :
		TR_165 = TR_112 ;
	7'h2d :
		TR_165 = TR_112 ;
	7'h2e :
		TR_165 = TR_112 ;
	7'h2f :
		TR_165 = TR_112 ;
	7'h30 :
		TR_165 = TR_112 ;
	7'h31 :
		TR_165 = TR_112 ;
	7'h32 :
		TR_165 = TR_112 ;
	7'h33 :
		TR_165 = TR_112 ;
	7'h34 :
		TR_165 = TR_112 ;
	7'h35 :
		TR_165 = TR_112 ;
	7'h36 :
		TR_165 = TR_112 ;
	7'h37 :
		TR_165 = TR_112 ;
	7'h38 :
		TR_165 = TR_112 ;
	7'h39 :
		TR_165 = TR_112 ;
	7'h3a :
		TR_165 = TR_112 ;
	7'h3b :
		TR_165 = TR_112 ;
	7'h3c :
		TR_165 = TR_112 ;
	7'h3d :
		TR_165 = TR_112 ;
	7'h3e :
		TR_165 = TR_112 ;
	7'h3f :
		TR_165 = TR_112 ;
	7'h40 :
		TR_165 = TR_112 ;
	7'h41 :
		TR_165 = TR_112 ;
	7'h42 :
		TR_165 = TR_112 ;
	7'h43 :
		TR_165 = TR_112 ;
	7'h44 :
		TR_165 = TR_112 ;
	7'h45 :
		TR_165 = TR_112 ;
	7'h46 :
		TR_165 = TR_112 ;
	7'h47 :
		TR_165 = TR_112 ;
	7'h48 :
		TR_165 = TR_112 ;
	7'h49 :
		TR_165 = TR_112 ;
	7'h4a :
		TR_165 = TR_112 ;
	7'h4b :
		TR_165 = TR_112 ;
	7'h4c :
		TR_165 = TR_112 ;
	7'h4d :
		TR_165 = TR_112 ;
	7'h4e :
		TR_165 = TR_112 ;
	7'h4f :
		TR_165 = TR_112 ;
	7'h50 :
		TR_165 = TR_112 ;
	7'h51 :
		TR_165 = TR_112 ;
	7'h52 :
		TR_165 = TR_112 ;
	7'h53 :
		TR_165 = TR_112 ;
	7'h54 :
		TR_165 = TR_112 ;
	7'h55 :
		TR_165 = TR_112 ;
	7'h56 :
		TR_165 = TR_112 ;
	7'h57 :
		TR_165 = TR_112 ;
	7'h58 :
		TR_165 = TR_112 ;
	7'h59 :
		TR_165 = TR_112 ;
	7'h5a :
		TR_165 = TR_112 ;
	7'h5b :
		TR_165 = TR_112 ;
	7'h5c :
		TR_165 = TR_112 ;
	7'h5d :
		TR_165 = TR_112 ;
	7'h5e :
		TR_165 = TR_112 ;
	7'h5f :
		TR_165 = TR_112 ;
	7'h60 :
		TR_165 = TR_112 ;
	7'h61 :
		TR_165 = TR_112 ;
	7'h62 :
		TR_165 = TR_112 ;
	7'h63 :
		TR_165 = TR_112 ;
	7'h64 :
		TR_165 = 9'h000 ;	// line#=../rle.cpp:80
	7'h65 :
		TR_165 = TR_112 ;
	7'h66 :
		TR_165 = TR_112 ;
	7'h67 :
		TR_165 = TR_112 ;
	7'h68 :
		TR_165 = TR_112 ;
	7'h69 :
		TR_165 = TR_112 ;
	7'h6a :
		TR_165 = TR_112 ;
	7'h6b :
		TR_165 = TR_112 ;
	7'h6c :
		TR_165 = TR_112 ;
	7'h6d :
		TR_165 = TR_112 ;
	7'h6e :
		TR_165 = TR_112 ;
	7'h6f :
		TR_165 = TR_112 ;
	7'h70 :
		TR_165 = TR_112 ;
	7'h71 :
		TR_165 = TR_112 ;
	7'h72 :
		TR_165 = TR_112 ;
	7'h73 :
		TR_165 = TR_112 ;
	7'h74 :
		TR_165 = TR_112 ;
	7'h75 :
		TR_165 = TR_112 ;
	7'h76 :
		TR_165 = TR_112 ;
	7'h77 :
		TR_165 = TR_112 ;
	7'h78 :
		TR_165 = TR_112 ;
	7'h79 :
		TR_165 = TR_112 ;
	7'h7a :
		TR_165 = TR_112 ;
	7'h7b :
		TR_165 = TR_112 ;
	7'h7c :
		TR_165 = TR_112 ;
	7'h7d :
		TR_165 = TR_112 ;
	7'h7e :
		TR_165 = TR_112 ;
	7'h7f :
		TR_165 = TR_112 ;
	default :
		TR_165 = 9'hx ;
	endcase
always @ ( TR_165 or U_173 or sub8u_71ot or U_183 or RG_rl_179 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_100_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h64 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_100_t = ( ( { 9{ M_180 } } & RG_rl_179 )
		| ( { 9{ U_173 } } & TR_165 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_100_en = ( M_180 | RG_rl_100_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_100_en )
		RG_rl_100 <= RG_rl_100_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_113 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_164 = TR_113 ;
	7'h01 :
		TR_164 = TR_113 ;
	7'h02 :
		TR_164 = TR_113 ;
	7'h03 :
		TR_164 = TR_113 ;
	7'h04 :
		TR_164 = TR_113 ;
	7'h05 :
		TR_164 = TR_113 ;
	7'h06 :
		TR_164 = TR_113 ;
	7'h07 :
		TR_164 = TR_113 ;
	7'h08 :
		TR_164 = TR_113 ;
	7'h09 :
		TR_164 = TR_113 ;
	7'h0a :
		TR_164 = TR_113 ;
	7'h0b :
		TR_164 = TR_113 ;
	7'h0c :
		TR_164 = TR_113 ;
	7'h0d :
		TR_164 = TR_113 ;
	7'h0e :
		TR_164 = TR_113 ;
	7'h0f :
		TR_164 = TR_113 ;
	7'h10 :
		TR_164 = TR_113 ;
	7'h11 :
		TR_164 = TR_113 ;
	7'h12 :
		TR_164 = TR_113 ;
	7'h13 :
		TR_164 = TR_113 ;
	7'h14 :
		TR_164 = TR_113 ;
	7'h15 :
		TR_164 = TR_113 ;
	7'h16 :
		TR_164 = TR_113 ;
	7'h17 :
		TR_164 = TR_113 ;
	7'h18 :
		TR_164 = TR_113 ;
	7'h19 :
		TR_164 = TR_113 ;
	7'h1a :
		TR_164 = TR_113 ;
	7'h1b :
		TR_164 = TR_113 ;
	7'h1c :
		TR_164 = TR_113 ;
	7'h1d :
		TR_164 = TR_113 ;
	7'h1e :
		TR_164 = TR_113 ;
	7'h1f :
		TR_164 = TR_113 ;
	7'h20 :
		TR_164 = TR_113 ;
	7'h21 :
		TR_164 = TR_113 ;
	7'h22 :
		TR_164 = TR_113 ;
	7'h23 :
		TR_164 = TR_113 ;
	7'h24 :
		TR_164 = TR_113 ;
	7'h25 :
		TR_164 = TR_113 ;
	7'h26 :
		TR_164 = TR_113 ;
	7'h27 :
		TR_164 = TR_113 ;
	7'h28 :
		TR_164 = TR_113 ;
	7'h29 :
		TR_164 = TR_113 ;
	7'h2a :
		TR_164 = TR_113 ;
	7'h2b :
		TR_164 = TR_113 ;
	7'h2c :
		TR_164 = TR_113 ;
	7'h2d :
		TR_164 = TR_113 ;
	7'h2e :
		TR_164 = TR_113 ;
	7'h2f :
		TR_164 = TR_113 ;
	7'h30 :
		TR_164 = TR_113 ;
	7'h31 :
		TR_164 = TR_113 ;
	7'h32 :
		TR_164 = TR_113 ;
	7'h33 :
		TR_164 = TR_113 ;
	7'h34 :
		TR_164 = TR_113 ;
	7'h35 :
		TR_164 = TR_113 ;
	7'h36 :
		TR_164 = TR_113 ;
	7'h37 :
		TR_164 = TR_113 ;
	7'h38 :
		TR_164 = TR_113 ;
	7'h39 :
		TR_164 = TR_113 ;
	7'h3a :
		TR_164 = TR_113 ;
	7'h3b :
		TR_164 = TR_113 ;
	7'h3c :
		TR_164 = TR_113 ;
	7'h3d :
		TR_164 = TR_113 ;
	7'h3e :
		TR_164 = TR_113 ;
	7'h3f :
		TR_164 = TR_113 ;
	7'h40 :
		TR_164 = TR_113 ;
	7'h41 :
		TR_164 = TR_113 ;
	7'h42 :
		TR_164 = TR_113 ;
	7'h43 :
		TR_164 = TR_113 ;
	7'h44 :
		TR_164 = TR_113 ;
	7'h45 :
		TR_164 = TR_113 ;
	7'h46 :
		TR_164 = TR_113 ;
	7'h47 :
		TR_164 = TR_113 ;
	7'h48 :
		TR_164 = TR_113 ;
	7'h49 :
		TR_164 = TR_113 ;
	7'h4a :
		TR_164 = TR_113 ;
	7'h4b :
		TR_164 = TR_113 ;
	7'h4c :
		TR_164 = TR_113 ;
	7'h4d :
		TR_164 = TR_113 ;
	7'h4e :
		TR_164 = TR_113 ;
	7'h4f :
		TR_164 = TR_113 ;
	7'h50 :
		TR_164 = TR_113 ;
	7'h51 :
		TR_164 = TR_113 ;
	7'h52 :
		TR_164 = TR_113 ;
	7'h53 :
		TR_164 = TR_113 ;
	7'h54 :
		TR_164 = TR_113 ;
	7'h55 :
		TR_164 = TR_113 ;
	7'h56 :
		TR_164 = TR_113 ;
	7'h57 :
		TR_164 = TR_113 ;
	7'h58 :
		TR_164 = TR_113 ;
	7'h59 :
		TR_164 = TR_113 ;
	7'h5a :
		TR_164 = TR_113 ;
	7'h5b :
		TR_164 = TR_113 ;
	7'h5c :
		TR_164 = TR_113 ;
	7'h5d :
		TR_164 = TR_113 ;
	7'h5e :
		TR_164 = TR_113 ;
	7'h5f :
		TR_164 = TR_113 ;
	7'h60 :
		TR_164 = TR_113 ;
	7'h61 :
		TR_164 = TR_113 ;
	7'h62 :
		TR_164 = TR_113 ;
	7'h63 :
		TR_164 = TR_113 ;
	7'h64 :
		TR_164 = TR_113 ;
	7'h65 :
		TR_164 = 9'h000 ;	// line#=../rle.cpp:80
	7'h66 :
		TR_164 = TR_113 ;
	7'h67 :
		TR_164 = TR_113 ;
	7'h68 :
		TR_164 = TR_113 ;
	7'h69 :
		TR_164 = TR_113 ;
	7'h6a :
		TR_164 = TR_113 ;
	7'h6b :
		TR_164 = TR_113 ;
	7'h6c :
		TR_164 = TR_113 ;
	7'h6d :
		TR_164 = TR_113 ;
	7'h6e :
		TR_164 = TR_113 ;
	7'h6f :
		TR_164 = TR_113 ;
	7'h70 :
		TR_164 = TR_113 ;
	7'h71 :
		TR_164 = TR_113 ;
	7'h72 :
		TR_164 = TR_113 ;
	7'h73 :
		TR_164 = TR_113 ;
	7'h74 :
		TR_164 = TR_113 ;
	7'h75 :
		TR_164 = TR_113 ;
	7'h76 :
		TR_164 = TR_113 ;
	7'h77 :
		TR_164 = TR_113 ;
	7'h78 :
		TR_164 = TR_113 ;
	7'h79 :
		TR_164 = TR_113 ;
	7'h7a :
		TR_164 = TR_113 ;
	7'h7b :
		TR_164 = TR_113 ;
	7'h7c :
		TR_164 = TR_113 ;
	7'h7d :
		TR_164 = TR_113 ;
	7'h7e :
		TR_164 = TR_113 ;
	7'h7f :
		TR_164 = TR_113 ;
	default :
		TR_164 = 9'hx ;
	endcase
always @ ( TR_164 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_48 or 
	U_174 or RG_rl_179 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_101_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h65 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_101_t = ( ( { 9{ ST1_03d } } & RG_rl_179 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_48 )
		| ( { 9{ U_173 } } & TR_164 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_101_en = ( ST1_03d | U_174 | RG_rl_101_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_101_en )
		RG_rl_101 <= RG_rl_101_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_114 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_163 = TR_114 ;
	7'h01 :
		TR_163 = TR_114 ;
	7'h02 :
		TR_163 = TR_114 ;
	7'h03 :
		TR_163 = TR_114 ;
	7'h04 :
		TR_163 = TR_114 ;
	7'h05 :
		TR_163 = TR_114 ;
	7'h06 :
		TR_163 = TR_114 ;
	7'h07 :
		TR_163 = TR_114 ;
	7'h08 :
		TR_163 = TR_114 ;
	7'h09 :
		TR_163 = TR_114 ;
	7'h0a :
		TR_163 = TR_114 ;
	7'h0b :
		TR_163 = TR_114 ;
	7'h0c :
		TR_163 = TR_114 ;
	7'h0d :
		TR_163 = TR_114 ;
	7'h0e :
		TR_163 = TR_114 ;
	7'h0f :
		TR_163 = TR_114 ;
	7'h10 :
		TR_163 = TR_114 ;
	7'h11 :
		TR_163 = TR_114 ;
	7'h12 :
		TR_163 = TR_114 ;
	7'h13 :
		TR_163 = TR_114 ;
	7'h14 :
		TR_163 = TR_114 ;
	7'h15 :
		TR_163 = TR_114 ;
	7'h16 :
		TR_163 = TR_114 ;
	7'h17 :
		TR_163 = TR_114 ;
	7'h18 :
		TR_163 = TR_114 ;
	7'h19 :
		TR_163 = TR_114 ;
	7'h1a :
		TR_163 = TR_114 ;
	7'h1b :
		TR_163 = TR_114 ;
	7'h1c :
		TR_163 = TR_114 ;
	7'h1d :
		TR_163 = TR_114 ;
	7'h1e :
		TR_163 = TR_114 ;
	7'h1f :
		TR_163 = TR_114 ;
	7'h20 :
		TR_163 = TR_114 ;
	7'h21 :
		TR_163 = TR_114 ;
	7'h22 :
		TR_163 = TR_114 ;
	7'h23 :
		TR_163 = TR_114 ;
	7'h24 :
		TR_163 = TR_114 ;
	7'h25 :
		TR_163 = TR_114 ;
	7'h26 :
		TR_163 = TR_114 ;
	7'h27 :
		TR_163 = TR_114 ;
	7'h28 :
		TR_163 = TR_114 ;
	7'h29 :
		TR_163 = TR_114 ;
	7'h2a :
		TR_163 = TR_114 ;
	7'h2b :
		TR_163 = TR_114 ;
	7'h2c :
		TR_163 = TR_114 ;
	7'h2d :
		TR_163 = TR_114 ;
	7'h2e :
		TR_163 = TR_114 ;
	7'h2f :
		TR_163 = TR_114 ;
	7'h30 :
		TR_163 = TR_114 ;
	7'h31 :
		TR_163 = TR_114 ;
	7'h32 :
		TR_163 = TR_114 ;
	7'h33 :
		TR_163 = TR_114 ;
	7'h34 :
		TR_163 = TR_114 ;
	7'h35 :
		TR_163 = TR_114 ;
	7'h36 :
		TR_163 = TR_114 ;
	7'h37 :
		TR_163 = TR_114 ;
	7'h38 :
		TR_163 = TR_114 ;
	7'h39 :
		TR_163 = TR_114 ;
	7'h3a :
		TR_163 = TR_114 ;
	7'h3b :
		TR_163 = TR_114 ;
	7'h3c :
		TR_163 = TR_114 ;
	7'h3d :
		TR_163 = TR_114 ;
	7'h3e :
		TR_163 = TR_114 ;
	7'h3f :
		TR_163 = TR_114 ;
	7'h40 :
		TR_163 = TR_114 ;
	7'h41 :
		TR_163 = TR_114 ;
	7'h42 :
		TR_163 = TR_114 ;
	7'h43 :
		TR_163 = TR_114 ;
	7'h44 :
		TR_163 = TR_114 ;
	7'h45 :
		TR_163 = TR_114 ;
	7'h46 :
		TR_163 = TR_114 ;
	7'h47 :
		TR_163 = TR_114 ;
	7'h48 :
		TR_163 = TR_114 ;
	7'h49 :
		TR_163 = TR_114 ;
	7'h4a :
		TR_163 = TR_114 ;
	7'h4b :
		TR_163 = TR_114 ;
	7'h4c :
		TR_163 = TR_114 ;
	7'h4d :
		TR_163 = TR_114 ;
	7'h4e :
		TR_163 = TR_114 ;
	7'h4f :
		TR_163 = TR_114 ;
	7'h50 :
		TR_163 = TR_114 ;
	7'h51 :
		TR_163 = TR_114 ;
	7'h52 :
		TR_163 = TR_114 ;
	7'h53 :
		TR_163 = TR_114 ;
	7'h54 :
		TR_163 = TR_114 ;
	7'h55 :
		TR_163 = TR_114 ;
	7'h56 :
		TR_163 = TR_114 ;
	7'h57 :
		TR_163 = TR_114 ;
	7'h58 :
		TR_163 = TR_114 ;
	7'h59 :
		TR_163 = TR_114 ;
	7'h5a :
		TR_163 = TR_114 ;
	7'h5b :
		TR_163 = TR_114 ;
	7'h5c :
		TR_163 = TR_114 ;
	7'h5d :
		TR_163 = TR_114 ;
	7'h5e :
		TR_163 = TR_114 ;
	7'h5f :
		TR_163 = TR_114 ;
	7'h60 :
		TR_163 = TR_114 ;
	7'h61 :
		TR_163 = TR_114 ;
	7'h62 :
		TR_163 = TR_114 ;
	7'h63 :
		TR_163 = TR_114 ;
	7'h64 :
		TR_163 = TR_114 ;
	7'h65 :
		TR_163 = TR_114 ;
	7'h66 :
		TR_163 = 9'h000 ;	// line#=../rle.cpp:80
	7'h67 :
		TR_163 = TR_114 ;
	7'h68 :
		TR_163 = TR_114 ;
	7'h69 :
		TR_163 = TR_114 ;
	7'h6a :
		TR_163 = TR_114 ;
	7'h6b :
		TR_163 = TR_114 ;
	7'h6c :
		TR_163 = TR_114 ;
	7'h6d :
		TR_163 = TR_114 ;
	7'h6e :
		TR_163 = TR_114 ;
	7'h6f :
		TR_163 = TR_114 ;
	7'h70 :
		TR_163 = TR_114 ;
	7'h71 :
		TR_163 = TR_114 ;
	7'h72 :
		TR_163 = TR_114 ;
	7'h73 :
		TR_163 = TR_114 ;
	7'h74 :
		TR_163 = TR_114 ;
	7'h75 :
		TR_163 = TR_114 ;
	7'h76 :
		TR_163 = TR_114 ;
	7'h77 :
		TR_163 = TR_114 ;
	7'h78 :
		TR_163 = TR_114 ;
	7'h79 :
		TR_163 = TR_114 ;
	7'h7a :
		TR_163 = TR_114 ;
	7'h7b :
		TR_163 = TR_114 ;
	7'h7c :
		TR_163 = TR_114 ;
	7'h7d :
		TR_163 = TR_114 ;
	7'h7e :
		TR_163 = TR_114 ;
	7'h7f :
		TR_163 = TR_114 ;
	default :
		TR_163 = 9'hx ;
	endcase
always @ ( TR_163 or U_173 or sub8u_71ot or U_183 or RG_rl_180 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_102_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h66 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_102_t = ( ( { 9{ M_180 } } & RG_rl_180 )
		| ( { 9{ U_173 } } & TR_163 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_102_en = ( M_180 | RG_rl_102_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_102_en )
		RG_rl_102 <= RG_rl_102_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_115 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_162 = TR_115 ;
	7'h01 :
		TR_162 = TR_115 ;
	7'h02 :
		TR_162 = TR_115 ;
	7'h03 :
		TR_162 = TR_115 ;
	7'h04 :
		TR_162 = TR_115 ;
	7'h05 :
		TR_162 = TR_115 ;
	7'h06 :
		TR_162 = TR_115 ;
	7'h07 :
		TR_162 = TR_115 ;
	7'h08 :
		TR_162 = TR_115 ;
	7'h09 :
		TR_162 = TR_115 ;
	7'h0a :
		TR_162 = TR_115 ;
	7'h0b :
		TR_162 = TR_115 ;
	7'h0c :
		TR_162 = TR_115 ;
	7'h0d :
		TR_162 = TR_115 ;
	7'h0e :
		TR_162 = TR_115 ;
	7'h0f :
		TR_162 = TR_115 ;
	7'h10 :
		TR_162 = TR_115 ;
	7'h11 :
		TR_162 = TR_115 ;
	7'h12 :
		TR_162 = TR_115 ;
	7'h13 :
		TR_162 = TR_115 ;
	7'h14 :
		TR_162 = TR_115 ;
	7'h15 :
		TR_162 = TR_115 ;
	7'h16 :
		TR_162 = TR_115 ;
	7'h17 :
		TR_162 = TR_115 ;
	7'h18 :
		TR_162 = TR_115 ;
	7'h19 :
		TR_162 = TR_115 ;
	7'h1a :
		TR_162 = TR_115 ;
	7'h1b :
		TR_162 = TR_115 ;
	7'h1c :
		TR_162 = TR_115 ;
	7'h1d :
		TR_162 = TR_115 ;
	7'h1e :
		TR_162 = TR_115 ;
	7'h1f :
		TR_162 = TR_115 ;
	7'h20 :
		TR_162 = TR_115 ;
	7'h21 :
		TR_162 = TR_115 ;
	7'h22 :
		TR_162 = TR_115 ;
	7'h23 :
		TR_162 = TR_115 ;
	7'h24 :
		TR_162 = TR_115 ;
	7'h25 :
		TR_162 = TR_115 ;
	7'h26 :
		TR_162 = TR_115 ;
	7'h27 :
		TR_162 = TR_115 ;
	7'h28 :
		TR_162 = TR_115 ;
	7'h29 :
		TR_162 = TR_115 ;
	7'h2a :
		TR_162 = TR_115 ;
	7'h2b :
		TR_162 = TR_115 ;
	7'h2c :
		TR_162 = TR_115 ;
	7'h2d :
		TR_162 = TR_115 ;
	7'h2e :
		TR_162 = TR_115 ;
	7'h2f :
		TR_162 = TR_115 ;
	7'h30 :
		TR_162 = TR_115 ;
	7'h31 :
		TR_162 = TR_115 ;
	7'h32 :
		TR_162 = TR_115 ;
	7'h33 :
		TR_162 = TR_115 ;
	7'h34 :
		TR_162 = TR_115 ;
	7'h35 :
		TR_162 = TR_115 ;
	7'h36 :
		TR_162 = TR_115 ;
	7'h37 :
		TR_162 = TR_115 ;
	7'h38 :
		TR_162 = TR_115 ;
	7'h39 :
		TR_162 = TR_115 ;
	7'h3a :
		TR_162 = TR_115 ;
	7'h3b :
		TR_162 = TR_115 ;
	7'h3c :
		TR_162 = TR_115 ;
	7'h3d :
		TR_162 = TR_115 ;
	7'h3e :
		TR_162 = TR_115 ;
	7'h3f :
		TR_162 = TR_115 ;
	7'h40 :
		TR_162 = TR_115 ;
	7'h41 :
		TR_162 = TR_115 ;
	7'h42 :
		TR_162 = TR_115 ;
	7'h43 :
		TR_162 = TR_115 ;
	7'h44 :
		TR_162 = TR_115 ;
	7'h45 :
		TR_162 = TR_115 ;
	7'h46 :
		TR_162 = TR_115 ;
	7'h47 :
		TR_162 = TR_115 ;
	7'h48 :
		TR_162 = TR_115 ;
	7'h49 :
		TR_162 = TR_115 ;
	7'h4a :
		TR_162 = TR_115 ;
	7'h4b :
		TR_162 = TR_115 ;
	7'h4c :
		TR_162 = TR_115 ;
	7'h4d :
		TR_162 = TR_115 ;
	7'h4e :
		TR_162 = TR_115 ;
	7'h4f :
		TR_162 = TR_115 ;
	7'h50 :
		TR_162 = TR_115 ;
	7'h51 :
		TR_162 = TR_115 ;
	7'h52 :
		TR_162 = TR_115 ;
	7'h53 :
		TR_162 = TR_115 ;
	7'h54 :
		TR_162 = TR_115 ;
	7'h55 :
		TR_162 = TR_115 ;
	7'h56 :
		TR_162 = TR_115 ;
	7'h57 :
		TR_162 = TR_115 ;
	7'h58 :
		TR_162 = TR_115 ;
	7'h59 :
		TR_162 = TR_115 ;
	7'h5a :
		TR_162 = TR_115 ;
	7'h5b :
		TR_162 = TR_115 ;
	7'h5c :
		TR_162 = TR_115 ;
	7'h5d :
		TR_162 = TR_115 ;
	7'h5e :
		TR_162 = TR_115 ;
	7'h5f :
		TR_162 = TR_115 ;
	7'h60 :
		TR_162 = TR_115 ;
	7'h61 :
		TR_162 = TR_115 ;
	7'h62 :
		TR_162 = TR_115 ;
	7'h63 :
		TR_162 = TR_115 ;
	7'h64 :
		TR_162 = TR_115 ;
	7'h65 :
		TR_162 = TR_115 ;
	7'h66 :
		TR_162 = TR_115 ;
	7'h67 :
		TR_162 = 9'h000 ;	// line#=../rle.cpp:80
	7'h68 :
		TR_162 = TR_115 ;
	7'h69 :
		TR_162 = TR_115 ;
	7'h6a :
		TR_162 = TR_115 ;
	7'h6b :
		TR_162 = TR_115 ;
	7'h6c :
		TR_162 = TR_115 ;
	7'h6d :
		TR_162 = TR_115 ;
	7'h6e :
		TR_162 = TR_115 ;
	7'h6f :
		TR_162 = TR_115 ;
	7'h70 :
		TR_162 = TR_115 ;
	7'h71 :
		TR_162 = TR_115 ;
	7'h72 :
		TR_162 = TR_115 ;
	7'h73 :
		TR_162 = TR_115 ;
	7'h74 :
		TR_162 = TR_115 ;
	7'h75 :
		TR_162 = TR_115 ;
	7'h76 :
		TR_162 = TR_115 ;
	7'h77 :
		TR_162 = TR_115 ;
	7'h78 :
		TR_162 = TR_115 ;
	7'h79 :
		TR_162 = TR_115 ;
	7'h7a :
		TR_162 = TR_115 ;
	7'h7b :
		TR_162 = TR_115 ;
	7'h7c :
		TR_162 = TR_115 ;
	7'h7d :
		TR_162 = TR_115 ;
	7'h7e :
		TR_162 = TR_115 ;
	7'h7f :
		TR_162 = TR_115 ;
	default :
		TR_162 = 9'hx ;
	endcase
always @ ( TR_162 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_49 or 
	U_174 or RG_rl_180 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_103_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h67 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_103_t = ( ( { 9{ ST1_03d } } & RG_rl_180 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_49 )
		| ( { 9{ U_173 } } & TR_162 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_103_en = ( ST1_03d | U_174 | RG_rl_103_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_103_en )
		RG_rl_103 <= RG_rl_103_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_116 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_161 = TR_116 ;
	7'h01 :
		TR_161 = TR_116 ;
	7'h02 :
		TR_161 = TR_116 ;
	7'h03 :
		TR_161 = TR_116 ;
	7'h04 :
		TR_161 = TR_116 ;
	7'h05 :
		TR_161 = TR_116 ;
	7'h06 :
		TR_161 = TR_116 ;
	7'h07 :
		TR_161 = TR_116 ;
	7'h08 :
		TR_161 = TR_116 ;
	7'h09 :
		TR_161 = TR_116 ;
	7'h0a :
		TR_161 = TR_116 ;
	7'h0b :
		TR_161 = TR_116 ;
	7'h0c :
		TR_161 = TR_116 ;
	7'h0d :
		TR_161 = TR_116 ;
	7'h0e :
		TR_161 = TR_116 ;
	7'h0f :
		TR_161 = TR_116 ;
	7'h10 :
		TR_161 = TR_116 ;
	7'h11 :
		TR_161 = TR_116 ;
	7'h12 :
		TR_161 = TR_116 ;
	7'h13 :
		TR_161 = TR_116 ;
	7'h14 :
		TR_161 = TR_116 ;
	7'h15 :
		TR_161 = TR_116 ;
	7'h16 :
		TR_161 = TR_116 ;
	7'h17 :
		TR_161 = TR_116 ;
	7'h18 :
		TR_161 = TR_116 ;
	7'h19 :
		TR_161 = TR_116 ;
	7'h1a :
		TR_161 = TR_116 ;
	7'h1b :
		TR_161 = TR_116 ;
	7'h1c :
		TR_161 = TR_116 ;
	7'h1d :
		TR_161 = TR_116 ;
	7'h1e :
		TR_161 = TR_116 ;
	7'h1f :
		TR_161 = TR_116 ;
	7'h20 :
		TR_161 = TR_116 ;
	7'h21 :
		TR_161 = TR_116 ;
	7'h22 :
		TR_161 = TR_116 ;
	7'h23 :
		TR_161 = TR_116 ;
	7'h24 :
		TR_161 = TR_116 ;
	7'h25 :
		TR_161 = TR_116 ;
	7'h26 :
		TR_161 = TR_116 ;
	7'h27 :
		TR_161 = TR_116 ;
	7'h28 :
		TR_161 = TR_116 ;
	7'h29 :
		TR_161 = TR_116 ;
	7'h2a :
		TR_161 = TR_116 ;
	7'h2b :
		TR_161 = TR_116 ;
	7'h2c :
		TR_161 = TR_116 ;
	7'h2d :
		TR_161 = TR_116 ;
	7'h2e :
		TR_161 = TR_116 ;
	7'h2f :
		TR_161 = TR_116 ;
	7'h30 :
		TR_161 = TR_116 ;
	7'h31 :
		TR_161 = TR_116 ;
	7'h32 :
		TR_161 = TR_116 ;
	7'h33 :
		TR_161 = TR_116 ;
	7'h34 :
		TR_161 = TR_116 ;
	7'h35 :
		TR_161 = TR_116 ;
	7'h36 :
		TR_161 = TR_116 ;
	7'h37 :
		TR_161 = TR_116 ;
	7'h38 :
		TR_161 = TR_116 ;
	7'h39 :
		TR_161 = TR_116 ;
	7'h3a :
		TR_161 = TR_116 ;
	7'h3b :
		TR_161 = TR_116 ;
	7'h3c :
		TR_161 = TR_116 ;
	7'h3d :
		TR_161 = TR_116 ;
	7'h3e :
		TR_161 = TR_116 ;
	7'h3f :
		TR_161 = TR_116 ;
	7'h40 :
		TR_161 = TR_116 ;
	7'h41 :
		TR_161 = TR_116 ;
	7'h42 :
		TR_161 = TR_116 ;
	7'h43 :
		TR_161 = TR_116 ;
	7'h44 :
		TR_161 = TR_116 ;
	7'h45 :
		TR_161 = TR_116 ;
	7'h46 :
		TR_161 = TR_116 ;
	7'h47 :
		TR_161 = TR_116 ;
	7'h48 :
		TR_161 = TR_116 ;
	7'h49 :
		TR_161 = TR_116 ;
	7'h4a :
		TR_161 = TR_116 ;
	7'h4b :
		TR_161 = TR_116 ;
	7'h4c :
		TR_161 = TR_116 ;
	7'h4d :
		TR_161 = TR_116 ;
	7'h4e :
		TR_161 = TR_116 ;
	7'h4f :
		TR_161 = TR_116 ;
	7'h50 :
		TR_161 = TR_116 ;
	7'h51 :
		TR_161 = TR_116 ;
	7'h52 :
		TR_161 = TR_116 ;
	7'h53 :
		TR_161 = TR_116 ;
	7'h54 :
		TR_161 = TR_116 ;
	7'h55 :
		TR_161 = TR_116 ;
	7'h56 :
		TR_161 = TR_116 ;
	7'h57 :
		TR_161 = TR_116 ;
	7'h58 :
		TR_161 = TR_116 ;
	7'h59 :
		TR_161 = TR_116 ;
	7'h5a :
		TR_161 = TR_116 ;
	7'h5b :
		TR_161 = TR_116 ;
	7'h5c :
		TR_161 = TR_116 ;
	7'h5d :
		TR_161 = TR_116 ;
	7'h5e :
		TR_161 = TR_116 ;
	7'h5f :
		TR_161 = TR_116 ;
	7'h60 :
		TR_161 = TR_116 ;
	7'h61 :
		TR_161 = TR_116 ;
	7'h62 :
		TR_161 = TR_116 ;
	7'h63 :
		TR_161 = TR_116 ;
	7'h64 :
		TR_161 = TR_116 ;
	7'h65 :
		TR_161 = TR_116 ;
	7'h66 :
		TR_161 = TR_116 ;
	7'h67 :
		TR_161 = TR_116 ;
	7'h68 :
		TR_161 = 9'h000 ;	// line#=../rle.cpp:80
	7'h69 :
		TR_161 = TR_116 ;
	7'h6a :
		TR_161 = TR_116 ;
	7'h6b :
		TR_161 = TR_116 ;
	7'h6c :
		TR_161 = TR_116 ;
	7'h6d :
		TR_161 = TR_116 ;
	7'h6e :
		TR_161 = TR_116 ;
	7'h6f :
		TR_161 = TR_116 ;
	7'h70 :
		TR_161 = TR_116 ;
	7'h71 :
		TR_161 = TR_116 ;
	7'h72 :
		TR_161 = TR_116 ;
	7'h73 :
		TR_161 = TR_116 ;
	7'h74 :
		TR_161 = TR_116 ;
	7'h75 :
		TR_161 = TR_116 ;
	7'h76 :
		TR_161 = TR_116 ;
	7'h77 :
		TR_161 = TR_116 ;
	7'h78 :
		TR_161 = TR_116 ;
	7'h79 :
		TR_161 = TR_116 ;
	7'h7a :
		TR_161 = TR_116 ;
	7'h7b :
		TR_161 = TR_116 ;
	7'h7c :
		TR_161 = TR_116 ;
	7'h7d :
		TR_161 = TR_116 ;
	7'h7e :
		TR_161 = TR_116 ;
	7'h7f :
		TR_161 = TR_116 ;
	default :
		TR_161 = 9'hx ;
	endcase
always @ ( TR_161 or U_173 or sub8u_71ot or U_183 or RG_rl_181 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_104_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h68 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_104_t = ( ( { 9{ M_180 } } & RG_rl_181 )
		| ( { 9{ U_173 } } & TR_161 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_104_en = ( M_180 | RG_rl_104_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_104_en )
		RG_rl_104 <= RG_rl_104_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_117 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_160 = TR_117 ;
	7'h01 :
		TR_160 = TR_117 ;
	7'h02 :
		TR_160 = TR_117 ;
	7'h03 :
		TR_160 = TR_117 ;
	7'h04 :
		TR_160 = TR_117 ;
	7'h05 :
		TR_160 = TR_117 ;
	7'h06 :
		TR_160 = TR_117 ;
	7'h07 :
		TR_160 = TR_117 ;
	7'h08 :
		TR_160 = TR_117 ;
	7'h09 :
		TR_160 = TR_117 ;
	7'h0a :
		TR_160 = TR_117 ;
	7'h0b :
		TR_160 = TR_117 ;
	7'h0c :
		TR_160 = TR_117 ;
	7'h0d :
		TR_160 = TR_117 ;
	7'h0e :
		TR_160 = TR_117 ;
	7'h0f :
		TR_160 = TR_117 ;
	7'h10 :
		TR_160 = TR_117 ;
	7'h11 :
		TR_160 = TR_117 ;
	7'h12 :
		TR_160 = TR_117 ;
	7'h13 :
		TR_160 = TR_117 ;
	7'h14 :
		TR_160 = TR_117 ;
	7'h15 :
		TR_160 = TR_117 ;
	7'h16 :
		TR_160 = TR_117 ;
	7'h17 :
		TR_160 = TR_117 ;
	7'h18 :
		TR_160 = TR_117 ;
	7'h19 :
		TR_160 = TR_117 ;
	7'h1a :
		TR_160 = TR_117 ;
	7'h1b :
		TR_160 = TR_117 ;
	7'h1c :
		TR_160 = TR_117 ;
	7'h1d :
		TR_160 = TR_117 ;
	7'h1e :
		TR_160 = TR_117 ;
	7'h1f :
		TR_160 = TR_117 ;
	7'h20 :
		TR_160 = TR_117 ;
	7'h21 :
		TR_160 = TR_117 ;
	7'h22 :
		TR_160 = TR_117 ;
	7'h23 :
		TR_160 = TR_117 ;
	7'h24 :
		TR_160 = TR_117 ;
	7'h25 :
		TR_160 = TR_117 ;
	7'h26 :
		TR_160 = TR_117 ;
	7'h27 :
		TR_160 = TR_117 ;
	7'h28 :
		TR_160 = TR_117 ;
	7'h29 :
		TR_160 = TR_117 ;
	7'h2a :
		TR_160 = TR_117 ;
	7'h2b :
		TR_160 = TR_117 ;
	7'h2c :
		TR_160 = TR_117 ;
	7'h2d :
		TR_160 = TR_117 ;
	7'h2e :
		TR_160 = TR_117 ;
	7'h2f :
		TR_160 = TR_117 ;
	7'h30 :
		TR_160 = TR_117 ;
	7'h31 :
		TR_160 = TR_117 ;
	7'h32 :
		TR_160 = TR_117 ;
	7'h33 :
		TR_160 = TR_117 ;
	7'h34 :
		TR_160 = TR_117 ;
	7'h35 :
		TR_160 = TR_117 ;
	7'h36 :
		TR_160 = TR_117 ;
	7'h37 :
		TR_160 = TR_117 ;
	7'h38 :
		TR_160 = TR_117 ;
	7'h39 :
		TR_160 = TR_117 ;
	7'h3a :
		TR_160 = TR_117 ;
	7'h3b :
		TR_160 = TR_117 ;
	7'h3c :
		TR_160 = TR_117 ;
	7'h3d :
		TR_160 = TR_117 ;
	7'h3e :
		TR_160 = TR_117 ;
	7'h3f :
		TR_160 = TR_117 ;
	7'h40 :
		TR_160 = TR_117 ;
	7'h41 :
		TR_160 = TR_117 ;
	7'h42 :
		TR_160 = TR_117 ;
	7'h43 :
		TR_160 = TR_117 ;
	7'h44 :
		TR_160 = TR_117 ;
	7'h45 :
		TR_160 = TR_117 ;
	7'h46 :
		TR_160 = TR_117 ;
	7'h47 :
		TR_160 = TR_117 ;
	7'h48 :
		TR_160 = TR_117 ;
	7'h49 :
		TR_160 = TR_117 ;
	7'h4a :
		TR_160 = TR_117 ;
	7'h4b :
		TR_160 = TR_117 ;
	7'h4c :
		TR_160 = TR_117 ;
	7'h4d :
		TR_160 = TR_117 ;
	7'h4e :
		TR_160 = TR_117 ;
	7'h4f :
		TR_160 = TR_117 ;
	7'h50 :
		TR_160 = TR_117 ;
	7'h51 :
		TR_160 = TR_117 ;
	7'h52 :
		TR_160 = TR_117 ;
	7'h53 :
		TR_160 = TR_117 ;
	7'h54 :
		TR_160 = TR_117 ;
	7'h55 :
		TR_160 = TR_117 ;
	7'h56 :
		TR_160 = TR_117 ;
	7'h57 :
		TR_160 = TR_117 ;
	7'h58 :
		TR_160 = TR_117 ;
	7'h59 :
		TR_160 = TR_117 ;
	7'h5a :
		TR_160 = TR_117 ;
	7'h5b :
		TR_160 = TR_117 ;
	7'h5c :
		TR_160 = TR_117 ;
	7'h5d :
		TR_160 = TR_117 ;
	7'h5e :
		TR_160 = TR_117 ;
	7'h5f :
		TR_160 = TR_117 ;
	7'h60 :
		TR_160 = TR_117 ;
	7'h61 :
		TR_160 = TR_117 ;
	7'h62 :
		TR_160 = TR_117 ;
	7'h63 :
		TR_160 = TR_117 ;
	7'h64 :
		TR_160 = TR_117 ;
	7'h65 :
		TR_160 = TR_117 ;
	7'h66 :
		TR_160 = TR_117 ;
	7'h67 :
		TR_160 = TR_117 ;
	7'h68 :
		TR_160 = TR_117 ;
	7'h69 :
		TR_160 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6a :
		TR_160 = TR_117 ;
	7'h6b :
		TR_160 = TR_117 ;
	7'h6c :
		TR_160 = TR_117 ;
	7'h6d :
		TR_160 = TR_117 ;
	7'h6e :
		TR_160 = TR_117 ;
	7'h6f :
		TR_160 = TR_117 ;
	7'h70 :
		TR_160 = TR_117 ;
	7'h71 :
		TR_160 = TR_117 ;
	7'h72 :
		TR_160 = TR_117 ;
	7'h73 :
		TR_160 = TR_117 ;
	7'h74 :
		TR_160 = TR_117 ;
	7'h75 :
		TR_160 = TR_117 ;
	7'h76 :
		TR_160 = TR_117 ;
	7'h77 :
		TR_160 = TR_117 ;
	7'h78 :
		TR_160 = TR_117 ;
	7'h79 :
		TR_160 = TR_117 ;
	7'h7a :
		TR_160 = TR_117 ;
	7'h7b :
		TR_160 = TR_117 ;
	7'h7c :
		TR_160 = TR_117 ;
	7'h7d :
		TR_160 = TR_117 ;
	7'h7e :
		TR_160 = TR_117 ;
	7'h7f :
		TR_160 = TR_117 ;
	default :
		TR_160 = 9'hx ;
	endcase
always @ ( TR_160 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_50 or 
	U_174 or RG_rl_181 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_105_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h69 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_105_t = ( ( { 9{ ST1_03d } } & RG_rl_181 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_50 )
		| ( { 9{ U_173 } } & TR_160 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_105_en = ( ST1_03d | U_174 | RG_rl_105_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_105_en )
		RG_rl_105 <= RG_rl_105_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_118 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_159 = TR_118 ;
	7'h01 :
		TR_159 = TR_118 ;
	7'h02 :
		TR_159 = TR_118 ;
	7'h03 :
		TR_159 = TR_118 ;
	7'h04 :
		TR_159 = TR_118 ;
	7'h05 :
		TR_159 = TR_118 ;
	7'h06 :
		TR_159 = TR_118 ;
	7'h07 :
		TR_159 = TR_118 ;
	7'h08 :
		TR_159 = TR_118 ;
	7'h09 :
		TR_159 = TR_118 ;
	7'h0a :
		TR_159 = TR_118 ;
	7'h0b :
		TR_159 = TR_118 ;
	7'h0c :
		TR_159 = TR_118 ;
	7'h0d :
		TR_159 = TR_118 ;
	7'h0e :
		TR_159 = TR_118 ;
	7'h0f :
		TR_159 = TR_118 ;
	7'h10 :
		TR_159 = TR_118 ;
	7'h11 :
		TR_159 = TR_118 ;
	7'h12 :
		TR_159 = TR_118 ;
	7'h13 :
		TR_159 = TR_118 ;
	7'h14 :
		TR_159 = TR_118 ;
	7'h15 :
		TR_159 = TR_118 ;
	7'h16 :
		TR_159 = TR_118 ;
	7'h17 :
		TR_159 = TR_118 ;
	7'h18 :
		TR_159 = TR_118 ;
	7'h19 :
		TR_159 = TR_118 ;
	7'h1a :
		TR_159 = TR_118 ;
	7'h1b :
		TR_159 = TR_118 ;
	7'h1c :
		TR_159 = TR_118 ;
	7'h1d :
		TR_159 = TR_118 ;
	7'h1e :
		TR_159 = TR_118 ;
	7'h1f :
		TR_159 = TR_118 ;
	7'h20 :
		TR_159 = TR_118 ;
	7'h21 :
		TR_159 = TR_118 ;
	7'h22 :
		TR_159 = TR_118 ;
	7'h23 :
		TR_159 = TR_118 ;
	7'h24 :
		TR_159 = TR_118 ;
	7'h25 :
		TR_159 = TR_118 ;
	7'h26 :
		TR_159 = TR_118 ;
	7'h27 :
		TR_159 = TR_118 ;
	7'h28 :
		TR_159 = TR_118 ;
	7'h29 :
		TR_159 = TR_118 ;
	7'h2a :
		TR_159 = TR_118 ;
	7'h2b :
		TR_159 = TR_118 ;
	7'h2c :
		TR_159 = TR_118 ;
	7'h2d :
		TR_159 = TR_118 ;
	7'h2e :
		TR_159 = TR_118 ;
	7'h2f :
		TR_159 = TR_118 ;
	7'h30 :
		TR_159 = TR_118 ;
	7'h31 :
		TR_159 = TR_118 ;
	7'h32 :
		TR_159 = TR_118 ;
	7'h33 :
		TR_159 = TR_118 ;
	7'h34 :
		TR_159 = TR_118 ;
	7'h35 :
		TR_159 = TR_118 ;
	7'h36 :
		TR_159 = TR_118 ;
	7'h37 :
		TR_159 = TR_118 ;
	7'h38 :
		TR_159 = TR_118 ;
	7'h39 :
		TR_159 = TR_118 ;
	7'h3a :
		TR_159 = TR_118 ;
	7'h3b :
		TR_159 = TR_118 ;
	7'h3c :
		TR_159 = TR_118 ;
	7'h3d :
		TR_159 = TR_118 ;
	7'h3e :
		TR_159 = TR_118 ;
	7'h3f :
		TR_159 = TR_118 ;
	7'h40 :
		TR_159 = TR_118 ;
	7'h41 :
		TR_159 = TR_118 ;
	7'h42 :
		TR_159 = TR_118 ;
	7'h43 :
		TR_159 = TR_118 ;
	7'h44 :
		TR_159 = TR_118 ;
	7'h45 :
		TR_159 = TR_118 ;
	7'h46 :
		TR_159 = TR_118 ;
	7'h47 :
		TR_159 = TR_118 ;
	7'h48 :
		TR_159 = TR_118 ;
	7'h49 :
		TR_159 = TR_118 ;
	7'h4a :
		TR_159 = TR_118 ;
	7'h4b :
		TR_159 = TR_118 ;
	7'h4c :
		TR_159 = TR_118 ;
	7'h4d :
		TR_159 = TR_118 ;
	7'h4e :
		TR_159 = TR_118 ;
	7'h4f :
		TR_159 = TR_118 ;
	7'h50 :
		TR_159 = TR_118 ;
	7'h51 :
		TR_159 = TR_118 ;
	7'h52 :
		TR_159 = TR_118 ;
	7'h53 :
		TR_159 = TR_118 ;
	7'h54 :
		TR_159 = TR_118 ;
	7'h55 :
		TR_159 = TR_118 ;
	7'h56 :
		TR_159 = TR_118 ;
	7'h57 :
		TR_159 = TR_118 ;
	7'h58 :
		TR_159 = TR_118 ;
	7'h59 :
		TR_159 = TR_118 ;
	7'h5a :
		TR_159 = TR_118 ;
	7'h5b :
		TR_159 = TR_118 ;
	7'h5c :
		TR_159 = TR_118 ;
	7'h5d :
		TR_159 = TR_118 ;
	7'h5e :
		TR_159 = TR_118 ;
	7'h5f :
		TR_159 = TR_118 ;
	7'h60 :
		TR_159 = TR_118 ;
	7'h61 :
		TR_159 = TR_118 ;
	7'h62 :
		TR_159 = TR_118 ;
	7'h63 :
		TR_159 = TR_118 ;
	7'h64 :
		TR_159 = TR_118 ;
	7'h65 :
		TR_159 = TR_118 ;
	7'h66 :
		TR_159 = TR_118 ;
	7'h67 :
		TR_159 = TR_118 ;
	7'h68 :
		TR_159 = TR_118 ;
	7'h69 :
		TR_159 = TR_118 ;
	7'h6a :
		TR_159 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6b :
		TR_159 = TR_118 ;
	7'h6c :
		TR_159 = TR_118 ;
	7'h6d :
		TR_159 = TR_118 ;
	7'h6e :
		TR_159 = TR_118 ;
	7'h6f :
		TR_159 = TR_118 ;
	7'h70 :
		TR_159 = TR_118 ;
	7'h71 :
		TR_159 = TR_118 ;
	7'h72 :
		TR_159 = TR_118 ;
	7'h73 :
		TR_159 = TR_118 ;
	7'h74 :
		TR_159 = TR_118 ;
	7'h75 :
		TR_159 = TR_118 ;
	7'h76 :
		TR_159 = TR_118 ;
	7'h77 :
		TR_159 = TR_118 ;
	7'h78 :
		TR_159 = TR_118 ;
	7'h79 :
		TR_159 = TR_118 ;
	7'h7a :
		TR_159 = TR_118 ;
	7'h7b :
		TR_159 = TR_118 ;
	7'h7c :
		TR_159 = TR_118 ;
	7'h7d :
		TR_159 = TR_118 ;
	7'h7e :
		TR_159 = TR_118 ;
	7'h7f :
		TR_159 = TR_118 ;
	default :
		TR_159 = 9'hx ;
	endcase
always @ ( TR_159 or U_173 or sub8u_71ot or U_183 or RG_rl_182 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_106_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h6a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_106_t = ( ( { 9{ M_180 } } & RG_rl_182 )
		| ( { 9{ U_173 } } & TR_159 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_106_en = ( M_180 | RG_rl_106_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_106_en )
		RG_rl_106 <= RG_rl_106_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_119 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_158 = TR_119 ;
	7'h01 :
		TR_158 = TR_119 ;
	7'h02 :
		TR_158 = TR_119 ;
	7'h03 :
		TR_158 = TR_119 ;
	7'h04 :
		TR_158 = TR_119 ;
	7'h05 :
		TR_158 = TR_119 ;
	7'h06 :
		TR_158 = TR_119 ;
	7'h07 :
		TR_158 = TR_119 ;
	7'h08 :
		TR_158 = TR_119 ;
	7'h09 :
		TR_158 = TR_119 ;
	7'h0a :
		TR_158 = TR_119 ;
	7'h0b :
		TR_158 = TR_119 ;
	7'h0c :
		TR_158 = TR_119 ;
	7'h0d :
		TR_158 = TR_119 ;
	7'h0e :
		TR_158 = TR_119 ;
	7'h0f :
		TR_158 = TR_119 ;
	7'h10 :
		TR_158 = TR_119 ;
	7'h11 :
		TR_158 = TR_119 ;
	7'h12 :
		TR_158 = TR_119 ;
	7'h13 :
		TR_158 = TR_119 ;
	7'h14 :
		TR_158 = TR_119 ;
	7'h15 :
		TR_158 = TR_119 ;
	7'h16 :
		TR_158 = TR_119 ;
	7'h17 :
		TR_158 = TR_119 ;
	7'h18 :
		TR_158 = TR_119 ;
	7'h19 :
		TR_158 = TR_119 ;
	7'h1a :
		TR_158 = TR_119 ;
	7'h1b :
		TR_158 = TR_119 ;
	7'h1c :
		TR_158 = TR_119 ;
	7'h1d :
		TR_158 = TR_119 ;
	7'h1e :
		TR_158 = TR_119 ;
	7'h1f :
		TR_158 = TR_119 ;
	7'h20 :
		TR_158 = TR_119 ;
	7'h21 :
		TR_158 = TR_119 ;
	7'h22 :
		TR_158 = TR_119 ;
	7'h23 :
		TR_158 = TR_119 ;
	7'h24 :
		TR_158 = TR_119 ;
	7'h25 :
		TR_158 = TR_119 ;
	7'h26 :
		TR_158 = TR_119 ;
	7'h27 :
		TR_158 = TR_119 ;
	7'h28 :
		TR_158 = TR_119 ;
	7'h29 :
		TR_158 = TR_119 ;
	7'h2a :
		TR_158 = TR_119 ;
	7'h2b :
		TR_158 = TR_119 ;
	7'h2c :
		TR_158 = TR_119 ;
	7'h2d :
		TR_158 = TR_119 ;
	7'h2e :
		TR_158 = TR_119 ;
	7'h2f :
		TR_158 = TR_119 ;
	7'h30 :
		TR_158 = TR_119 ;
	7'h31 :
		TR_158 = TR_119 ;
	7'h32 :
		TR_158 = TR_119 ;
	7'h33 :
		TR_158 = TR_119 ;
	7'h34 :
		TR_158 = TR_119 ;
	7'h35 :
		TR_158 = TR_119 ;
	7'h36 :
		TR_158 = TR_119 ;
	7'h37 :
		TR_158 = TR_119 ;
	7'h38 :
		TR_158 = TR_119 ;
	7'h39 :
		TR_158 = TR_119 ;
	7'h3a :
		TR_158 = TR_119 ;
	7'h3b :
		TR_158 = TR_119 ;
	7'h3c :
		TR_158 = TR_119 ;
	7'h3d :
		TR_158 = TR_119 ;
	7'h3e :
		TR_158 = TR_119 ;
	7'h3f :
		TR_158 = TR_119 ;
	7'h40 :
		TR_158 = TR_119 ;
	7'h41 :
		TR_158 = TR_119 ;
	7'h42 :
		TR_158 = TR_119 ;
	7'h43 :
		TR_158 = TR_119 ;
	7'h44 :
		TR_158 = TR_119 ;
	7'h45 :
		TR_158 = TR_119 ;
	7'h46 :
		TR_158 = TR_119 ;
	7'h47 :
		TR_158 = TR_119 ;
	7'h48 :
		TR_158 = TR_119 ;
	7'h49 :
		TR_158 = TR_119 ;
	7'h4a :
		TR_158 = TR_119 ;
	7'h4b :
		TR_158 = TR_119 ;
	7'h4c :
		TR_158 = TR_119 ;
	7'h4d :
		TR_158 = TR_119 ;
	7'h4e :
		TR_158 = TR_119 ;
	7'h4f :
		TR_158 = TR_119 ;
	7'h50 :
		TR_158 = TR_119 ;
	7'h51 :
		TR_158 = TR_119 ;
	7'h52 :
		TR_158 = TR_119 ;
	7'h53 :
		TR_158 = TR_119 ;
	7'h54 :
		TR_158 = TR_119 ;
	7'h55 :
		TR_158 = TR_119 ;
	7'h56 :
		TR_158 = TR_119 ;
	7'h57 :
		TR_158 = TR_119 ;
	7'h58 :
		TR_158 = TR_119 ;
	7'h59 :
		TR_158 = TR_119 ;
	7'h5a :
		TR_158 = TR_119 ;
	7'h5b :
		TR_158 = TR_119 ;
	7'h5c :
		TR_158 = TR_119 ;
	7'h5d :
		TR_158 = TR_119 ;
	7'h5e :
		TR_158 = TR_119 ;
	7'h5f :
		TR_158 = TR_119 ;
	7'h60 :
		TR_158 = TR_119 ;
	7'h61 :
		TR_158 = TR_119 ;
	7'h62 :
		TR_158 = TR_119 ;
	7'h63 :
		TR_158 = TR_119 ;
	7'h64 :
		TR_158 = TR_119 ;
	7'h65 :
		TR_158 = TR_119 ;
	7'h66 :
		TR_158 = TR_119 ;
	7'h67 :
		TR_158 = TR_119 ;
	7'h68 :
		TR_158 = TR_119 ;
	7'h69 :
		TR_158 = TR_119 ;
	7'h6a :
		TR_158 = TR_119 ;
	7'h6b :
		TR_158 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6c :
		TR_158 = TR_119 ;
	7'h6d :
		TR_158 = TR_119 ;
	7'h6e :
		TR_158 = TR_119 ;
	7'h6f :
		TR_158 = TR_119 ;
	7'h70 :
		TR_158 = TR_119 ;
	7'h71 :
		TR_158 = TR_119 ;
	7'h72 :
		TR_158 = TR_119 ;
	7'h73 :
		TR_158 = TR_119 ;
	7'h74 :
		TR_158 = TR_119 ;
	7'h75 :
		TR_158 = TR_119 ;
	7'h76 :
		TR_158 = TR_119 ;
	7'h77 :
		TR_158 = TR_119 ;
	7'h78 :
		TR_158 = TR_119 ;
	7'h79 :
		TR_158 = TR_119 ;
	7'h7a :
		TR_158 = TR_119 ;
	7'h7b :
		TR_158 = TR_119 ;
	7'h7c :
		TR_158 = TR_119 ;
	7'h7d :
		TR_158 = TR_119 ;
	7'h7e :
		TR_158 = TR_119 ;
	7'h7f :
		TR_158 = TR_119 ;
	default :
		TR_158 = 9'hx ;
	endcase
always @ ( TR_158 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_51 or 
	U_174 or RG_rl_182 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_107_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h6b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_107_t = ( ( { 9{ ST1_03d } } & RG_rl_182 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_51 )
		| ( { 9{ U_173 } } & TR_158 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_107_en = ( ST1_03d | U_174 | RG_rl_107_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_107_en )
		RG_rl_107 <= RG_rl_107_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_120 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_157 = TR_120 ;
	7'h01 :
		TR_157 = TR_120 ;
	7'h02 :
		TR_157 = TR_120 ;
	7'h03 :
		TR_157 = TR_120 ;
	7'h04 :
		TR_157 = TR_120 ;
	7'h05 :
		TR_157 = TR_120 ;
	7'h06 :
		TR_157 = TR_120 ;
	7'h07 :
		TR_157 = TR_120 ;
	7'h08 :
		TR_157 = TR_120 ;
	7'h09 :
		TR_157 = TR_120 ;
	7'h0a :
		TR_157 = TR_120 ;
	7'h0b :
		TR_157 = TR_120 ;
	7'h0c :
		TR_157 = TR_120 ;
	7'h0d :
		TR_157 = TR_120 ;
	7'h0e :
		TR_157 = TR_120 ;
	7'h0f :
		TR_157 = TR_120 ;
	7'h10 :
		TR_157 = TR_120 ;
	7'h11 :
		TR_157 = TR_120 ;
	7'h12 :
		TR_157 = TR_120 ;
	7'h13 :
		TR_157 = TR_120 ;
	7'h14 :
		TR_157 = TR_120 ;
	7'h15 :
		TR_157 = TR_120 ;
	7'h16 :
		TR_157 = TR_120 ;
	7'h17 :
		TR_157 = TR_120 ;
	7'h18 :
		TR_157 = TR_120 ;
	7'h19 :
		TR_157 = TR_120 ;
	7'h1a :
		TR_157 = TR_120 ;
	7'h1b :
		TR_157 = TR_120 ;
	7'h1c :
		TR_157 = TR_120 ;
	7'h1d :
		TR_157 = TR_120 ;
	7'h1e :
		TR_157 = TR_120 ;
	7'h1f :
		TR_157 = TR_120 ;
	7'h20 :
		TR_157 = TR_120 ;
	7'h21 :
		TR_157 = TR_120 ;
	7'h22 :
		TR_157 = TR_120 ;
	7'h23 :
		TR_157 = TR_120 ;
	7'h24 :
		TR_157 = TR_120 ;
	7'h25 :
		TR_157 = TR_120 ;
	7'h26 :
		TR_157 = TR_120 ;
	7'h27 :
		TR_157 = TR_120 ;
	7'h28 :
		TR_157 = TR_120 ;
	7'h29 :
		TR_157 = TR_120 ;
	7'h2a :
		TR_157 = TR_120 ;
	7'h2b :
		TR_157 = TR_120 ;
	7'h2c :
		TR_157 = TR_120 ;
	7'h2d :
		TR_157 = TR_120 ;
	7'h2e :
		TR_157 = TR_120 ;
	7'h2f :
		TR_157 = TR_120 ;
	7'h30 :
		TR_157 = TR_120 ;
	7'h31 :
		TR_157 = TR_120 ;
	7'h32 :
		TR_157 = TR_120 ;
	7'h33 :
		TR_157 = TR_120 ;
	7'h34 :
		TR_157 = TR_120 ;
	7'h35 :
		TR_157 = TR_120 ;
	7'h36 :
		TR_157 = TR_120 ;
	7'h37 :
		TR_157 = TR_120 ;
	7'h38 :
		TR_157 = TR_120 ;
	7'h39 :
		TR_157 = TR_120 ;
	7'h3a :
		TR_157 = TR_120 ;
	7'h3b :
		TR_157 = TR_120 ;
	7'h3c :
		TR_157 = TR_120 ;
	7'h3d :
		TR_157 = TR_120 ;
	7'h3e :
		TR_157 = TR_120 ;
	7'h3f :
		TR_157 = TR_120 ;
	7'h40 :
		TR_157 = TR_120 ;
	7'h41 :
		TR_157 = TR_120 ;
	7'h42 :
		TR_157 = TR_120 ;
	7'h43 :
		TR_157 = TR_120 ;
	7'h44 :
		TR_157 = TR_120 ;
	7'h45 :
		TR_157 = TR_120 ;
	7'h46 :
		TR_157 = TR_120 ;
	7'h47 :
		TR_157 = TR_120 ;
	7'h48 :
		TR_157 = TR_120 ;
	7'h49 :
		TR_157 = TR_120 ;
	7'h4a :
		TR_157 = TR_120 ;
	7'h4b :
		TR_157 = TR_120 ;
	7'h4c :
		TR_157 = TR_120 ;
	7'h4d :
		TR_157 = TR_120 ;
	7'h4e :
		TR_157 = TR_120 ;
	7'h4f :
		TR_157 = TR_120 ;
	7'h50 :
		TR_157 = TR_120 ;
	7'h51 :
		TR_157 = TR_120 ;
	7'h52 :
		TR_157 = TR_120 ;
	7'h53 :
		TR_157 = TR_120 ;
	7'h54 :
		TR_157 = TR_120 ;
	7'h55 :
		TR_157 = TR_120 ;
	7'h56 :
		TR_157 = TR_120 ;
	7'h57 :
		TR_157 = TR_120 ;
	7'h58 :
		TR_157 = TR_120 ;
	7'h59 :
		TR_157 = TR_120 ;
	7'h5a :
		TR_157 = TR_120 ;
	7'h5b :
		TR_157 = TR_120 ;
	7'h5c :
		TR_157 = TR_120 ;
	7'h5d :
		TR_157 = TR_120 ;
	7'h5e :
		TR_157 = TR_120 ;
	7'h5f :
		TR_157 = TR_120 ;
	7'h60 :
		TR_157 = TR_120 ;
	7'h61 :
		TR_157 = TR_120 ;
	7'h62 :
		TR_157 = TR_120 ;
	7'h63 :
		TR_157 = TR_120 ;
	7'h64 :
		TR_157 = TR_120 ;
	7'h65 :
		TR_157 = TR_120 ;
	7'h66 :
		TR_157 = TR_120 ;
	7'h67 :
		TR_157 = TR_120 ;
	7'h68 :
		TR_157 = TR_120 ;
	7'h69 :
		TR_157 = TR_120 ;
	7'h6a :
		TR_157 = TR_120 ;
	7'h6b :
		TR_157 = TR_120 ;
	7'h6c :
		TR_157 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6d :
		TR_157 = TR_120 ;
	7'h6e :
		TR_157 = TR_120 ;
	7'h6f :
		TR_157 = TR_120 ;
	7'h70 :
		TR_157 = TR_120 ;
	7'h71 :
		TR_157 = TR_120 ;
	7'h72 :
		TR_157 = TR_120 ;
	7'h73 :
		TR_157 = TR_120 ;
	7'h74 :
		TR_157 = TR_120 ;
	7'h75 :
		TR_157 = TR_120 ;
	7'h76 :
		TR_157 = TR_120 ;
	7'h77 :
		TR_157 = TR_120 ;
	7'h78 :
		TR_157 = TR_120 ;
	7'h79 :
		TR_157 = TR_120 ;
	7'h7a :
		TR_157 = TR_120 ;
	7'h7b :
		TR_157 = TR_120 ;
	7'h7c :
		TR_157 = TR_120 ;
	7'h7d :
		TR_157 = TR_120 ;
	7'h7e :
		TR_157 = TR_120 ;
	7'h7f :
		TR_157 = TR_120 ;
	default :
		TR_157 = 9'hx ;
	endcase
always @ ( TR_157 or U_173 or sub8u_71ot or U_183 or RG_rl_183 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_108_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h6c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_108_t = ( ( { 9{ M_180 } } & RG_rl_183 )
		| ( { 9{ U_173 } } & TR_157 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_108_en = ( M_180 | RG_rl_108_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_108_en )
		RG_rl_108 <= RG_rl_108_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_121 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_156 = TR_121 ;
	7'h01 :
		TR_156 = TR_121 ;
	7'h02 :
		TR_156 = TR_121 ;
	7'h03 :
		TR_156 = TR_121 ;
	7'h04 :
		TR_156 = TR_121 ;
	7'h05 :
		TR_156 = TR_121 ;
	7'h06 :
		TR_156 = TR_121 ;
	7'h07 :
		TR_156 = TR_121 ;
	7'h08 :
		TR_156 = TR_121 ;
	7'h09 :
		TR_156 = TR_121 ;
	7'h0a :
		TR_156 = TR_121 ;
	7'h0b :
		TR_156 = TR_121 ;
	7'h0c :
		TR_156 = TR_121 ;
	7'h0d :
		TR_156 = TR_121 ;
	7'h0e :
		TR_156 = TR_121 ;
	7'h0f :
		TR_156 = TR_121 ;
	7'h10 :
		TR_156 = TR_121 ;
	7'h11 :
		TR_156 = TR_121 ;
	7'h12 :
		TR_156 = TR_121 ;
	7'h13 :
		TR_156 = TR_121 ;
	7'h14 :
		TR_156 = TR_121 ;
	7'h15 :
		TR_156 = TR_121 ;
	7'h16 :
		TR_156 = TR_121 ;
	7'h17 :
		TR_156 = TR_121 ;
	7'h18 :
		TR_156 = TR_121 ;
	7'h19 :
		TR_156 = TR_121 ;
	7'h1a :
		TR_156 = TR_121 ;
	7'h1b :
		TR_156 = TR_121 ;
	7'h1c :
		TR_156 = TR_121 ;
	7'h1d :
		TR_156 = TR_121 ;
	7'h1e :
		TR_156 = TR_121 ;
	7'h1f :
		TR_156 = TR_121 ;
	7'h20 :
		TR_156 = TR_121 ;
	7'h21 :
		TR_156 = TR_121 ;
	7'h22 :
		TR_156 = TR_121 ;
	7'h23 :
		TR_156 = TR_121 ;
	7'h24 :
		TR_156 = TR_121 ;
	7'h25 :
		TR_156 = TR_121 ;
	7'h26 :
		TR_156 = TR_121 ;
	7'h27 :
		TR_156 = TR_121 ;
	7'h28 :
		TR_156 = TR_121 ;
	7'h29 :
		TR_156 = TR_121 ;
	7'h2a :
		TR_156 = TR_121 ;
	7'h2b :
		TR_156 = TR_121 ;
	7'h2c :
		TR_156 = TR_121 ;
	7'h2d :
		TR_156 = TR_121 ;
	7'h2e :
		TR_156 = TR_121 ;
	7'h2f :
		TR_156 = TR_121 ;
	7'h30 :
		TR_156 = TR_121 ;
	7'h31 :
		TR_156 = TR_121 ;
	7'h32 :
		TR_156 = TR_121 ;
	7'h33 :
		TR_156 = TR_121 ;
	7'h34 :
		TR_156 = TR_121 ;
	7'h35 :
		TR_156 = TR_121 ;
	7'h36 :
		TR_156 = TR_121 ;
	7'h37 :
		TR_156 = TR_121 ;
	7'h38 :
		TR_156 = TR_121 ;
	7'h39 :
		TR_156 = TR_121 ;
	7'h3a :
		TR_156 = TR_121 ;
	7'h3b :
		TR_156 = TR_121 ;
	7'h3c :
		TR_156 = TR_121 ;
	7'h3d :
		TR_156 = TR_121 ;
	7'h3e :
		TR_156 = TR_121 ;
	7'h3f :
		TR_156 = TR_121 ;
	7'h40 :
		TR_156 = TR_121 ;
	7'h41 :
		TR_156 = TR_121 ;
	7'h42 :
		TR_156 = TR_121 ;
	7'h43 :
		TR_156 = TR_121 ;
	7'h44 :
		TR_156 = TR_121 ;
	7'h45 :
		TR_156 = TR_121 ;
	7'h46 :
		TR_156 = TR_121 ;
	7'h47 :
		TR_156 = TR_121 ;
	7'h48 :
		TR_156 = TR_121 ;
	7'h49 :
		TR_156 = TR_121 ;
	7'h4a :
		TR_156 = TR_121 ;
	7'h4b :
		TR_156 = TR_121 ;
	7'h4c :
		TR_156 = TR_121 ;
	7'h4d :
		TR_156 = TR_121 ;
	7'h4e :
		TR_156 = TR_121 ;
	7'h4f :
		TR_156 = TR_121 ;
	7'h50 :
		TR_156 = TR_121 ;
	7'h51 :
		TR_156 = TR_121 ;
	7'h52 :
		TR_156 = TR_121 ;
	7'h53 :
		TR_156 = TR_121 ;
	7'h54 :
		TR_156 = TR_121 ;
	7'h55 :
		TR_156 = TR_121 ;
	7'h56 :
		TR_156 = TR_121 ;
	7'h57 :
		TR_156 = TR_121 ;
	7'h58 :
		TR_156 = TR_121 ;
	7'h59 :
		TR_156 = TR_121 ;
	7'h5a :
		TR_156 = TR_121 ;
	7'h5b :
		TR_156 = TR_121 ;
	7'h5c :
		TR_156 = TR_121 ;
	7'h5d :
		TR_156 = TR_121 ;
	7'h5e :
		TR_156 = TR_121 ;
	7'h5f :
		TR_156 = TR_121 ;
	7'h60 :
		TR_156 = TR_121 ;
	7'h61 :
		TR_156 = TR_121 ;
	7'h62 :
		TR_156 = TR_121 ;
	7'h63 :
		TR_156 = TR_121 ;
	7'h64 :
		TR_156 = TR_121 ;
	7'h65 :
		TR_156 = TR_121 ;
	7'h66 :
		TR_156 = TR_121 ;
	7'h67 :
		TR_156 = TR_121 ;
	7'h68 :
		TR_156 = TR_121 ;
	7'h69 :
		TR_156 = TR_121 ;
	7'h6a :
		TR_156 = TR_121 ;
	7'h6b :
		TR_156 = TR_121 ;
	7'h6c :
		TR_156 = TR_121 ;
	7'h6d :
		TR_156 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6e :
		TR_156 = TR_121 ;
	7'h6f :
		TR_156 = TR_121 ;
	7'h70 :
		TR_156 = TR_121 ;
	7'h71 :
		TR_156 = TR_121 ;
	7'h72 :
		TR_156 = TR_121 ;
	7'h73 :
		TR_156 = TR_121 ;
	7'h74 :
		TR_156 = TR_121 ;
	7'h75 :
		TR_156 = TR_121 ;
	7'h76 :
		TR_156 = TR_121 ;
	7'h77 :
		TR_156 = TR_121 ;
	7'h78 :
		TR_156 = TR_121 ;
	7'h79 :
		TR_156 = TR_121 ;
	7'h7a :
		TR_156 = TR_121 ;
	7'h7b :
		TR_156 = TR_121 ;
	7'h7c :
		TR_156 = TR_121 ;
	7'h7d :
		TR_156 = TR_121 ;
	7'h7e :
		TR_156 = TR_121 ;
	7'h7f :
		TR_156 = TR_121 ;
	default :
		TR_156 = 9'hx ;
	endcase
always @ ( TR_156 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_52 or 
	U_174 or RG_rl_183 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_109_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h6d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_109_t = ( ( { 9{ ST1_03d } } & RG_rl_183 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_52 )
		| ( { 9{ U_173 } } & TR_156 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_109_en = ( ST1_03d | U_174 | RG_rl_109_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_109_en )
		RG_rl_109 <= RG_rl_109_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_122 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_155 = TR_122 ;
	7'h01 :
		TR_155 = TR_122 ;
	7'h02 :
		TR_155 = TR_122 ;
	7'h03 :
		TR_155 = TR_122 ;
	7'h04 :
		TR_155 = TR_122 ;
	7'h05 :
		TR_155 = TR_122 ;
	7'h06 :
		TR_155 = TR_122 ;
	7'h07 :
		TR_155 = TR_122 ;
	7'h08 :
		TR_155 = TR_122 ;
	7'h09 :
		TR_155 = TR_122 ;
	7'h0a :
		TR_155 = TR_122 ;
	7'h0b :
		TR_155 = TR_122 ;
	7'h0c :
		TR_155 = TR_122 ;
	7'h0d :
		TR_155 = TR_122 ;
	7'h0e :
		TR_155 = TR_122 ;
	7'h0f :
		TR_155 = TR_122 ;
	7'h10 :
		TR_155 = TR_122 ;
	7'h11 :
		TR_155 = TR_122 ;
	7'h12 :
		TR_155 = TR_122 ;
	7'h13 :
		TR_155 = TR_122 ;
	7'h14 :
		TR_155 = TR_122 ;
	7'h15 :
		TR_155 = TR_122 ;
	7'h16 :
		TR_155 = TR_122 ;
	7'h17 :
		TR_155 = TR_122 ;
	7'h18 :
		TR_155 = TR_122 ;
	7'h19 :
		TR_155 = TR_122 ;
	7'h1a :
		TR_155 = TR_122 ;
	7'h1b :
		TR_155 = TR_122 ;
	7'h1c :
		TR_155 = TR_122 ;
	7'h1d :
		TR_155 = TR_122 ;
	7'h1e :
		TR_155 = TR_122 ;
	7'h1f :
		TR_155 = TR_122 ;
	7'h20 :
		TR_155 = TR_122 ;
	7'h21 :
		TR_155 = TR_122 ;
	7'h22 :
		TR_155 = TR_122 ;
	7'h23 :
		TR_155 = TR_122 ;
	7'h24 :
		TR_155 = TR_122 ;
	7'h25 :
		TR_155 = TR_122 ;
	7'h26 :
		TR_155 = TR_122 ;
	7'h27 :
		TR_155 = TR_122 ;
	7'h28 :
		TR_155 = TR_122 ;
	7'h29 :
		TR_155 = TR_122 ;
	7'h2a :
		TR_155 = TR_122 ;
	7'h2b :
		TR_155 = TR_122 ;
	7'h2c :
		TR_155 = TR_122 ;
	7'h2d :
		TR_155 = TR_122 ;
	7'h2e :
		TR_155 = TR_122 ;
	7'h2f :
		TR_155 = TR_122 ;
	7'h30 :
		TR_155 = TR_122 ;
	7'h31 :
		TR_155 = TR_122 ;
	7'h32 :
		TR_155 = TR_122 ;
	7'h33 :
		TR_155 = TR_122 ;
	7'h34 :
		TR_155 = TR_122 ;
	7'h35 :
		TR_155 = TR_122 ;
	7'h36 :
		TR_155 = TR_122 ;
	7'h37 :
		TR_155 = TR_122 ;
	7'h38 :
		TR_155 = TR_122 ;
	7'h39 :
		TR_155 = TR_122 ;
	7'h3a :
		TR_155 = TR_122 ;
	7'h3b :
		TR_155 = TR_122 ;
	7'h3c :
		TR_155 = TR_122 ;
	7'h3d :
		TR_155 = TR_122 ;
	7'h3e :
		TR_155 = TR_122 ;
	7'h3f :
		TR_155 = TR_122 ;
	7'h40 :
		TR_155 = TR_122 ;
	7'h41 :
		TR_155 = TR_122 ;
	7'h42 :
		TR_155 = TR_122 ;
	7'h43 :
		TR_155 = TR_122 ;
	7'h44 :
		TR_155 = TR_122 ;
	7'h45 :
		TR_155 = TR_122 ;
	7'h46 :
		TR_155 = TR_122 ;
	7'h47 :
		TR_155 = TR_122 ;
	7'h48 :
		TR_155 = TR_122 ;
	7'h49 :
		TR_155 = TR_122 ;
	7'h4a :
		TR_155 = TR_122 ;
	7'h4b :
		TR_155 = TR_122 ;
	7'h4c :
		TR_155 = TR_122 ;
	7'h4d :
		TR_155 = TR_122 ;
	7'h4e :
		TR_155 = TR_122 ;
	7'h4f :
		TR_155 = TR_122 ;
	7'h50 :
		TR_155 = TR_122 ;
	7'h51 :
		TR_155 = TR_122 ;
	7'h52 :
		TR_155 = TR_122 ;
	7'h53 :
		TR_155 = TR_122 ;
	7'h54 :
		TR_155 = TR_122 ;
	7'h55 :
		TR_155 = TR_122 ;
	7'h56 :
		TR_155 = TR_122 ;
	7'h57 :
		TR_155 = TR_122 ;
	7'h58 :
		TR_155 = TR_122 ;
	7'h59 :
		TR_155 = TR_122 ;
	7'h5a :
		TR_155 = TR_122 ;
	7'h5b :
		TR_155 = TR_122 ;
	7'h5c :
		TR_155 = TR_122 ;
	7'h5d :
		TR_155 = TR_122 ;
	7'h5e :
		TR_155 = TR_122 ;
	7'h5f :
		TR_155 = TR_122 ;
	7'h60 :
		TR_155 = TR_122 ;
	7'h61 :
		TR_155 = TR_122 ;
	7'h62 :
		TR_155 = TR_122 ;
	7'h63 :
		TR_155 = TR_122 ;
	7'h64 :
		TR_155 = TR_122 ;
	7'h65 :
		TR_155 = TR_122 ;
	7'h66 :
		TR_155 = TR_122 ;
	7'h67 :
		TR_155 = TR_122 ;
	7'h68 :
		TR_155 = TR_122 ;
	7'h69 :
		TR_155 = TR_122 ;
	7'h6a :
		TR_155 = TR_122 ;
	7'h6b :
		TR_155 = TR_122 ;
	7'h6c :
		TR_155 = TR_122 ;
	7'h6d :
		TR_155 = TR_122 ;
	7'h6e :
		TR_155 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6f :
		TR_155 = TR_122 ;
	7'h70 :
		TR_155 = TR_122 ;
	7'h71 :
		TR_155 = TR_122 ;
	7'h72 :
		TR_155 = TR_122 ;
	7'h73 :
		TR_155 = TR_122 ;
	7'h74 :
		TR_155 = TR_122 ;
	7'h75 :
		TR_155 = TR_122 ;
	7'h76 :
		TR_155 = TR_122 ;
	7'h77 :
		TR_155 = TR_122 ;
	7'h78 :
		TR_155 = TR_122 ;
	7'h79 :
		TR_155 = TR_122 ;
	7'h7a :
		TR_155 = TR_122 ;
	7'h7b :
		TR_155 = TR_122 ;
	7'h7c :
		TR_155 = TR_122 ;
	7'h7d :
		TR_155 = TR_122 ;
	7'h7e :
		TR_155 = TR_122 ;
	7'h7f :
		TR_155 = TR_122 ;
	default :
		TR_155 = 9'hx ;
	endcase
always @ ( TR_155 or U_173 or sub8u_71ot or U_183 or RG_rl_184 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_110_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h6e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_110_t = ( ( { 9{ M_180 } } & RG_rl_184 )
		| ( { 9{ U_173 } } & TR_155 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_110_en = ( M_180 | RG_rl_110_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_110_en )
		RG_rl_110 <= RG_rl_110_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_123 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_154 = TR_123 ;
	7'h01 :
		TR_154 = TR_123 ;
	7'h02 :
		TR_154 = TR_123 ;
	7'h03 :
		TR_154 = TR_123 ;
	7'h04 :
		TR_154 = TR_123 ;
	7'h05 :
		TR_154 = TR_123 ;
	7'h06 :
		TR_154 = TR_123 ;
	7'h07 :
		TR_154 = TR_123 ;
	7'h08 :
		TR_154 = TR_123 ;
	7'h09 :
		TR_154 = TR_123 ;
	7'h0a :
		TR_154 = TR_123 ;
	7'h0b :
		TR_154 = TR_123 ;
	7'h0c :
		TR_154 = TR_123 ;
	7'h0d :
		TR_154 = TR_123 ;
	7'h0e :
		TR_154 = TR_123 ;
	7'h0f :
		TR_154 = TR_123 ;
	7'h10 :
		TR_154 = TR_123 ;
	7'h11 :
		TR_154 = TR_123 ;
	7'h12 :
		TR_154 = TR_123 ;
	7'h13 :
		TR_154 = TR_123 ;
	7'h14 :
		TR_154 = TR_123 ;
	7'h15 :
		TR_154 = TR_123 ;
	7'h16 :
		TR_154 = TR_123 ;
	7'h17 :
		TR_154 = TR_123 ;
	7'h18 :
		TR_154 = TR_123 ;
	7'h19 :
		TR_154 = TR_123 ;
	7'h1a :
		TR_154 = TR_123 ;
	7'h1b :
		TR_154 = TR_123 ;
	7'h1c :
		TR_154 = TR_123 ;
	7'h1d :
		TR_154 = TR_123 ;
	7'h1e :
		TR_154 = TR_123 ;
	7'h1f :
		TR_154 = TR_123 ;
	7'h20 :
		TR_154 = TR_123 ;
	7'h21 :
		TR_154 = TR_123 ;
	7'h22 :
		TR_154 = TR_123 ;
	7'h23 :
		TR_154 = TR_123 ;
	7'h24 :
		TR_154 = TR_123 ;
	7'h25 :
		TR_154 = TR_123 ;
	7'h26 :
		TR_154 = TR_123 ;
	7'h27 :
		TR_154 = TR_123 ;
	7'h28 :
		TR_154 = TR_123 ;
	7'h29 :
		TR_154 = TR_123 ;
	7'h2a :
		TR_154 = TR_123 ;
	7'h2b :
		TR_154 = TR_123 ;
	7'h2c :
		TR_154 = TR_123 ;
	7'h2d :
		TR_154 = TR_123 ;
	7'h2e :
		TR_154 = TR_123 ;
	7'h2f :
		TR_154 = TR_123 ;
	7'h30 :
		TR_154 = TR_123 ;
	7'h31 :
		TR_154 = TR_123 ;
	7'h32 :
		TR_154 = TR_123 ;
	7'h33 :
		TR_154 = TR_123 ;
	7'h34 :
		TR_154 = TR_123 ;
	7'h35 :
		TR_154 = TR_123 ;
	7'h36 :
		TR_154 = TR_123 ;
	7'h37 :
		TR_154 = TR_123 ;
	7'h38 :
		TR_154 = TR_123 ;
	7'h39 :
		TR_154 = TR_123 ;
	7'h3a :
		TR_154 = TR_123 ;
	7'h3b :
		TR_154 = TR_123 ;
	7'h3c :
		TR_154 = TR_123 ;
	7'h3d :
		TR_154 = TR_123 ;
	7'h3e :
		TR_154 = TR_123 ;
	7'h3f :
		TR_154 = TR_123 ;
	7'h40 :
		TR_154 = TR_123 ;
	7'h41 :
		TR_154 = TR_123 ;
	7'h42 :
		TR_154 = TR_123 ;
	7'h43 :
		TR_154 = TR_123 ;
	7'h44 :
		TR_154 = TR_123 ;
	7'h45 :
		TR_154 = TR_123 ;
	7'h46 :
		TR_154 = TR_123 ;
	7'h47 :
		TR_154 = TR_123 ;
	7'h48 :
		TR_154 = TR_123 ;
	7'h49 :
		TR_154 = TR_123 ;
	7'h4a :
		TR_154 = TR_123 ;
	7'h4b :
		TR_154 = TR_123 ;
	7'h4c :
		TR_154 = TR_123 ;
	7'h4d :
		TR_154 = TR_123 ;
	7'h4e :
		TR_154 = TR_123 ;
	7'h4f :
		TR_154 = TR_123 ;
	7'h50 :
		TR_154 = TR_123 ;
	7'h51 :
		TR_154 = TR_123 ;
	7'h52 :
		TR_154 = TR_123 ;
	7'h53 :
		TR_154 = TR_123 ;
	7'h54 :
		TR_154 = TR_123 ;
	7'h55 :
		TR_154 = TR_123 ;
	7'h56 :
		TR_154 = TR_123 ;
	7'h57 :
		TR_154 = TR_123 ;
	7'h58 :
		TR_154 = TR_123 ;
	7'h59 :
		TR_154 = TR_123 ;
	7'h5a :
		TR_154 = TR_123 ;
	7'h5b :
		TR_154 = TR_123 ;
	7'h5c :
		TR_154 = TR_123 ;
	7'h5d :
		TR_154 = TR_123 ;
	7'h5e :
		TR_154 = TR_123 ;
	7'h5f :
		TR_154 = TR_123 ;
	7'h60 :
		TR_154 = TR_123 ;
	7'h61 :
		TR_154 = TR_123 ;
	7'h62 :
		TR_154 = TR_123 ;
	7'h63 :
		TR_154 = TR_123 ;
	7'h64 :
		TR_154 = TR_123 ;
	7'h65 :
		TR_154 = TR_123 ;
	7'h66 :
		TR_154 = TR_123 ;
	7'h67 :
		TR_154 = TR_123 ;
	7'h68 :
		TR_154 = TR_123 ;
	7'h69 :
		TR_154 = TR_123 ;
	7'h6a :
		TR_154 = TR_123 ;
	7'h6b :
		TR_154 = TR_123 ;
	7'h6c :
		TR_154 = TR_123 ;
	7'h6d :
		TR_154 = TR_123 ;
	7'h6e :
		TR_154 = TR_123 ;
	7'h6f :
		TR_154 = 9'h000 ;	// line#=../rle.cpp:80
	7'h70 :
		TR_154 = TR_123 ;
	7'h71 :
		TR_154 = TR_123 ;
	7'h72 :
		TR_154 = TR_123 ;
	7'h73 :
		TR_154 = TR_123 ;
	7'h74 :
		TR_154 = TR_123 ;
	7'h75 :
		TR_154 = TR_123 ;
	7'h76 :
		TR_154 = TR_123 ;
	7'h77 :
		TR_154 = TR_123 ;
	7'h78 :
		TR_154 = TR_123 ;
	7'h79 :
		TR_154 = TR_123 ;
	7'h7a :
		TR_154 = TR_123 ;
	7'h7b :
		TR_154 = TR_123 ;
	7'h7c :
		TR_154 = TR_123 ;
	7'h7d :
		TR_154 = TR_123 ;
	7'h7e :
		TR_154 = TR_123 ;
	7'h7f :
		TR_154 = TR_123 ;
	default :
		TR_154 = 9'hx ;
	endcase
always @ ( TR_154 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_53 or 
	U_174 or RG_rl_184 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_111_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h6f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_111_t = ( ( { 9{ ST1_03d } } & RG_rl_184 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_53 )
		| ( { 9{ U_173 } } & TR_154 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_111_en = ( ST1_03d | U_174 | RG_rl_111_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_111_en )
		RG_rl_111 <= RG_rl_111_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_124 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_153 = TR_124 ;
	7'h01 :
		TR_153 = TR_124 ;
	7'h02 :
		TR_153 = TR_124 ;
	7'h03 :
		TR_153 = TR_124 ;
	7'h04 :
		TR_153 = TR_124 ;
	7'h05 :
		TR_153 = TR_124 ;
	7'h06 :
		TR_153 = TR_124 ;
	7'h07 :
		TR_153 = TR_124 ;
	7'h08 :
		TR_153 = TR_124 ;
	7'h09 :
		TR_153 = TR_124 ;
	7'h0a :
		TR_153 = TR_124 ;
	7'h0b :
		TR_153 = TR_124 ;
	7'h0c :
		TR_153 = TR_124 ;
	7'h0d :
		TR_153 = TR_124 ;
	7'h0e :
		TR_153 = TR_124 ;
	7'h0f :
		TR_153 = TR_124 ;
	7'h10 :
		TR_153 = TR_124 ;
	7'h11 :
		TR_153 = TR_124 ;
	7'h12 :
		TR_153 = TR_124 ;
	7'h13 :
		TR_153 = TR_124 ;
	7'h14 :
		TR_153 = TR_124 ;
	7'h15 :
		TR_153 = TR_124 ;
	7'h16 :
		TR_153 = TR_124 ;
	7'h17 :
		TR_153 = TR_124 ;
	7'h18 :
		TR_153 = TR_124 ;
	7'h19 :
		TR_153 = TR_124 ;
	7'h1a :
		TR_153 = TR_124 ;
	7'h1b :
		TR_153 = TR_124 ;
	7'h1c :
		TR_153 = TR_124 ;
	7'h1d :
		TR_153 = TR_124 ;
	7'h1e :
		TR_153 = TR_124 ;
	7'h1f :
		TR_153 = TR_124 ;
	7'h20 :
		TR_153 = TR_124 ;
	7'h21 :
		TR_153 = TR_124 ;
	7'h22 :
		TR_153 = TR_124 ;
	7'h23 :
		TR_153 = TR_124 ;
	7'h24 :
		TR_153 = TR_124 ;
	7'h25 :
		TR_153 = TR_124 ;
	7'h26 :
		TR_153 = TR_124 ;
	7'h27 :
		TR_153 = TR_124 ;
	7'h28 :
		TR_153 = TR_124 ;
	7'h29 :
		TR_153 = TR_124 ;
	7'h2a :
		TR_153 = TR_124 ;
	7'h2b :
		TR_153 = TR_124 ;
	7'h2c :
		TR_153 = TR_124 ;
	7'h2d :
		TR_153 = TR_124 ;
	7'h2e :
		TR_153 = TR_124 ;
	7'h2f :
		TR_153 = TR_124 ;
	7'h30 :
		TR_153 = TR_124 ;
	7'h31 :
		TR_153 = TR_124 ;
	7'h32 :
		TR_153 = TR_124 ;
	7'h33 :
		TR_153 = TR_124 ;
	7'h34 :
		TR_153 = TR_124 ;
	7'h35 :
		TR_153 = TR_124 ;
	7'h36 :
		TR_153 = TR_124 ;
	7'h37 :
		TR_153 = TR_124 ;
	7'h38 :
		TR_153 = TR_124 ;
	7'h39 :
		TR_153 = TR_124 ;
	7'h3a :
		TR_153 = TR_124 ;
	7'h3b :
		TR_153 = TR_124 ;
	7'h3c :
		TR_153 = TR_124 ;
	7'h3d :
		TR_153 = TR_124 ;
	7'h3e :
		TR_153 = TR_124 ;
	7'h3f :
		TR_153 = TR_124 ;
	7'h40 :
		TR_153 = TR_124 ;
	7'h41 :
		TR_153 = TR_124 ;
	7'h42 :
		TR_153 = TR_124 ;
	7'h43 :
		TR_153 = TR_124 ;
	7'h44 :
		TR_153 = TR_124 ;
	7'h45 :
		TR_153 = TR_124 ;
	7'h46 :
		TR_153 = TR_124 ;
	7'h47 :
		TR_153 = TR_124 ;
	7'h48 :
		TR_153 = TR_124 ;
	7'h49 :
		TR_153 = TR_124 ;
	7'h4a :
		TR_153 = TR_124 ;
	7'h4b :
		TR_153 = TR_124 ;
	7'h4c :
		TR_153 = TR_124 ;
	7'h4d :
		TR_153 = TR_124 ;
	7'h4e :
		TR_153 = TR_124 ;
	7'h4f :
		TR_153 = TR_124 ;
	7'h50 :
		TR_153 = TR_124 ;
	7'h51 :
		TR_153 = TR_124 ;
	7'h52 :
		TR_153 = TR_124 ;
	7'h53 :
		TR_153 = TR_124 ;
	7'h54 :
		TR_153 = TR_124 ;
	7'h55 :
		TR_153 = TR_124 ;
	7'h56 :
		TR_153 = TR_124 ;
	7'h57 :
		TR_153 = TR_124 ;
	7'h58 :
		TR_153 = TR_124 ;
	7'h59 :
		TR_153 = TR_124 ;
	7'h5a :
		TR_153 = TR_124 ;
	7'h5b :
		TR_153 = TR_124 ;
	7'h5c :
		TR_153 = TR_124 ;
	7'h5d :
		TR_153 = TR_124 ;
	7'h5e :
		TR_153 = TR_124 ;
	7'h5f :
		TR_153 = TR_124 ;
	7'h60 :
		TR_153 = TR_124 ;
	7'h61 :
		TR_153 = TR_124 ;
	7'h62 :
		TR_153 = TR_124 ;
	7'h63 :
		TR_153 = TR_124 ;
	7'h64 :
		TR_153 = TR_124 ;
	7'h65 :
		TR_153 = TR_124 ;
	7'h66 :
		TR_153 = TR_124 ;
	7'h67 :
		TR_153 = TR_124 ;
	7'h68 :
		TR_153 = TR_124 ;
	7'h69 :
		TR_153 = TR_124 ;
	7'h6a :
		TR_153 = TR_124 ;
	7'h6b :
		TR_153 = TR_124 ;
	7'h6c :
		TR_153 = TR_124 ;
	7'h6d :
		TR_153 = TR_124 ;
	7'h6e :
		TR_153 = TR_124 ;
	7'h6f :
		TR_153 = TR_124 ;
	7'h70 :
		TR_153 = 9'h000 ;	// line#=../rle.cpp:80
	7'h71 :
		TR_153 = TR_124 ;
	7'h72 :
		TR_153 = TR_124 ;
	7'h73 :
		TR_153 = TR_124 ;
	7'h74 :
		TR_153 = TR_124 ;
	7'h75 :
		TR_153 = TR_124 ;
	7'h76 :
		TR_153 = TR_124 ;
	7'h77 :
		TR_153 = TR_124 ;
	7'h78 :
		TR_153 = TR_124 ;
	7'h79 :
		TR_153 = TR_124 ;
	7'h7a :
		TR_153 = TR_124 ;
	7'h7b :
		TR_153 = TR_124 ;
	7'h7c :
		TR_153 = TR_124 ;
	7'h7d :
		TR_153 = TR_124 ;
	7'h7e :
		TR_153 = TR_124 ;
	7'h7f :
		TR_153 = TR_124 ;
	default :
		TR_153 = 9'hx ;
	endcase
always @ ( TR_153 or U_173 or sub8u_71ot or U_183 or RG_rl_185 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_112_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h70 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_112_t = ( ( { 9{ M_180 } } & RG_rl_185 )
		| ( { 9{ U_173 } } & TR_153 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_112_en = ( M_180 | RG_rl_112_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_112_en )
		RG_rl_112 <= RG_rl_112_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_125 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_152 = TR_125 ;
	7'h01 :
		TR_152 = TR_125 ;
	7'h02 :
		TR_152 = TR_125 ;
	7'h03 :
		TR_152 = TR_125 ;
	7'h04 :
		TR_152 = TR_125 ;
	7'h05 :
		TR_152 = TR_125 ;
	7'h06 :
		TR_152 = TR_125 ;
	7'h07 :
		TR_152 = TR_125 ;
	7'h08 :
		TR_152 = TR_125 ;
	7'h09 :
		TR_152 = TR_125 ;
	7'h0a :
		TR_152 = TR_125 ;
	7'h0b :
		TR_152 = TR_125 ;
	7'h0c :
		TR_152 = TR_125 ;
	7'h0d :
		TR_152 = TR_125 ;
	7'h0e :
		TR_152 = TR_125 ;
	7'h0f :
		TR_152 = TR_125 ;
	7'h10 :
		TR_152 = TR_125 ;
	7'h11 :
		TR_152 = TR_125 ;
	7'h12 :
		TR_152 = TR_125 ;
	7'h13 :
		TR_152 = TR_125 ;
	7'h14 :
		TR_152 = TR_125 ;
	7'h15 :
		TR_152 = TR_125 ;
	7'h16 :
		TR_152 = TR_125 ;
	7'h17 :
		TR_152 = TR_125 ;
	7'h18 :
		TR_152 = TR_125 ;
	7'h19 :
		TR_152 = TR_125 ;
	7'h1a :
		TR_152 = TR_125 ;
	7'h1b :
		TR_152 = TR_125 ;
	7'h1c :
		TR_152 = TR_125 ;
	7'h1d :
		TR_152 = TR_125 ;
	7'h1e :
		TR_152 = TR_125 ;
	7'h1f :
		TR_152 = TR_125 ;
	7'h20 :
		TR_152 = TR_125 ;
	7'h21 :
		TR_152 = TR_125 ;
	7'h22 :
		TR_152 = TR_125 ;
	7'h23 :
		TR_152 = TR_125 ;
	7'h24 :
		TR_152 = TR_125 ;
	7'h25 :
		TR_152 = TR_125 ;
	7'h26 :
		TR_152 = TR_125 ;
	7'h27 :
		TR_152 = TR_125 ;
	7'h28 :
		TR_152 = TR_125 ;
	7'h29 :
		TR_152 = TR_125 ;
	7'h2a :
		TR_152 = TR_125 ;
	7'h2b :
		TR_152 = TR_125 ;
	7'h2c :
		TR_152 = TR_125 ;
	7'h2d :
		TR_152 = TR_125 ;
	7'h2e :
		TR_152 = TR_125 ;
	7'h2f :
		TR_152 = TR_125 ;
	7'h30 :
		TR_152 = TR_125 ;
	7'h31 :
		TR_152 = TR_125 ;
	7'h32 :
		TR_152 = TR_125 ;
	7'h33 :
		TR_152 = TR_125 ;
	7'h34 :
		TR_152 = TR_125 ;
	7'h35 :
		TR_152 = TR_125 ;
	7'h36 :
		TR_152 = TR_125 ;
	7'h37 :
		TR_152 = TR_125 ;
	7'h38 :
		TR_152 = TR_125 ;
	7'h39 :
		TR_152 = TR_125 ;
	7'h3a :
		TR_152 = TR_125 ;
	7'h3b :
		TR_152 = TR_125 ;
	7'h3c :
		TR_152 = TR_125 ;
	7'h3d :
		TR_152 = TR_125 ;
	7'h3e :
		TR_152 = TR_125 ;
	7'h3f :
		TR_152 = TR_125 ;
	7'h40 :
		TR_152 = TR_125 ;
	7'h41 :
		TR_152 = TR_125 ;
	7'h42 :
		TR_152 = TR_125 ;
	7'h43 :
		TR_152 = TR_125 ;
	7'h44 :
		TR_152 = TR_125 ;
	7'h45 :
		TR_152 = TR_125 ;
	7'h46 :
		TR_152 = TR_125 ;
	7'h47 :
		TR_152 = TR_125 ;
	7'h48 :
		TR_152 = TR_125 ;
	7'h49 :
		TR_152 = TR_125 ;
	7'h4a :
		TR_152 = TR_125 ;
	7'h4b :
		TR_152 = TR_125 ;
	7'h4c :
		TR_152 = TR_125 ;
	7'h4d :
		TR_152 = TR_125 ;
	7'h4e :
		TR_152 = TR_125 ;
	7'h4f :
		TR_152 = TR_125 ;
	7'h50 :
		TR_152 = TR_125 ;
	7'h51 :
		TR_152 = TR_125 ;
	7'h52 :
		TR_152 = TR_125 ;
	7'h53 :
		TR_152 = TR_125 ;
	7'h54 :
		TR_152 = TR_125 ;
	7'h55 :
		TR_152 = TR_125 ;
	7'h56 :
		TR_152 = TR_125 ;
	7'h57 :
		TR_152 = TR_125 ;
	7'h58 :
		TR_152 = TR_125 ;
	7'h59 :
		TR_152 = TR_125 ;
	7'h5a :
		TR_152 = TR_125 ;
	7'h5b :
		TR_152 = TR_125 ;
	7'h5c :
		TR_152 = TR_125 ;
	7'h5d :
		TR_152 = TR_125 ;
	7'h5e :
		TR_152 = TR_125 ;
	7'h5f :
		TR_152 = TR_125 ;
	7'h60 :
		TR_152 = TR_125 ;
	7'h61 :
		TR_152 = TR_125 ;
	7'h62 :
		TR_152 = TR_125 ;
	7'h63 :
		TR_152 = TR_125 ;
	7'h64 :
		TR_152 = TR_125 ;
	7'h65 :
		TR_152 = TR_125 ;
	7'h66 :
		TR_152 = TR_125 ;
	7'h67 :
		TR_152 = TR_125 ;
	7'h68 :
		TR_152 = TR_125 ;
	7'h69 :
		TR_152 = TR_125 ;
	7'h6a :
		TR_152 = TR_125 ;
	7'h6b :
		TR_152 = TR_125 ;
	7'h6c :
		TR_152 = TR_125 ;
	7'h6d :
		TR_152 = TR_125 ;
	7'h6e :
		TR_152 = TR_125 ;
	7'h6f :
		TR_152 = TR_125 ;
	7'h70 :
		TR_152 = TR_125 ;
	7'h71 :
		TR_152 = 9'h000 ;	// line#=../rle.cpp:80
	7'h72 :
		TR_152 = TR_125 ;
	7'h73 :
		TR_152 = TR_125 ;
	7'h74 :
		TR_152 = TR_125 ;
	7'h75 :
		TR_152 = TR_125 ;
	7'h76 :
		TR_152 = TR_125 ;
	7'h77 :
		TR_152 = TR_125 ;
	7'h78 :
		TR_152 = TR_125 ;
	7'h79 :
		TR_152 = TR_125 ;
	7'h7a :
		TR_152 = TR_125 ;
	7'h7b :
		TR_152 = TR_125 ;
	7'h7c :
		TR_152 = TR_125 ;
	7'h7d :
		TR_152 = TR_125 ;
	7'h7e :
		TR_152 = TR_125 ;
	7'h7f :
		TR_152 = TR_125 ;
	default :
		TR_152 = 9'hx ;
	endcase
always @ ( TR_152 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_54 or 
	U_174 or RG_rl_185 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_113_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h71 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_113_t = ( ( { 9{ ST1_03d } } & RG_rl_185 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_54 )
		| ( { 9{ U_173 } } & TR_152 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_113_en = ( ST1_03d | U_174 | RG_rl_113_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_113_en )
		RG_rl_113 <= RG_rl_113_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_126 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_151 = TR_126 ;
	7'h01 :
		TR_151 = TR_126 ;
	7'h02 :
		TR_151 = TR_126 ;
	7'h03 :
		TR_151 = TR_126 ;
	7'h04 :
		TR_151 = TR_126 ;
	7'h05 :
		TR_151 = TR_126 ;
	7'h06 :
		TR_151 = TR_126 ;
	7'h07 :
		TR_151 = TR_126 ;
	7'h08 :
		TR_151 = TR_126 ;
	7'h09 :
		TR_151 = TR_126 ;
	7'h0a :
		TR_151 = TR_126 ;
	7'h0b :
		TR_151 = TR_126 ;
	7'h0c :
		TR_151 = TR_126 ;
	7'h0d :
		TR_151 = TR_126 ;
	7'h0e :
		TR_151 = TR_126 ;
	7'h0f :
		TR_151 = TR_126 ;
	7'h10 :
		TR_151 = TR_126 ;
	7'h11 :
		TR_151 = TR_126 ;
	7'h12 :
		TR_151 = TR_126 ;
	7'h13 :
		TR_151 = TR_126 ;
	7'h14 :
		TR_151 = TR_126 ;
	7'h15 :
		TR_151 = TR_126 ;
	7'h16 :
		TR_151 = TR_126 ;
	7'h17 :
		TR_151 = TR_126 ;
	7'h18 :
		TR_151 = TR_126 ;
	7'h19 :
		TR_151 = TR_126 ;
	7'h1a :
		TR_151 = TR_126 ;
	7'h1b :
		TR_151 = TR_126 ;
	7'h1c :
		TR_151 = TR_126 ;
	7'h1d :
		TR_151 = TR_126 ;
	7'h1e :
		TR_151 = TR_126 ;
	7'h1f :
		TR_151 = TR_126 ;
	7'h20 :
		TR_151 = TR_126 ;
	7'h21 :
		TR_151 = TR_126 ;
	7'h22 :
		TR_151 = TR_126 ;
	7'h23 :
		TR_151 = TR_126 ;
	7'h24 :
		TR_151 = TR_126 ;
	7'h25 :
		TR_151 = TR_126 ;
	7'h26 :
		TR_151 = TR_126 ;
	7'h27 :
		TR_151 = TR_126 ;
	7'h28 :
		TR_151 = TR_126 ;
	7'h29 :
		TR_151 = TR_126 ;
	7'h2a :
		TR_151 = TR_126 ;
	7'h2b :
		TR_151 = TR_126 ;
	7'h2c :
		TR_151 = TR_126 ;
	7'h2d :
		TR_151 = TR_126 ;
	7'h2e :
		TR_151 = TR_126 ;
	7'h2f :
		TR_151 = TR_126 ;
	7'h30 :
		TR_151 = TR_126 ;
	7'h31 :
		TR_151 = TR_126 ;
	7'h32 :
		TR_151 = TR_126 ;
	7'h33 :
		TR_151 = TR_126 ;
	7'h34 :
		TR_151 = TR_126 ;
	7'h35 :
		TR_151 = TR_126 ;
	7'h36 :
		TR_151 = TR_126 ;
	7'h37 :
		TR_151 = TR_126 ;
	7'h38 :
		TR_151 = TR_126 ;
	7'h39 :
		TR_151 = TR_126 ;
	7'h3a :
		TR_151 = TR_126 ;
	7'h3b :
		TR_151 = TR_126 ;
	7'h3c :
		TR_151 = TR_126 ;
	7'h3d :
		TR_151 = TR_126 ;
	7'h3e :
		TR_151 = TR_126 ;
	7'h3f :
		TR_151 = TR_126 ;
	7'h40 :
		TR_151 = TR_126 ;
	7'h41 :
		TR_151 = TR_126 ;
	7'h42 :
		TR_151 = TR_126 ;
	7'h43 :
		TR_151 = TR_126 ;
	7'h44 :
		TR_151 = TR_126 ;
	7'h45 :
		TR_151 = TR_126 ;
	7'h46 :
		TR_151 = TR_126 ;
	7'h47 :
		TR_151 = TR_126 ;
	7'h48 :
		TR_151 = TR_126 ;
	7'h49 :
		TR_151 = TR_126 ;
	7'h4a :
		TR_151 = TR_126 ;
	7'h4b :
		TR_151 = TR_126 ;
	7'h4c :
		TR_151 = TR_126 ;
	7'h4d :
		TR_151 = TR_126 ;
	7'h4e :
		TR_151 = TR_126 ;
	7'h4f :
		TR_151 = TR_126 ;
	7'h50 :
		TR_151 = TR_126 ;
	7'h51 :
		TR_151 = TR_126 ;
	7'h52 :
		TR_151 = TR_126 ;
	7'h53 :
		TR_151 = TR_126 ;
	7'h54 :
		TR_151 = TR_126 ;
	7'h55 :
		TR_151 = TR_126 ;
	7'h56 :
		TR_151 = TR_126 ;
	7'h57 :
		TR_151 = TR_126 ;
	7'h58 :
		TR_151 = TR_126 ;
	7'h59 :
		TR_151 = TR_126 ;
	7'h5a :
		TR_151 = TR_126 ;
	7'h5b :
		TR_151 = TR_126 ;
	7'h5c :
		TR_151 = TR_126 ;
	7'h5d :
		TR_151 = TR_126 ;
	7'h5e :
		TR_151 = TR_126 ;
	7'h5f :
		TR_151 = TR_126 ;
	7'h60 :
		TR_151 = TR_126 ;
	7'h61 :
		TR_151 = TR_126 ;
	7'h62 :
		TR_151 = TR_126 ;
	7'h63 :
		TR_151 = TR_126 ;
	7'h64 :
		TR_151 = TR_126 ;
	7'h65 :
		TR_151 = TR_126 ;
	7'h66 :
		TR_151 = TR_126 ;
	7'h67 :
		TR_151 = TR_126 ;
	7'h68 :
		TR_151 = TR_126 ;
	7'h69 :
		TR_151 = TR_126 ;
	7'h6a :
		TR_151 = TR_126 ;
	7'h6b :
		TR_151 = TR_126 ;
	7'h6c :
		TR_151 = TR_126 ;
	7'h6d :
		TR_151 = TR_126 ;
	7'h6e :
		TR_151 = TR_126 ;
	7'h6f :
		TR_151 = TR_126 ;
	7'h70 :
		TR_151 = TR_126 ;
	7'h71 :
		TR_151 = TR_126 ;
	7'h72 :
		TR_151 = 9'h000 ;	// line#=../rle.cpp:80
	7'h73 :
		TR_151 = TR_126 ;
	7'h74 :
		TR_151 = TR_126 ;
	7'h75 :
		TR_151 = TR_126 ;
	7'h76 :
		TR_151 = TR_126 ;
	7'h77 :
		TR_151 = TR_126 ;
	7'h78 :
		TR_151 = TR_126 ;
	7'h79 :
		TR_151 = TR_126 ;
	7'h7a :
		TR_151 = TR_126 ;
	7'h7b :
		TR_151 = TR_126 ;
	7'h7c :
		TR_151 = TR_126 ;
	7'h7d :
		TR_151 = TR_126 ;
	7'h7e :
		TR_151 = TR_126 ;
	7'h7f :
		TR_151 = TR_126 ;
	default :
		TR_151 = 9'hx ;
	endcase
always @ ( TR_151 or U_173 or sub8u_71ot or U_183 or RG_rl_186 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_114_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h72 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_114_t = ( ( { 9{ M_180 } } & RG_rl_186 )
		| ( { 9{ U_173 } } & TR_151 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_114_en = ( M_180 | RG_rl_114_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_114_en )
		RG_rl_114 <= RG_rl_114_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_127 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_150 = TR_127 ;
	7'h01 :
		TR_150 = TR_127 ;
	7'h02 :
		TR_150 = TR_127 ;
	7'h03 :
		TR_150 = TR_127 ;
	7'h04 :
		TR_150 = TR_127 ;
	7'h05 :
		TR_150 = TR_127 ;
	7'h06 :
		TR_150 = TR_127 ;
	7'h07 :
		TR_150 = TR_127 ;
	7'h08 :
		TR_150 = TR_127 ;
	7'h09 :
		TR_150 = TR_127 ;
	7'h0a :
		TR_150 = TR_127 ;
	7'h0b :
		TR_150 = TR_127 ;
	7'h0c :
		TR_150 = TR_127 ;
	7'h0d :
		TR_150 = TR_127 ;
	7'h0e :
		TR_150 = TR_127 ;
	7'h0f :
		TR_150 = TR_127 ;
	7'h10 :
		TR_150 = TR_127 ;
	7'h11 :
		TR_150 = TR_127 ;
	7'h12 :
		TR_150 = TR_127 ;
	7'h13 :
		TR_150 = TR_127 ;
	7'h14 :
		TR_150 = TR_127 ;
	7'h15 :
		TR_150 = TR_127 ;
	7'h16 :
		TR_150 = TR_127 ;
	7'h17 :
		TR_150 = TR_127 ;
	7'h18 :
		TR_150 = TR_127 ;
	7'h19 :
		TR_150 = TR_127 ;
	7'h1a :
		TR_150 = TR_127 ;
	7'h1b :
		TR_150 = TR_127 ;
	7'h1c :
		TR_150 = TR_127 ;
	7'h1d :
		TR_150 = TR_127 ;
	7'h1e :
		TR_150 = TR_127 ;
	7'h1f :
		TR_150 = TR_127 ;
	7'h20 :
		TR_150 = TR_127 ;
	7'h21 :
		TR_150 = TR_127 ;
	7'h22 :
		TR_150 = TR_127 ;
	7'h23 :
		TR_150 = TR_127 ;
	7'h24 :
		TR_150 = TR_127 ;
	7'h25 :
		TR_150 = TR_127 ;
	7'h26 :
		TR_150 = TR_127 ;
	7'h27 :
		TR_150 = TR_127 ;
	7'h28 :
		TR_150 = TR_127 ;
	7'h29 :
		TR_150 = TR_127 ;
	7'h2a :
		TR_150 = TR_127 ;
	7'h2b :
		TR_150 = TR_127 ;
	7'h2c :
		TR_150 = TR_127 ;
	7'h2d :
		TR_150 = TR_127 ;
	7'h2e :
		TR_150 = TR_127 ;
	7'h2f :
		TR_150 = TR_127 ;
	7'h30 :
		TR_150 = TR_127 ;
	7'h31 :
		TR_150 = TR_127 ;
	7'h32 :
		TR_150 = TR_127 ;
	7'h33 :
		TR_150 = TR_127 ;
	7'h34 :
		TR_150 = TR_127 ;
	7'h35 :
		TR_150 = TR_127 ;
	7'h36 :
		TR_150 = TR_127 ;
	7'h37 :
		TR_150 = TR_127 ;
	7'h38 :
		TR_150 = TR_127 ;
	7'h39 :
		TR_150 = TR_127 ;
	7'h3a :
		TR_150 = TR_127 ;
	7'h3b :
		TR_150 = TR_127 ;
	7'h3c :
		TR_150 = TR_127 ;
	7'h3d :
		TR_150 = TR_127 ;
	7'h3e :
		TR_150 = TR_127 ;
	7'h3f :
		TR_150 = TR_127 ;
	7'h40 :
		TR_150 = TR_127 ;
	7'h41 :
		TR_150 = TR_127 ;
	7'h42 :
		TR_150 = TR_127 ;
	7'h43 :
		TR_150 = TR_127 ;
	7'h44 :
		TR_150 = TR_127 ;
	7'h45 :
		TR_150 = TR_127 ;
	7'h46 :
		TR_150 = TR_127 ;
	7'h47 :
		TR_150 = TR_127 ;
	7'h48 :
		TR_150 = TR_127 ;
	7'h49 :
		TR_150 = TR_127 ;
	7'h4a :
		TR_150 = TR_127 ;
	7'h4b :
		TR_150 = TR_127 ;
	7'h4c :
		TR_150 = TR_127 ;
	7'h4d :
		TR_150 = TR_127 ;
	7'h4e :
		TR_150 = TR_127 ;
	7'h4f :
		TR_150 = TR_127 ;
	7'h50 :
		TR_150 = TR_127 ;
	7'h51 :
		TR_150 = TR_127 ;
	7'h52 :
		TR_150 = TR_127 ;
	7'h53 :
		TR_150 = TR_127 ;
	7'h54 :
		TR_150 = TR_127 ;
	7'h55 :
		TR_150 = TR_127 ;
	7'h56 :
		TR_150 = TR_127 ;
	7'h57 :
		TR_150 = TR_127 ;
	7'h58 :
		TR_150 = TR_127 ;
	7'h59 :
		TR_150 = TR_127 ;
	7'h5a :
		TR_150 = TR_127 ;
	7'h5b :
		TR_150 = TR_127 ;
	7'h5c :
		TR_150 = TR_127 ;
	7'h5d :
		TR_150 = TR_127 ;
	7'h5e :
		TR_150 = TR_127 ;
	7'h5f :
		TR_150 = TR_127 ;
	7'h60 :
		TR_150 = TR_127 ;
	7'h61 :
		TR_150 = TR_127 ;
	7'h62 :
		TR_150 = TR_127 ;
	7'h63 :
		TR_150 = TR_127 ;
	7'h64 :
		TR_150 = TR_127 ;
	7'h65 :
		TR_150 = TR_127 ;
	7'h66 :
		TR_150 = TR_127 ;
	7'h67 :
		TR_150 = TR_127 ;
	7'h68 :
		TR_150 = TR_127 ;
	7'h69 :
		TR_150 = TR_127 ;
	7'h6a :
		TR_150 = TR_127 ;
	7'h6b :
		TR_150 = TR_127 ;
	7'h6c :
		TR_150 = TR_127 ;
	7'h6d :
		TR_150 = TR_127 ;
	7'h6e :
		TR_150 = TR_127 ;
	7'h6f :
		TR_150 = TR_127 ;
	7'h70 :
		TR_150 = TR_127 ;
	7'h71 :
		TR_150 = TR_127 ;
	7'h72 :
		TR_150 = TR_127 ;
	7'h73 :
		TR_150 = 9'h000 ;	// line#=../rle.cpp:80
	7'h74 :
		TR_150 = TR_127 ;
	7'h75 :
		TR_150 = TR_127 ;
	7'h76 :
		TR_150 = TR_127 ;
	7'h77 :
		TR_150 = TR_127 ;
	7'h78 :
		TR_150 = TR_127 ;
	7'h79 :
		TR_150 = TR_127 ;
	7'h7a :
		TR_150 = TR_127 ;
	7'h7b :
		TR_150 = TR_127 ;
	7'h7c :
		TR_150 = TR_127 ;
	7'h7d :
		TR_150 = TR_127 ;
	7'h7e :
		TR_150 = TR_127 ;
	7'h7f :
		TR_150 = TR_127 ;
	default :
		TR_150 = 9'hx ;
	endcase
always @ ( TR_150 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_55 or 
	U_174 or RG_rl_186 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_115_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h73 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_115_t = ( ( { 9{ ST1_03d } } & RG_rl_186 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_55 )
		| ( { 9{ U_173 } } & TR_150 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_115_en = ( ST1_03d | U_174 | RG_rl_115_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_115_en )
		RG_rl_115 <= RG_rl_115_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_128 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_149 = TR_128 ;
	7'h01 :
		TR_149 = TR_128 ;
	7'h02 :
		TR_149 = TR_128 ;
	7'h03 :
		TR_149 = TR_128 ;
	7'h04 :
		TR_149 = TR_128 ;
	7'h05 :
		TR_149 = TR_128 ;
	7'h06 :
		TR_149 = TR_128 ;
	7'h07 :
		TR_149 = TR_128 ;
	7'h08 :
		TR_149 = TR_128 ;
	7'h09 :
		TR_149 = TR_128 ;
	7'h0a :
		TR_149 = TR_128 ;
	7'h0b :
		TR_149 = TR_128 ;
	7'h0c :
		TR_149 = TR_128 ;
	7'h0d :
		TR_149 = TR_128 ;
	7'h0e :
		TR_149 = TR_128 ;
	7'h0f :
		TR_149 = TR_128 ;
	7'h10 :
		TR_149 = TR_128 ;
	7'h11 :
		TR_149 = TR_128 ;
	7'h12 :
		TR_149 = TR_128 ;
	7'h13 :
		TR_149 = TR_128 ;
	7'h14 :
		TR_149 = TR_128 ;
	7'h15 :
		TR_149 = TR_128 ;
	7'h16 :
		TR_149 = TR_128 ;
	7'h17 :
		TR_149 = TR_128 ;
	7'h18 :
		TR_149 = TR_128 ;
	7'h19 :
		TR_149 = TR_128 ;
	7'h1a :
		TR_149 = TR_128 ;
	7'h1b :
		TR_149 = TR_128 ;
	7'h1c :
		TR_149 = TR_128 ;
	7'h1d :
		TR_149 = TR_128 ;
	7'h1e :
		TR_149 = TR_128 ;
	7'h1f :
		TR_149 = TR_128 ;
	7'h20 :
		TR_149 = TR_128 ;
	7'h21 :
		TR_149 = TR_128 ;
	7'h22 :
		TR_149 = TR_128 ;
	7'h23 :
		TR_149 = TR_128 ;
	7'h24 :
		TR_149 = TR_128 ;
	7'h25 :
		TR_149 = TR_128 ;
	7'h26 :
		TR_149 = TR_128 ;
	7'h27 :
		TR_149 = TR_128 ;
	7'h28 :
		TR_149 = TR_128 ;
	7'h29 :
		TR_149 = TR_128 ;
	7'h2a :
		TR_149 = TR_128 ;
	7'h2b :
		TR_149 = TR_128 ;
	7'h2c :
		TR_149 = TR_128 ;
	7'h2d :
		TR_149 = TR_128 ;
	7'h2e :
		TR_149 = TR_128 ;
	7'h2f :
		TR_149 = TR_128 ;
	7'h30 :
		TR_149 = TR_128 ;
	7'h31 :
		TR_149 = TR_128 ;
	7'h32 :
		TR_149 = TR_128 ;
	7'h33 :
		TR_149 = TR_128 ;
	7'h34 :
		TR_149 = TR_128 ;
	7'h35 :
		TR_149 = TR_128 ;
	7'h36 :
		TR_149 = TR_128 ;
	7'h37 :
		TR_149 = TR_128 ;
	7'h38 :
		TR_149 = TR_128 ;
	7'h39 :
		TR_149 = TR_128 ;
	7'h3a :
		TR_149 = TR_128 ;
	7'h3b :
		TR_149 = TR_128 ;
	7'h3c :
		TR_149 = TR_128 ;
	7'h3d :
		TR_149 = TR_128 ;
	7'h3e :
		TR_149 = TR_128 ;
	7'h3f :
		TR_149 = TR_128 ;
	7'h40 :
		TR_149 = TR_128 ;
	7'h41 :
		TR_149 = TR_128 ;
	7'h42 :
		TR_149 = TR_128 ;
	7'h43 :
		TR_149 = TR_128 ;
	7'h44 :
		TR_149 = TR_128 ;
	7'h45 :
		TR_149 = TR_128 ;
	7'h46 :
		TR_149 = TR_128 ;
	7'h47 :
		TR_149 = TR_128 ;
	7'h48 :
		TR_149 = TR_128 ;
	7'h49 :
		TR_149 = TR_128 ;
	7'h4a :
		TR_149 = TR_128 ;
	7'h4b :
		TR_149 = TR_128 ;
	7'h4c :
		TR_149 = TR_128 ;
	7'h4d :
		TR_149 = TR_128 ;
	7'h4e :
		TR_149 = TR_128 ;
	7'h4f :
		TR_149 = TR_128 ;
	7'h50 :
		TR_149 = TR_128 ;
	7'h51 :
		TR_149 = TR_128 ;
	7'h52 :
		TR_149 = TR_128 ;
	7'h53 :
		TR_149 = TR_128 ;
	7'h54 :
		TR_149 = TR_128 ;
	7'h55 :
		TR_149 = TR_128 ;
	7'h56 :
		TR_149 = TR_128 ;
	7'h57 :
		TR_149 = TR_128 ;
	7'h58 :
		TR_149 = TR_128 ;
	7'h59 :
		TR_149 = TR_128 ;
	7'h5a :
		TR_149 = TR_128 ;
	7'h5b :
		TR_149 = TR_128 ;
	7'h5c :
		TR_149 = TR_128 ;
	7'h5d :
		TR_149 = TR_128 ;
	7'h5e :
		TR_149 = TR_128 ;
	7'h5f :
		TR_149 = TR_128 ;
	7'h60 :
		TR_149 = TR_128 ;
	7'h61 :
		TR_149 = TR_128 ;
	7'h62 :
		TR_149 = TR_128 ;
	7'h63 :
		TR_149 = TR_128 ;
	7'h64 :
		TR_149 = TR_128 ;
	7'h65 :
		TR_149 = TR_128 ;
	7'h66 :
		TR_149 = TR_128 ;
	7'h67 :
		TR_149 = TR_128 ;
	7'h68 :
		TR_149 = TR_128 ;
	7'h69 :
		TR_149 = TR_128 ;
	7'h6a :
		TR_149 = TR_128 ;
	7'h6b :
		TR_149 = TR_128 ;
	7'h6c :
		TR_149 = TR_128 ;
	7'h6d :
		TR_149 = TR_128 ;
	7'h6e :
		TR_149 = TR_128 ;
	7'h6f :
		TR_149 = TR_128 ;
	7'h70 :
		TR_149 = TR_128 ;
	7'h71 :
		TR_149 = TR_128 ;
	7'h72 :
		TR_149 = TR_128 ;
	7'h73 :
		TR_149 = TR_128 ;
	7'h74 :
		TR_149 = 9'h000 ;	// line#=../rle.cpp:80
	7'h75 :
		TR_149 = TR_128 ;
	7'h76 :
		TR_149 = TR_128 ;
	7'h77 :
		TR_149 = TR_128 ;
	7'h78 :
		TR_149 = TR_128 ;
	7'h79 :
		TR_149 = TR_128 ;
	7'h7a :
		TR_149 = TR_128 ;
	7'h7b :
		TR_149 = TR_128 ;
	7'h7c :
		TR_149 = TR_128 ;
	7'h7d :
		TR_149 = TR_128 ;
	7'h7e :
		TR_149 = TR_128 ;
	7'h7f :
		TR_149 = TR_128 ;
	default :
		TR_149 = 9'hx ;
	endcase
always @ ( TR_149 or U_173 or sub8u_71ot or U_183 or RG_rl_187 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_116_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h74 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_116_t = ( ( { 9{ M_180 } } & RG_rl_187 )
		| ( { 9{ U_173 } } & TR_149 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_116_en = ( M_180 | RG_rl_116_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_116_en )
		RG_rl_116 <= RG_rl_116_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_129 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_148 = TR_129 ;
	7'h01 :
		TR_148 = TR_129 ;
	7'h02 :
		TR_148 = TR_129 ;
	7'h03 :
		TR_148 = TR_129 ;
	7'h04 :
		TR_148 = TR_129 ;
	7'h05 :
		TR_148 = TR_129 ;
	7'h06 :
		TR_148 = TR_129 ;
	7'h07 :
		TR_148 = TR_129 ;
	7'h08 :
		TR_148 = TR_129 ;
	7'h09 :
		TR_148 = TR_129 ;
	7'h0a :
		TR_148 = TR_129 ;
	7'h0b :
		TR_148 = TR_129 ;
	7'h0c :
		TR_148 = TR_129 ;
	7'h0d :
		TR_148 = TR_129 ;
	7'h0e :
		TR_148 = TR_129 ;
	7'h0f :
		TR_148 = TR_129 ;
	7'h10 :
		TR_148 = TR_129 ;
	7'h11 :
		TR_148 = TR_129 ;
	7'h12 :
		TR_148 = TR_129 ;
	7'h13 :
		TR_148 = TR_129 ;
	7'h14 :
		TR_148 = TR_129 ;
	7'h15 :
		TR_148 = TR_129 ;
	7'h16 :
		TR_148 = TR_129 ;
	7'h17 :
		TR_148 = TR_129 ;
	7'h18 :
		TR_148 = TR_129 ;
	7'h19 :
		TR_148 = TR_129 ;
	7'h1a :
		TR_148 = TR_129 ;
	7'h1b :
		TR_148 = TR_129 ;
	7'h1c :
		TR_148 = TR_129 ;
	7'h1d :
		TR_148 = TR_129 ;
	7'h1e :
		TR_148 = TR_129 ;
	7'h1f :
		TR_148 = TR_129 ;
	7'h20 :
		TR_148 = TR_129 ;
	7'h21 :
		TR_148 = TR_129 ;
	7'h22 :
		TR_148 = TR_129 ;
	7'h23 :
		TR_148 = TR_129 ;
	7'h24 :
		TR_148 = TR_129 ;
	7'h25 :
		TR_148 = TR_129 ;
	7'h26 :
		TR_148 = TR_129 ;
	7'h27 :
		TR_148 = TR_129 ;
	7'h28 :
		TR_148 = TR_129 ;
	7'h29 :
		TR_148 = TR_129 ;
	7'h2a :
		TR_148 = TR_129 ;
	7'h2b :
		TR_148 = TR_129 ;
	7'h2c :
		TR_148 = TR_129 ;
	7'h2d :
		TR_148 = TR_129 ;
	7'h2e :
		TR_148 = TR_129 ;
	7'h2f :
		TR_148 = TR_129 ;
	7'h30 :
		TR_148 = TR_129 ;
	7'h31 :
		TR_148 = TR_129 ;
	7'h32 :
		TR_148 = TR_129 ;
	7'h33 :
		TR_148 = TR_129 ;
	7'h34 :
		TR_148 = TR_129 ;
	7'h35 :
		TR_148 = TR_129 ;
	7'h36 :
		TR_148 = TR_129 ;
	7'h37 :
		TR_148 = TR_129 ;
	7'h38 :
		TR_148 = TR_129 ;
	7'h39 :
		TR_148 = TR_129 ;
	7'h3a :
		TR_148 = TR_129 ;
	7'h3b :
		TR_148 = TR_129 ;
	7'h3c :
		TR_148 = TR_129 ;
	7'h3d :
		TR_148 = TR_129 ;
	7'h3e :
		TR_148 = TR_129 ;
	7'h3f :
		TR_148 = TR_129 ;
	7'h40 :
		TR_148 = TR_129 ;
	7'h41 :
		TR_148 = TR_129 ;
	7'h42 :
		TR_148 = TR_129 ;
	7'h43 :
		TR_148 = TR_129 ;
	7'h44 :
		TR_148 = TR_129 ;
	7'h45 :
		TR_148 = TR_129 ;
	7'h46 :
		TR_148 = TR_129 ;
	7'h47 :
		TR_148 = TR_129 ;
	7'h48 :
		TR_148 = TR_129 ;
	7'h49 :
		TR_148 = TR_129 ;
	7'h4a :
		TR_148 = TR_129 ;
	7'h4b :
		TR_148 = TR_129 ;
	7'h4c :
		TR_148 = TR_129 ;
	7'h4d :
		TR_148 = TR_129 ;
	7'h4e :
		TR_148 = TR_129 ;
	7'h4f :
		TR_148 = TR_129 ;
	7'h50 :
		TR_148 = TR_129 ;
	7'h51 :
		TR_148 = TR_129 ;
	7'h52 :
		TR_148 = TR_129 ;
	7'h53 :
		TR_148 = TR_129 ;
	7'h54 :
		TR_148 = TR_129 ;
	7'h55 :
		TR_148 = TR_129 ;
	7'h56 :
		TR_148 = TR_129 ;
	7'h57 :
		TR_148 = TR_129 ;
	7'h58 :
		TR_148 = TR_129 ;
	7'h59 :
		TR_148 = TR_129 ;
	7'h5a :
		TR_148 = TR_129 ;
	7'h5b :
		TR_148 = TR_129 ;
	7'h5c :
		TR_148 = TR_129 ;
	7'h5d :
		TR_148 = TR_129 ;
	7'h5e :
		TR_148 = TR_129 ;
	7'h5f :
		TR_148 = TR_129 ;
	7'h60 :
		TR_148 = TR_129 ;
	7'h61 :
		TR_148 = TR_129 ;
	7'h62 :
		TR_148 = TR_129 ;
	7'h63 :
		TR_148 = TR_129 ;
	7'h64 :
		TR_148 = TR_129 ;
	7'h65 :
		TR_148 = TR_129 ;
	7'h66 :
		TR_148 = TR_129 ;
	7'h67 :
		TR_148 = TR_129 ;
	7'h68 :
		TR_148 = TR_129 ;
	7'h69 :
		TR_148 = TR_129 ;
	7'h6a :
		TR_148 = TR_129 ;
	7'h6b :
		TR_148 = TR_129 ;
	7'h6c :
		TR_148 = TR_129 ;
	7'h6d :
		TR_148 = TR_129 ;
	7'h6e :
		TR_148 = TR_129 ;
	7'h6f :
		TR_148 = TR_129 ;
	7'h70 :
		TR_148 = TR_129 ;
	7'h71 :
		TR_148 = TR_129 ;
	7'h72 :
		TR_148 = TR_129 ;
	7'h73 :
		TR_148 = TR_129 ;
	7'h74 :
		TR_148 = TR_129 ;
	7'h75 :
		TR_148 = 9'h000 ;	// line#=../rle.cpp:80
	7'h76 :
		TR_148 = TR_129 ;
	7'h77 :
		TR_148 = TR_129 ;
	7'h78 :
		TR_148 = TR_129 ;
	7'h79 :
		TR_148 = TR_129 ;
	7'h7a :
		TR_148 = TR_129 ;
	7'h7b :
		TR_148 = TR_129 ;
	7'h7c :
		TR_148 = TR_129 ;
	7'h7d :
		TR_148 = TR_129 ;
	7'h7e :
		TR_148 = TR_129 ;
	7'h7f :
		TR_148 = TR_129 ;
	default :
		TR_148 = 9'hx ;
	endcase
always @ ( TR_148 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_56 or 
	U_174 or RG_rl_187 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_117_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h75 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_117_t = ( ( { 9{ ST1_03d } } & RG_rl_187 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_56 )
		| ( { 9{ U_173 } } & TR_148 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_117_en = ( ST1_03d | U_174 | RG_rl_117_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_117_en )
		RG_rl_117 <= RG_rl_117_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_130 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_147 = TR_130 ;
	7'h01 :
		TR_147 = TR_130 ;
	7'h02 :
		TR_147 = TR_130 ;
	7'h03 :
		TR_147 = TR_130 ;
	7'h04 :
		TR_147 = TR_130 ;
	7'h05 :
		TR_147 = TR_130 ;
	7'h06 :
		TR_147 = TR_130 ;
	7'h07 :
		TR_147 = TR_130 ;
	7'h08 :
		TR_147 = TR_130 ;
	7'h09 :
		TR_147 = TR_130 ;
	7'h0a :
		TR_147 = TR_130 ;
	7'h0b :
		TR_147 = TR_130 ;
	7'h0c :
		TR_147 = TR_130 ;
	7'h0d :
		TR_147 = TR_130 ;
	7'h0e :
		TR_147 = TR_130 ;
	7'h0f :
		TR_147 = TR_130 ;
	7'h10 :
		TR_147 = TR_130 ;
	7'h11 :
		TR_147 = TR_130 ;
	7'h12 :
		TR_147 = TR_130 ;
	7'h13 :
		TR_147 = TR_130 ;
	7'h14 :
		TR_147 = TR_130 ;
	7'h15 :
		TR_147 = TR_130 ;
	7'h16 :
		TR_147 = TR_130 ;
	7'h17 :
		TR_147 = TR_130 ;
	7'h18 :
		TR_147 = TR_130 ;
	7'h19 :
		TR_147 = TR_130 ;
	7'h1a :
		TR_147 = TR_130 ;
	7'h1b :
		TR_147 = TR_130 ;
	7'h1c :
		TR_147 = TR_130 ;
	7'h1d :
		TR_147 = TR_130 ;
	7'h1e :
		TR_147 = TR_130 ;
	7'h1f :
		TR_147 = TR_130 ;
	7'h20 :
		TR_147 = TR_130 ;
	7'h21 :
		TR_147 = TR_130 ;
	7'h22 :
		TR_147 = TR_130 ;
	7'h23 :
		TR_147 = TR_130 ;
	7'h24 :
		TR_147 = TR_130 ;
	7'h25 :
		TR_147 = TR_130 ;
	7'h26 :
		TR_147 = TR_130 ;
	7'h27 :
		TR_147 = TR_130 ;
	7'h28 :
		TR_147 = TR_130 ;
	7'h29 :
		TR_147 = TR_130 ;
	7'h2a :
		TR_147 = TR_130 ;
	7'h2b :
		TR_147 = TR_130 ;
	7'h2c :
		TR_147 = TR_130 ;
	7'h2d :
		TR_147 = TR_130 ;
	7'h2e :
		TR_147 = TR_130 ;
	7'h2f :
		TR_147 = TR_130 ;
	7'h30 :
		TR_147 = TR_130 ;
	7'h31 :
		TR_147 = TR_130 ;
	7'h32 :
		TR_147 = TR_130 ;
	7'h33 :
		TR_147 = TR_130 ;
	7'h34 :
		TR_147 = TR_130 ;
	7'h35 :
		TR_147 = TR_130 ;
	7'h36 :
		TR_147 = TR_130 ;
	7'h37 :
		TR_147 = TR_130 ;
	7'h38 :
		TR_147 = TR_130 ;
	7'h39 :
		TR_147 = TR_130 ;
	7'h3a :
		TR_147 = TR_130 ;
	7'h3b :
		TR_147 = TR_130 ;
	7'h3c :
		TR_147 = TR_130 ;
	7'h3d :
		TR_147 = TR_130 ;
	7'h3e :
		TR_147 = TR_130 ;
	7'h3f :
		TR_147 = TR_130 ;
	7'h40 :
		TR_147 = TR_130 ;
	7'h41 :
		TR_147 = TR_130 ;
	7'h42 :
		TR_147 = TR_130 ;
	7'h43 :
		TR_147 = TR_130 ;
	7'h44 :
		TR_147 = TR_130 ;
	7'h45 :
		TR_147 = TR_130 ;
	7'h46 :
		TR_147 = TR_130 ;
	7'h47 :
		TR_147 = TR_130 ;
	7'h48 :
		TR_147 = TR_130 ;
	7'h49 :
		TR_147 = TR_130 ;
	7'h4a :
		TR_147 = TR_130 ;
	7'h4b :
		TR_147 = TR_130 ;
	7'h4c :
		TR_147 = TR_130 ;
	7'h4d :
		TR_147 = TR_130 ;
	7'h4e :
		TR_147 = TR_130 ;
	7'h4f :
		TR_147 = TR_130 ;
	7'h50 :
		TR_147 = TR_130 ;
	7'h51 :
		TR_147 = TR_130 ;
	7'h52 :
		TR_147 = TR_130 ;
	7'h53 :
		TR_147 = TR_130 ;
	7'h54 :
		TR_147 = TR_130 ;
	7'h55 :
		TR_147 = TR_130 ;
	7'h56 :
		TR_147 = TR_130 ;
	7'h57 :
		TR_147 = TR_130 ;
	7'h58 :
		TR_147 = TR_130 ;
	7'h59 :
		TR_147 = TR_130 ;
	7'h5a :
		TR_147 = TR_130 ;
	7'h5b :
		TR_147 = TR_130 ;
	7'h5c :
		TR_147 = TR_130 ;
	7'h5d :
		TR_147 = TR_130 ;
	7'h5e :
		TR_147 = TR_130 ;
	7'h5f :
		TR_147 = TR_130 ;
	7'h60 :
		TR_147 = TR_130 ;
	7'h61 :
		TR_147 = TR_130 ;
	7'h62 :
		TR_147 = TR_130 ;
	7'h63 :
		TR_147 = TR_130 ;
	7'h64 :
		TR_147 = TR_130 ;
	7'h65 :
		TR_147 = TR_130 ;
	7'h66 :
		TR_147 = TR_130 ;
	7'h67 :
		TR_147 = TR_130 ;
	7'h68 :
		TR_147 = TR_130 ;
	7'h69 :
		TR_147 = TR_130 ;
	7'h6a :
		TR_147 = TR_130 ;
	7'h6b :
		TR_147 = TR_130 ;
	7'h6c :
		TR_147 = TR_130 ;
	7'h6d :
		TR_147 = TR_130 ;
	7'h6e :
		TR_147 = TR_130 ;
	7'h6f :
		TR_147 = TR_130 ;
	7'h70 :
		TR_147 = TR_130 ;
	7'h71 :
		TR_147 = TR_130 ;
	7'h72 :
		TR_147 = TR_130 ;
	7'h73 :
		TR_147 = TR_130 ;
	7'h74 :
		TR_147 = TR_130 ;
	7'h75 :
		TR_147 = TR_130 ;
	7'h76 :
		TR_147 = 9'h000 ;	// line#=../rle.cpp:80
	7'h77 :
		TR_147 = TR_130 ;
	7'h78 :
		TR_147 = TR_130 ;
	7'h79 :
		TR_147 = TR_130 ;
	7'h7a :
		TR_147 = TR_130 ;
	7'h7b :
		TR_147 = TR_130 ;
	7'h7c :
		TR_147 = TR_130 ;
	7'h7d :
		TR_147 = TR_130 ;
	7'h7e :
		TR_147 = TR_130 ;
	7'h7f :
		TR_147 = TR_130 ;
	default :
		TR_147 = 9'hx ;
	endcase
always @ ( TR_147 or U_173 or sub8u_71ot or U_183 or RG_rl_188 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_118_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h76 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_118_t = ( ( { 9{ M_180 } } & RG_rl_188 )
		| ( { 9{ U_173 } } & TR_147 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_118_en = ( M_180 | RG_rl_118_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_118_en )
		RG_rl_118 <= RG_rl_118_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_131 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_146 = TR_131 ;
	7'h01 :
		TR_146 = TR_131 ;
	7'h02 :
		TR_146 = TR_131 ;
	7'h03 :
		TR_146 = TR_131 ;
	7'h04 :
		TR_146 = TR_131 ;
	7'h05 :
		TR_146 = TR_131 ;
	7'h06 :
		TR_146 = TR_131 ;
	7'h07 :
		TR_146 = TR_131 ;
	7'h08 :
		TR_146 = TR_131 ;
	7'h09 :
		TR_146 = TR_131 ;
	7'h0a :
		TR_146 = TR_131 ;
	7'h0b :
		TR_146 = TR_131 ;
	7'h0c :
		TR_146 = TR_131 ;
	7'h0d :
		TR_146 = TR_131 ;
	7'h0e :
		TR_146 = TR_131 ;
	7'h0f :
		TR_146 = TR_131 ;
	7'h10 :
		TR_146 = TR_131 ;
	7'h11 :
		TR_146 = TR_131 ;
	7'h12 :
		TR_146 = TR_131 ;
	7'h13 :
		TR_146 = TR_131 ;
	7'h14 :
		TR_146 = TR_131 ;
	7'h15 :
		TR_146 = TR_131 ;
	7'h16 :
		TR_146 = TR_131 ;
	7'h17 :
		TR_146 = TR_131 ;
	7'h18 :
		TR_146 = TR_131 ;
	7'h19 :
		TR_146 = TR_131 ;
	7'h1a :
		TR_146 = TR_131 ;
	7'h1b :
		TR_146 = TR_131 ;
	7'h1c :
		TR_146 = TR_131 ;
	7'h1d :
		TR_146 = TR_131 ;
	7'h1e :
		TR_146 = TR_131 ;
	7'h1f :
		TR_146 = TR_131 ;
	7'h20 :
		TR_146 = TR_131 ;
	7'h21 :
		TR_146 = TR_131 ;
	7'h22 :
		TR_146 = TR_131 ;
	7'h23 :
		TR_146 = TR_131 ;
	7'h24 :
		TR_146 = TR_131 ;
	7'h25 :
		TR_146 = TR_131 ;
	7'h26 :
		TR_146 = TR_131 ;
	7'h27 :
		TR_146 = TR_131 ;
	7'h28 :
		TR_146 = TR_131 ;
	7'h29 :
		TR_146 = TR_131 ;
	7'h2a :
		TR_146 = TR_131 ;
	7'h2b :
		TR_146 = TR_131 ;
	7'h2c :
		TR_146 = TR_131 ;
	7'h2d :
		TR_146 = TR_131 ;
	7'h2e :
		TR_146 = TR_131 ;
	7'h2f :
		TR_146 = TR_131 ;
	7'h30 :
		TR_146 = TR_131 ;
	7'h31 :
		TR_146 = TR_131 ;
	7'h32 :
		TR_146 = TR_131 ;
	7'h33 :
		TR_146 = TR_131 ;
	7'h34 :
		TR_146 = TR_131 ;
	7'h35 :
		TR_146 = TR_131 ;
	7'h36 :
		TR_146 = TR_131 ;
	7'h37 :
		TR_146 = TR_131 ;
	7'h38 :
		TR_146 = TR_131 ;
	7'h39 :
		TR_146 = TR_131 ;
	7'h3a :
		TR_146 = TR_131 ;
	7'h3b :
		TR_146 = TR_131 ;
	7'h3c :
		TR_146 = TR_131 ;
	7'h3d :
		TR_146 = TR_131 ;
	7'h3e :
		TR_146 = TR_131 ;
	7'h3f :
		TR_146 = TR_131 ;
	7'h40 :
		TR_146 = TR_131 ;
	7'h41 :
		TR_146 = TR_131 ;
	7'h42 :
		TR_146 = TR_131 ;
	7'h43 :
		TR_146 = TR_131 ;
	7'h44 :
		TR_146 = TR_131 ;
	7'h45 :
		TR_146 = TR_131 ;
	7'h46 :
		TR_146 = TR_131 ;
	7'h47 :
		TR_146 = TR_131 ;
	7'h48 :
		TR_146 = TR_131 ;
	7'h49 :
		TR_146 = TR_131 ;
	7'h4a :
		TR_146 = TR_131 ;
	7'h4b :
		TR_146 = TR_131 ;
	7'h4c :
		TR_146 = TR_131 ;
	7'h4d :
		TR_146 = TR_131 ;
	7'h4e :
		TR_146 = TR_131 ;
	7'h4f :
		TR_146 = TR_131 ;
	7'h50 :
		TR_146 = TR_131 ;
	7'h51 :
		TR_146 = TR_131 ;
	7'h52 :
		TR_146 = TR_131 ;
	7'h53 :
		TR_146 = TR_131 ;
	7'h54 :
		TR_146 = TR_131 ;
	7'h55 :
		TR_146 = TR_131 ;
	7'h56 :
		TR_146 = TR_131 ;
	7'h57 :
		TR_146 = TR_131 ;
	7'h58 :
		TR_146 = TR_131 ;
	7'h59 :
		TR_146 = TR_131 ;
	7'h5a :
		TR_146 = TR_131 ;
	7'h5b :
		TR_146 = TR_131 ;
	7'h5c :
		TR_146 = TR_131 ;
	7'h5d :
		TR_146 = TR_131 ;
	7'h5e :
		TR_146 = TR_131 ;
	7'h5f :
		TR_146 = TR_131 ;
	7'h60 :
		TR_146 = TR_131 ;
	7'h61 :
		TR_146 = TR_131 ;
	7'h62 :
		TR_146 = TR_131 ;
	7'h63 :
		TR_146 = TR_131 ;
	7'h64 :
		TR_146 = TR_131 ;
	7'h65 :
		TR_146 = TR_131 ;
	7'h66 :
		TR_146 = TR_131 ;
	7'h67 :
		TR_146 = TR_131 ;
	7'h68 :
		TR_146 = TR_131 ;
	7'h69 :
		TR_146 = TR_131 ;
	7'h6a :
		TR_146 = TR_131 ;
	7'h6b :
		TR_146 = TR_131 ;
	7'h6c :
		TR_146 = TR_131 ;
	7'h6d :
		TR_146 = TR_131 ;
	7'h6e :
		TR_146 = TR_131 ;
	7'h6f :
		TR_146 = TR_131 ;
	7'h70 :
		TR_146 = TR_131 ;
	7'h71 :
		TR_146 = TR_131 ;
	7'h72 :
		TR_146 = TR_131 ;
	7'h73 :
		TR_146 = TR_131 ;
	7'h74 :
		TR_146 = TR_131 ;
	7'h75 :
		TR_146 = TR_131 ;
	7'h76 :
		TR_146 = TR_131 ;
	7'h77 :
		TR_146 = 9'h000 ;	// line#=../rle.cpp:80
	7'h78 :
		TR_146 = TR_131 ;
	7'h79 :
		TR_146 = TR_131 ;
	7'h7a :
		TR_146 = TR_131 ;
	7'h7b :
		TR_146 = TR_131 ;
	7'h7c :
		TR_146 = TR_131 ;
	7'h7d :
		TR_146 = TR_131 ;
	7'h7e :
		TR_146 = TR_131 ;
	7'h7f :
		TR_146 = TR_131 ;
	default :
		TR_146 = 9'hx ;
	endcase
always @ ( TR_146 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_57 or 
	U_174 or RG_rl_188 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_119_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h77 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_119_t = ( ( { 9{ ST1_03d } } & RG_rl_188 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_57 )
		| ( { 9{ U_173 } } & TR_146 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_119_en = ( ST1_03d | U_174 | RG_rl_119_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_119_en )
		RG_rl_119 <= RG_rl_119_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_132 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_145 = TR_132 ;
	7'h01 :
		TR_145 = TR_132 ;
	7'h02 :
		TR_145 = TR_132 ;
	7'h03 :
		TR_145 = TR_132 ;
	7'h04 :
		TR_145 = TR_132 ;
	7'h05 :
		TR_145 = TR_132 ;
	7'h06 :
		TR_145 = TR_132 ;
	7'h07 :
		TR_145 = TR_132 ;
	7'h08 :
		TR_145 = TR_132 ;
	7'h09 :
		TR_145 = TR_132 ;
	7'h0a :
		TR_145 = TR_132 ;
	7'h0b :
		TR_145 = TR_132 ;
	7'h0c :
		TR_145 = TR_132 ;
	7'h0d :
		TR_145 = TR_132 ;
	7'h0e :
		TR_145 = TR_132 ;
	7'h0f :
		TR_145 = TR_132 ;
	7'h10 :
		TR_145 = TR_132 ;
	7'h11 :
		TR_145 = TR_132 ;
	7'h12 :
		TR_145 = TR_132 ;
	7'h13 :
		TR_145 = TR_132 ;
	7'h14 :
		TR_145 = TR_132 ;
	7'h15 :
		TR_145 = TR_132 ;
	7'h16 :
		TR_145 = TR_132 ;
	7'h17 :
		TR_145 = TR_132 ;
	7'h18 :
		TR_145 = TR_132 ;
	7'h19 :
		TR_145 = TR_132 ;
	7'h1a :
		TR_145 = TR_132 ;
	7'h1b :
		TR_145 = TR_132 ;
	7'h1c :
		TR_145 = TR_132 ;
	7'h1d :
		TR_145 = TR_132 ;
	7'h1e :
		TR_145 = TR_132 ;
	7'h1f :
		TR_145 = TR_132 ;
	7'h20 :
		TR_145 = TR_132 ;
	7'h21 :
		TR_145 = TR_132 ;
	7'h22 :
		TR_145 = TR_132 ;
	7'h23 :
		TR_145 = TR_132 ;
	7'h24 :
		TR_145 = TR_132 ;
	7'h25 :
		TR_145 = TR_132 ;
	7'h26 :
		TR_145 = TR_132 ;
	7'h27 :
		TR_145 = TR_132 ;
	7'h28 :
		TR_145 = TR_132 ;
	7'h29 :
		TR_145 = TR_132 ;
	7'h2a :
		TR_145 = TR_132 ;
	7'h2b :
		TR_145 = TR_132 ;
	7'h2c :
		TR_145 = TR_132 ;
	7'h2d :
		TR_145 = TR_132 ;
	7'h2e :
		TR_145 = TR_132 ;
	7'h2f :
		TR_145 = TR_132 ;
	7'h30 :
		TR_145 = TR_132 ;
	7'h31 :
		TR_145 = TR_132 ;
	7'h32 :
		TR_145 = TR_132 ;
	7'h33 :
		TR_145 = TR_132 ;
	7'h34 :
		TR_145 = TR_132 ;
	7'h35 :
		TR_145 = TR_132 ;
	7'h36 :
		TR_145 = TR_132 ;
	7'h37 :
		TR_145 = TR_132 ;
	7'h38 :
		TR_145 = TR_132 ;
	7'h39 :
		TR_145 = TR_132 ;
	7'h3a :
		TR_145 = TR_132 ;
	7'h3b :
		TR_145 = TR_132 ;
	7'h3c :
		TR_145 = TR_132 ;
	7'h3d :
		TR_145 = TR_132 ;
	7'h3e :
		TR_145 = TR_132 ;
	7'h3f :
		TR_145 = TR_132 ;
	7'h40 :
		TR_145 = TR_132 ;
	7'h41 :
		TR_145 = TR_132 ;
	7'h42 :
		TR_145 = TR_132 ;
	7'h43 :
		TR_145 = TR_132 ;
	7'h44 :
		TR_145 = TR_132 ;
	7'h45 :
		TR_145 = TR_132 ;
	7'h46 :
		TR_145 = TR_132 ;
	7'h47 :
		TR_145 = TR_132 ;
	7'h48 :
		TR_145 = TR_132 ;
	7'h49 :
		TR_145 = TR_132 ;
	7'h4a :
		TR_145 = TR_132 ;
	7'h4b :
		TR_145 = TR_132 ;
	7'h4c :
		TR_145 = TR_132 ;
	7'h4d :
		TR_145 = TR_132 ;
	7'h4e :
		TR_145 = TR_132 ;
	7'h4f :
		TR_145 = TR_132 ;
	7'h50 :
		TR_145 = TR_132 ;
	7'h51 :
		TR_145 = TR_132 ;
	7'h52 :
		TR_145 = TR_132 ;
	7'h53 :
		TR_145 = TR_132 ;
	7'h54 :
		TR_145 = TR_132 ;
	7'h55 :
		TR_145 = TR_132 ;
	7'h56 :
		TR_145 = TR_132 ;
	7'h57 :
		TR_145 = TR_132 ;
	7'h58 :
		TR_145 = TR_132 ;
	7'h59 :
		TR_145 = TR_132 ;
	7'h5a :
		TR_145 = TR_132 ;
	7'h5b :
		TR_145 = TR_132 ;
	7'h5c :
		TR_145 = TR_132 ;
	7'h5d :
		TR_145 = TR_132 ;
	7'h5e :
		TR_145 = TR_132 ;
	7'h5f :
		TR_145 = TR_132 ;
	7'h60 :
		TR_145 = TR_132 ;
	7'h61 :
		TR_145 = TR_132 ;
	7'h62 :
		TR_145 = TR_132 ;
	7'h63 :
		TR_145 = TR_132 ;
	7'h64 :
		TR_145 = TR_132 ;
	7'h65 :
		TR_145 = TR_132 ;
	7'h66 :
		TR_145 = TR_132 ;
	7'h67 :
		TR_145 = TR_132 ;
	7'h68 :
		TR_145 = TR_132 ;
	7'h69 :
		TR_145 = TR_132 ;
	7'h6a :
		TR_145 = TR_132 ;
	7'h6b :
		TR_145 = TR_132 ;
	7'h6c :
		TR_145 = TR_132 ;
	7'h6d :
		TR_145 = TR_132 ;
	7'h6e :
		TR_145 = TR_132 ;
	7'h6f :
		TR_145 = TR_132 ;
	7'h70 :
		TR_145 = TR_132 ;
	7'h71 :
		TR_145 = TR_132 ;
	7'h72 :
		TR_145 = TR_132 ;
	7'h73 :
		TR_145 = TR_132 ;
	7'h74 :
		TR_145 = TR_132 ;
	7'h75 :
		TR_145 = TR_132 ;
	7'h76 :
		TR_145 = TR_132 ;
	7'h77 :
		TR_145 = TR_132 ;
	7'h78 :
		TR_145 = 9'h000 ;	// line#=../rle.cpp:80
	7'h79 :
		TR_145 = TR_132 ;
	7'h7a :
		TR_145 = TR_132 ;
	7'h7b :
		TR_145 = TR_132 ;
	7'h7c :
		TR_145 = TR_132 ;
	7'h7d :
		TR_145 = TR_132 ;
	7'h7e :
		TR_145 = TR_132 ;
	7'h7f :
		TR_145 = TR_132 ;
	default :
		TR_145 = 9'hx ;
	endcase
always @ ( TR_145 or U_173 or sub8u_71ot or U_183 or RG_rl_189 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_120_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h78 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_120_t = ( ( { 9{ M_180 } } & RG_rl_189 )
		| ( { 9{ U_173 } } & TR_145 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_120_en = ( M_180 | RG_rl_120_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_120_en )
		RG_rl_120 <= RG_rl_120_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_133 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_144 = TR_133 ;
	7'h01 :
		TR_144 = TR_133 ;
	7'h02 :
		TR_144 = TR_133 ;
	7'h03 :
		TR_144 = TR_133 ;
	7'h04 :
		TR_144 = TR_133 ;
	7'h05 :
		TR_144 = TR_133 ;
	7'h06 :
		TR_144 = TR_133 ;
	7'h07 :
		TR_144 = TR_133 ;
	7'h08 :
		TR_144 = TR_133 ;
	7'h09 :
		TR_144 = TR_133 ;
	7'h0a :
		TR_144 = TR_133 ;
	7'h0b :
		TR_144 = TR_133 ;
	7'h0c :
		TR_144 = TR_133 ;
	7'h0d :
		TR_144 = TR_133 ;
	7'h0e :
		TR_144 = TR_133 ;
	7'h0f :
		TR_144 = TR_133 ;
	7'h10 :
		TR_144 = TR_133 ;
	7'h11 :
		TR_144 = TR_133 ;
	7'h12 :
		TR_144 = TR_133 ;
	7'h13 :
		TR_144 = TR_133 ;
	7'h14 :
		TR_144 = TR_133 ;
	7'h15 :
		TR_144 = TR_133 ;
	7'h16 :
		TR_144 = TR_133 ;
	7'h17 :
		TR_144 = TR_133 ;
	7'h18 :
		TR_144 = TR_133 ;
	7'h19 :
		TR_144 = TR_133 ;
	7'h1a :
		TR_144 = TR_133 ;
	7'h1b :
		TR_144 = TR_133 ;
	7'h1c :
		TR_144 = TR_133 ;
	7'h1d :
		TR_144 = TR_133 ;
	7'h1e :
		TR_144 = TR_133 ;
	7'h1f :
		TR_144 = TR_133 ;
	7'h20 :
		TR_144 = TR_133 ;
	7'h21 :
		TR_144 = TR_133 ;
	7'h22 :
		TR_144 = TR_133 ;
	7'h23 :
		TR_144 = TR_133 ;
	7'h24 :
		TR_144 = TR_133 ;
	7'h25 :
		TR_144 = TR_133 ;
	7'h26 :
		TR_144 = TR_133 ;
	7'h27 :
		TR_144 = TR_133 ;
	7'h28 :
		TR_144 = TR_133 ;
	7'h29 :
		TR_144 = TR_133 ;
	7'h2a :
		TR_144 = TR_133 ;
	7'h2b :
		TR_144 = TR_133 ;
	7'h2c :
		TR_144 = TR_133 ;
	7'h2d :
		TR_144 = TR_133 ;
	7'h2e :
		TR_144 = TR_133 ;
	7'h2f :
		TR_144 = TR_133 ;
	7'h30 :
		TR_144 = TR_133 ;
	7'h31 :
		TR_144 = TR_133 ;
	7'h32 :
		TR_144 = TR_133 ;
	7'h33 :
		TR_144 = TR_133 ;
	7'h34 :
		TR_144 = TR_133 ;
	7'h35 :
		TR_144 = TR_133 ;
	7'h36 :
		TR_144 = TR_133 ;
	7'h37 :
		TR_144 = TR_133 ;
	7'h38 :
		TR_144 = TR_133 ;
	7'h39 :
		TR_144 = TR_133 ;
	7'h3a :
		TR_144 = TR_133 ;
	7'h3b :
		TR_144 = TR_133 ;
	7'h3c :
		TR_144 = TR_133 ;
	7'h3d :
		TR_144 = TR_133 ;
	7'h3e :
		TR_144 = TR_133 ;
	7'h3f :
		TR_144 = TR_133 ;
	7'h40 :
		TR_144 = TR_133 ;
	7'h41 :
		TR_144 = TR_133 ;
	7'h42 :
		TR_144 = TR_133 ;
	7'h43 :
		TR_144 = TR_133 ;
	7'h44 :
		TR_144 = TR_133 ;
	7'h45 :
		TR_144 = TR_133 ;
	7'h46 :
		TR_144 = TR_133 ;
	7'h47 :
		TR_144 = TR_133 ;
	7'h48 :
		TR_144 = TR_133 ;
	7'h49 :
		TR_144 = TR_133 ;
	7'h4a :
		TR_144 = TR_133 ;
	7'h4b :
		TR_144 = TR_133 ;
	7'h4c :
		TR_144 = TR_133 ;
	7'h4d :
		TR_144 = TR_133 ;
	7'h4e :
		TR_144 = TR_133 ;
	7'h4f :
		TR_144 = TR_133 ;
	7'h50 :
		TR_144 = TR_133 ;
	7'h51 :
		TR_144 = TR_133 ;
	7'h52 :
		TR_144 = TR_133 ;
	7'h53 :
		TR_144 = TR_133 ;
	7'h54 :
		TR_144 = TR_133 ;
	7'h55 :
		TR_144 = TR_133 ;
	7'h56 :
		TR_144 = TR_133 ;
	7'h57 :
		TR_144 = TR_133 ;
	7'h58 :
		TR_144 = TR_133 ;
	7'h59 :
		TR_144 = TR_133 ;
	7'h5a :
		TR_144 = TR_133 ;
	7'h5b :
		TR_144 = TR_133 ;
	7'h5c :
		TR_144 = TR_133 ;
	7'h5d :
		TR_144 = TR_133 ;
	7'h5e :
		TR_144 = TR_133 ;
	7'h5f :
		TR_144 = TR_133 ;
	7'h60 :
		TR_144 = TR_133 ;
	7'h61 :
		TR_144 = TR_133 ;
	7'h62 :
		TR_144 = TR_133 ;
	7'h63 :
		TR_144 = TR_133 ;
	7'h64 :
		TR_144 = TR_133 ;
	7'h65 :
		TR_144 = TR_133 ;
	7'h66 :
		TR_144 = TR_133 ;
	7'h67 :
		TR_144 = TR_133 ;
	7'h68 :
		TR_144 = TR_133 ;
	7'h69 :
		TR_144 = TR_133 ;
	7'h6a :
		TR_144 = TR_133 ;
	7'h6b :
		TR_144 = TR_133 ;
	7'h6c :
		TR_144 = TR_133 ;
	7'h6d :
		TR_144 = TR_133 ;
	7'h6e :
		TR_144 = TR_133 ;
	7'h6f :
		TR_144 = TR_133 ;
	7'h70 :
		TR_144 = TR_133 ;
	7'h71 :
		TR_144 = TR_133 ;
	7'h72 :
		TR_144 = TR_133 ;
	7'h73 :
		TR_144 = TR_133 ;
	7'h74 :
		TR_144 = TR_133 ;
	7'h75 :
		TR_144 = TR_133 ;
	7'h76 :
		TR_144 = TR_133 ;
	7'h77 :
		TR_144 = TR_133 ;
	7'h78 :
		TR_144 = TR_133 ;
	7'h79 :
		TR_144 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7a :
		TR_144 = TR_133 ;
	7'h7b :
		TR_144 = TR_133 ;
	7'h7c :
		TR_144 = TR_133 ;
	7'h7d :
		TR_144 = TR_133 ;
	7'h7e :
		TR_144 = TR_133 ;
	7'h7f :
		TR_144 = TR_133 ;
	default :
		TR_144 = 9'hx ;
	endcase
always @ ( TR_144 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_58 or 
	U_174 or RG_rl_189 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_121_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h79 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_121_t = ( ( { 9{ ST1_03d } } & RG_rl_189 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_58 )
		| ( { 9{ U_173 } } & TR_144 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_121_en = ( ST1_03d | U_174 | RG_rl_121_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_121_en )
		RG_rl_121 <= RG_rl_121_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_134 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_143 = TR_134 ;
	7'h01 :
		TR_143 = TR_134 ;
	7'h02 :
		TR_143 = TR_134 ;
	7'h03 :
		TR_143 = TR_134 ;
	7'h04 :
		TR_143 = TR_134 ;
	7'h05 :
		TR_143 = TR_134 ;
	7'h06 :
		TR_143 = TR_134 ;
	7'h07 :
		TR_143 = TR_134 ;
	7'h08 :
		TR_143 = TR_134 ;
	7'h09 :
		TR_143 = TR_134 ;
	7'h0a :
		TR_143 = TR_134 ;
	7'h0b :
		TR_143 = TR_134 ;
	7'h0c :
		TR_143 = TR_134 ;
	7'h0d :
		TR_143 = TR_134 ;
	7'h0e :
		TR_143 = TR_134 ;
	7'h0f :
		TR_143 = TR_134 ;
	7'h10 :
		TR_143 = TR_134 ;
	7'h11 :
		TR_143 = TR_134 ;
	7'h12 :
		TR_143 = TR_134 ;
	7'h13 :
		TR_143 = TR_134 ;
	7'h14 :
		TR_143 = TR_134 ;
	7'h15 :
		TR_143 = TR_134 ;
	7'h16 :
		TR_143 = TR_134 ;
	7'h17 :
		TR_143 = TR_134 ;
	7'h18 :
		TR_143 = TR_134 ;
	7'h19 :
		TR_143 = TR_134 ;
	7'h1a :
		TR_143 = TR_134 ;
	7'h1b :
		TR_143 = TR_134 ;
	7'h1c :
		TR_143 = TR_134 ;
	7'h1d :
		TR_143 = TR_134 ;
	7'h1e :
		TR_143 = TR_134 ;
	7'h1f :
		TR_143 = TR_134 ;
	7'h20 :
		TR_143 = TR_134 ;
	7'h21 :
		TR_143 = TR_134 ;
	7'h22 :
		TR_143 = TR_134 ;
	7'h23 :
		TR_143 = TR_134 ;
	7'h24 :
		TR_143 = TR_134 ;
	7'h25 :
		TR_143 = TR_134 ;
	7'h26 :
		TR_143 = TR_134 ;
	7'h27 :
		TR_143 = TR_134 ;
	7'h28 :
		TR_143 = TR_134 ;
	7'h29 :
		TR_143 = TR_134 ;
	7'h2a :
		TR_143 = TR_134 ;
	7'h2b :
		TR_143 = TR_134 ;
	7'h2c :
		TR_143 = TR_134 ;
	7'h2d :
		TR_143 = TR_134 ;
	7'h2e :
		TR_143 = TR_134 ;
	7'h2f :
		TR_143 = TR_134 ;
	7'h30 :
		TR_143 = TR_134 ;
	7'h31 :
		TR_143 = TR_134 ;
	7'h32 :
		TR_143 = TR_134 ;
	7'h33 :
		TR_143 = TR_134 ;
	7'h34 :
		TR_143 = TR_134 ;
	7'h35 :
		TR_143 = TR_134 ;
	7'h36 :
		TR_143 = TR_134 ;
	7'h37 :
		TR_143 = TR_134 ;
	7'h38 :
		TR_143 = TR_134 ;
	7'h39 :
		TR_143 = TR_134 ;
	7'h3a :
		TR_143 = TR_134 ;
	7'h3b :
		TR_143 = TR_134 ;
	7'h3c :
		TR_143 = TR_134 ;
	7'h3d :
		TR_143 = TR_134 ;
	7'h3e :
		TR_143 = TR_134 ;
	7'h3f :
		TR_143 = TR_134 ;
	7'h40 :
		TR_143 = TR_134 ;
	7'h41 :
		TR_143 = TR_134 ;
	7'h42 :
		TR_143 = TR_134 ;
	7'h43 :
		TR_143 = TR_134 ;
	7'h44 :
		TR_143 = TR_134 ;
	7'h45 :
		TR_143 = TR_134 ;
	7'h46 :
		TR_143 = TR_134 ;
	7'h47 :
		TR_143 = TR_134 ;
	7'h48 :
		TR_143 = TR_134 ;
	7'h49 :
		TR_143 = TR_134 ;
	7'h4a :
		TR_143 = TR_134 ;
	7'h4b :
		TR_143 = TR_134 ;
	7'h4c :
		TR_143 = TR_134 ;
	7'h4d :
		TR_143 = TR_134 ;
	7'h4e :
		TR_143 = TR_134 ;
	7'h4f :
		TR_143 = TR_134 ;
	7'h50 :
		TR_143 = TR_134 ;
	7'h51 :
		TR_143 = TR_134 ;
	7'h52 :
		TR_143 = TR_134 ;
	7'h53 :
		TR_143 = TR_134 ;
	7'h54 :
		TR_143 = TR_134 ;
	7'h55 :
		TR_143 = TR_134 ;
	7'h56 :
		TR_143 = TR_134 ;
	7'h57 :
		TR_143 = TR_134 ;
	7'h58 :
		TR_143 = TR_134 ;
	7'h59 :
		TR_143 = TR_134 ;
	7'h5a :
		TR_143 = TR_134 ;
	7'h5b :
		TR_143 = TR_134 ;
	7'h5c :
		TR_143 = TR_134 ;
	7'h5d :
		TR_143 = TR_134 ;
	7'h5e :
		TR_143 = TR_134 ;
	7'h5f :
		TR_143 = TR_134 ;
	7'h60 :
		TR_143 = TR_134 ;
	7'h61 :
		TR_143 = TR_134 ;
	7'h62 :
		TR_143 = TR_134 ;
	7'h63 :
		TR_143 = TR_134 ;
	7'h64 :
		TR_143 = TR_134 ;
	7'h65 :
		TR_143 = TR_134 ;
	7'h66 :
		TR_143 = TR_134 ;
	7'h67 :
		TR_143 = TR_134 ;
	7'h68 :
		TR_143 = TR_134 ;
	7'h69 :
		TR_143 = TR_134 ;
	7'h6a :
		TR_143 = TR_134 ;
	7'h6b :
		TR_143 = TR_134 ;
	7'h6c :
		TR_143 = TR_134 ;
	7'h6d :
		TR_143 = TR_134 ;
	7'h6e :
		TR_143 = TR_134 ;
	7'h6f :
		TR_143 = TR_134 ;
	7'h70 :
		TR_143 = TR_134 ;
	7'h71 :
		TR_143 = TR_134 ;
	7'h72 :
		TR_143 = TR_134 ;
	7'h73 :
		TR_143 = TR_134 ;
	7'h74 :
		TR_143 = TR_134 ;
	7'h75 :
		TR_143 = TR_134 ;
	7'h76 :
		TR_143 = TR_134 ;
	7'h77 :
		TR_143 = TR_134 ;
	7'h78 :
		TR_143 = TR_134 ;
	7'h79 :
		TR_143 = TR_134 ;
	7'h7a :
		TR_143 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7b :
		TR_143 = TR_134 ;
	7'h7c :
		TR_143 = TR_134 ;
	7'h7d :
		TR_143 = TR_134 ;
	7'h7e :
		TR_143 = TR_134 ;
	7'h7f :
		TR_143 = TR_134 ;
	default :
		TR_143 = 9'hx ;
	endcase
always @ ( TR_143 or U_173 or sub8u_71ot or U_183 or RG_rl_190 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_122_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h7a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_122_t = ( ( { 9{ M_180 } } & RG_rl_190 )
		| ( { 9{ U_173 } } & TR_143 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_122_en = ( M_180 | RG_rl_122_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_122_en )
		RG_rl_122 <= RG_rl_122_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_135 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_142 = TR_135 ;
	7'h01 :
		TR_142 = TR_135 ;
	7'h02 :
		TR_142 = TR_135 ;
	7'h03 :
		TR_142 = TR_135 ;
	7'h04 :
		TR_142 = TR_135 ;
	7'h05 :
		TR_142 = TR_135 ;
	7'h06 :
		TR_142 = TR_135 ;
	7'h07 :
		TR_142 = TR_135 ;
	7'h08 :
		TR_142 = TR_135 ;
	7'h09 :
		TR_142 = TR_135 ;
	7'h0a :
		TR_142 = TR_135 ;
	7'h0b :
		TR_142 = TR_135 ;
	7'h0c :
		TR_142 = TR_135 ;
	7'h0d :
		TR_142 = TR_135 ;
	7'h0e :
		TR_142 = TR_135 ;
	7'h0f :
		TR_142 = TR_135 ;
	7'h10 :
		TR_142 = TR_135 ;
	7'h11 :
		TR_142 = TR_135 ;
	7'h12 :
		TR_142 = TR_135 ;
	7'h13 :
		TR_142 = TR_135 ;
	7'h14 :
		TR_142 = TR_135 ;
	7'h15 :
		TR_142 = TR_135 ;
	7'h16 :
		TR_142 = TR_135 ;
	7'h17 :
		TR_142 = TR_135 ;
	7'h18 :
		TR_142 = TR_135 ;
	7'h19 :
		TR_142 = TR_135 ;
	7'h1a :
		TR_142 = TR_135 ;
	7'h1b :
		TR_142 = TR_135 ;
	7'h1c :
		TR_142 = TR_135 ;
	7'h1d :
		TR_142 = TR_135 ;
	7'h1e :
		TR_142 = TR_135 ;
	7'h1f :
		TR_142 = TR_135 ;
	7'h20 :
		TR_142 = TR_135 ;
	7'h21 :
		TR_142 = TR_135 ;
	7'h22 :
		TR_142 = TR_135 ;
	7'h23 :
		TR_142 = TR_135 ;
	7'h24 :
		TR_142 = TR_135 ;
	7'h25 :
		TR_142 = TR_135 ;
	7'h26 :
		TR_142 = TR_135 ;
	7'h27 :
		TR_142 = TR_135 ;
	7'h28 :
		TR_142 = TR_135 ;
	7'h29 :
		TR_142 = TR_135 ;
	7'h2a :
		TR_142 = TR_135 ;
	7'h2b :
		TR_142 = TR_135 ;
	7'h2c :
		TR_142 = TR_135 ;
	7'h2d :
		TR_142 = TR_135 ;
	7'h2e :
		TR_142 = TR_135 ;
	7'h2f :
		TR_142 = TR_135 ;
	7'h30 :
		TR_142 = TR_135 ;
	7'h31 :
		TR_142 = TR_135 ;
	7'h32 :
		TR_142 = TR_135 ;
	7'h33 :
		TR_142 = TR_135 ;
	7'h34 :
		TR_142 = TR_135 ;
	7'h35 :
		TR_142 = TR_135 ;
	7'h36 :
		TR_142 = TR_135 ;
	7'h37 :
		TR_142 = TR_135 ;
	7'h38 :
		TR_142 = TR_135 ;
	7'h39 :
		TR_142 = TR_135 ;
	7'h3a :
		TR_142 = TR_135 ;
	7'h3b :
		TR_142 = TR_135 ;
	7'h3c :
		TR_142 = TR_135 ;
	7'h3d :
		TR_142 = TR_135 ;
	7'h3e :
		TR_142 = TR_135 ;
	7'h3f :
		TR_142 = TR_135 ;
	7'h40 :
		TR_142 = TR_135 ;
	7'h41 :
		TR_142 = TR_135 ;
	7'h42 :
		TR_142 = TR_135 ;
	7'h43 :
		TR_142 = TR_135 ;
	7'h44 :
		TR_142 = TR_135 ;
	7'h45 :
		TR_142 = TR_135 ;
	7'h46 :
		TR_142 = TR_135 ;
	7'h47 :
		TR_142 = TR_135 ;
	7'h48 :
		TR_142 = TR_135 ;
	7'h49 :
		TR_142 = TR_135 ;
	7'h4a :
		TR_142 = TR_135 ;
	7'h4b :
		TR_142 = TR_135 ;
	7'h4c :
		TR_142 = TR_135 ;
	7'h4d :
		TR_142 = TR_135 ;
	7'h4e :
		TR_142 = TR_135 ;
	7'h4f :
		TR_142 = TR_135 ;
	7'h50 :
		TR_142 = TR_135 ;
	7'h51 :
		TR_142 = TR_135 ;
	7'h52 :
		TR_142 = TR_135 ;
	7'h53 :
		TR_142 = TR_135 ;
	7'h54 :
		TR_142 = TR_135 ;
	7'h55 :
		TR_142 = TR_135 ;
	7'h56 :
		TR_142 = TR_135 ;
	7'h57 :
		TR_142 = TR_135 ;
	7'h58 :
		TR_142 = TR_135 ;
	7'h59 :
		TR_142 = TR_135 ;
	7'h5a :
		TR_142 = TR_135 ;
	7'h5b :
		TR_142 = TR_135 ;
	7'h5c :
		TR_142 = TR_135 ;
	7'h5d :
		TR_142 = TR_135 ;
	7'h5e :
		TR_142 = TR_135 ;
	7'h5f :
		TR_142 = TR_135 ;
	7'h60 :
		TR_142 = TR_135 ;
	7'h61 :
		TR_142 = TR_135 ;
	7'h62 :
		TR_142 = TR_135 ;
	7'h63 :
		TR_142 = TR_135 ;
	7'h64 :
		TR_142 = TR_135 ;
	7'h65 :
		TR_142 = TR_135 ;
	7'h66 :
		TR_142 = TR_135 ;
	7'h67 :
		TR_142 = TR_135 ;
	7'h68 :
		TR_142 = TR_135 ;
	7'h69 :
		TR_142 = TR_135 ;
	7'h6a :
		TR_142 = TR_135 ;
	7'h6b :
		TR_142 = TR_135 ;
	7'h6c :
		TR_142 = TR_135 ;
	7'h6d :
		TR_142 = TR_135 ;
	7'h6e :
		TR_142 = TR_135 ;
	7'h6f :
		TR_142 = TR_135 ;
	7'h70 :
		TR_142 = TR_135 ;
	7'h71 :
		TR_142 = TR_135 ;
	7'h72 :
		TR_142 = TR_135 ;
	7'h73 :
		TR_142 = TR_135 ;
	7'h74 :
		TR_142 = TR_135 ;
	7'h75 :
		TR_142 = TR_135 ;
	7'h76 :
		TR_142 = TR_135 ;
	7'h77 :
		TR_142 = TR_135 ;
	7'h78 :
		TR_142 = TR_135 ;
	7'h79 :
		TR_142 = TR_135 ;
	7'h7a :
		TR_142 = TR_135 ;
	7'h7b :
		TR_142 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7c :
		TR_142 = TR_135 ;
	7'h7d :
		TR_142 = TR_135 ;
	7'h7e :
		TR_142 = TR_135 ;
	7'h7f :
		TR_142 = TR_135 ;
	default :
		TR_142 = 9'hx ;
	endcase
always @ ( TR_142 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_59 or 
	U_174 or RG_rl_190 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_123_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h7b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_123_t = ( ( { 9{ ST1_03d } } & RG_rl_190 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_59 )
		| ( { 9{ U_173 } } & TR_142 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_123_en = ( ST1_03d | U_174 | RG_rl_123_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_123_en )
		RG_rl_123 <= RG_rl_123_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_136 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_141 = TR_136 ;
	7'h01 :
		TR_141 = TR_136 ;
	7'h02 :
		TR_141 = TR_136 ;
	7'h03 :
		TR_141 = TR_136 ;
	7'h04 :
		TR_141 = TR_136 ;
	7'h05 :
		TR_141 = TR_136 ;
	7'h06 :
		TR_141 = TR_136 ;
	7'h07 :
		TR_141 = TR_136 ;
	7'h08 :
		TR_141 = TR_136 ;
	7'h09 :
		TR_141 = TR_136 ;
	7'h0a :
		TR_141 = TR_136 ;
	7'h0b :
		TR_141 = TR_136 ;
	7'h0c :
		TR_141 = TR_136 ;
	7'h0d :
		TR_141 = TR_136 ;
	7'h0e :
		TR_141 = TR_136 ;
	7'h0f :
		TR_141 = TR_136 ;
	7'h10 :
		TR_141 = TR_136 ;
	7'h11 :
		TR_141 = TR_136 ;
	7'h12 :
		TR_141 = TR_136 ;
	7'h13 :
		TR_141 = TR_136 ;
	7'h14 :
		TR_141 = TR_136 ;
	7'h15 :
		TR_141 = TR_136 ;
	7'h16 :
		TR_141 = TR_136 ;
	7'h17 :
		TR_141 = TR_136 ;
	7'h18 :
		TR_141 = TR_136 ;
	7'h19 :
		TR_141 = TR_136 ;
	7'h1a :
		TR_141 = TR_136 ;
	7'h1b :
		TR_141 = TR_136 ;
	7'h1c :
		TR_141 = TR_136 ;
	7'h1d :
		TR_141 = TR_136 ;
	7'h1e :
		TR_141 = TR_136 ;
	7'h1f :
		TR_141 = TR_136 ;
	7'h20 :
		TR_141 = TR_136 ;
	7'h21 :
		TR_141 = TR_136 ;
	7'h22 :
		TR_141 = TR_136 ;
	7'h23 :
		TR_141 = TR_136 ;
	7'h24 :
		TR_141 = TR_136 ;
	7'h25 :
		TR_141 = TR_136 ;
	7'h26 :
		TR_141 = TR_136 ;
	7'h27 :
		TR_141 = TR_136 ;
	7'h28 :
		TR_141 = TR_136 ;
	7'h29 :
		TR_141 = TR_136 ;
	7'h2a :
		TR_141 = TR_136 ;
	7'h2b :
		TR_141 = TR_136 ;
	7'h2c :
		TR_141 = TR_136 ;
	7'h2d :
		TR_141 = TR_136 ;
	7'h2e :
		TR_141 = TR_136 ;
	7'h2f :
		TR_141 = TR_136 ;
	7'h30 :
		TR_141 = TR_136 ;
	7'h31 :
		TR_141 = TR_136 ;
	7'h32 :
		TR_141 = TR_136 ;
	7'h33 :
		TR_141 = TR_136 ;
	7'h34 :
		TR_141 = TR_136 ;
	7'h35 :
		TR_141 = TR_136 ;
	7'h36 :
		TR_141 = TR_136 ;
	7'h37 :
		TR_141 = TR_136 ;
	7'h38 :
		TR_141 = TR_136 ;
	7'h39 :
		TR_141 = TR_136 ;
	7'h3a :
		TR_141 = TR_136 ;
	7'h3b :
		TR_141 = TR_136 ;
	7'h3c :
		TR_141 = TR_136 ;
	7'h3d :
		TR_141 = TR_136 ;
	7'h3e :
		TR_141 = TR_136 ;
	7'h3f :
		TR_141 = TR_136 ;
	7'h40 :
		TR_141 = TR_136 ;
	7'h41 :
		TR_141 = TR_136 ;
	7'h42 :
		TR_141 = TR_136 ;
	7'h43 :
		TR_141 = TR_136 ;
	7'h44 :
		TR_141 = TR_136 ;
	7'h45 :
		TR_141 = TR_136 ;
	7'h46 :
		TR_141 = TR_136 ;
	7'h47 :
		TR_141 = TR_136 ;
	7'h48 :
		TR_141 = TR_136 ;
	7'h49 :
		TR_141 = TR_136 ;
	7'h4a :
		TR_141 = TR_136 ;
	7'h4b :
		TR_141 = TR_136 ;
	7'h4c :
		TR_141 = TR_136 ;
	7'h4d :
		TR_141 = TR_136 ;
	7'h4e :
		TR_141 = TR_136 ;
	7'h4f :
		TR_141 = TR_136 ;
	7'h50 :
		TR_141 = TR_136 ;
	7'h51 :
		TR_141 = TR_136 ;
	7'h52 :
		TR_141 = TR_136 ;
	7'h53 :
		TR_141 = TR_136 ;
	7'h54 :
		TR_141 = TR_136 ;
	7'h55 :
		TR_141 = TR_136 ;
	7'h56 :
		TR_141 = TR_136 ;
	7'h57 :
		TR_141 = TR_136 ;
	7'h58 :
		TR_141 = TR_136 ;
	7'h59 :
		TR_141 = TR_136 ;
	7'h5a :
		TR_141 = TR_136 ;
	7'h5b :
		TR_141 = TR_136 ;
	7'h5c :
		TR_141 = TR_136 ;
	7'h5d :
		TR_141 = TR_136 ;
	7'h5e :
		TR_141 = TR_136 ;
	7'h5f :
		TR_141 = TR_136 ;
	7'h60 :
		TR_141 = TR_136 ;
	7'h61 :
		TR_141 = TR_136 ;
	7'h62 :
		TR_141 = TR_136 ;
	7'h63 :
		TR_141 = TR_136 ;
	7'h64 :
		TR_141 = TR_136 ;
	7'h65 :
		TR_141 = TR_136 ;
	7'h66 :
		TR_141 = TR_136 ;
	7'h67 :
		TR_141 = TR_136 ;
	7'h68 :
		TR_141 = TR_136 ;
	7'h69 :
		TR_141 = TR_136 ;
	7'h6a :
		TR_141 = TR_136 ;
	7'h6b :
		TR_141 = TR_136 ;
	7'h6c :
		TR_141 = TR_136 ;
	7'h6d :
		TR_141 = TR_136 ;
	7'h6e :
		TR_141 = TR_136 ;
	7'h6f :
		TR_141 = TR_136 ;
	7'h70 :
		TR_141 = TR_136 ;
	7'h71 :
		TR_141 = TR_136 ;
	7'h72 :
		TR_141 = TR_136 ;
	7'h73 :
		TR_141 = TR_136 ;
	7'h74 :
		TR_141 = TR_136 ;
	7'h75 :
		TR_141 = TR_136 ;
	7'h76 :
		TR_141 = TR_136 ;
	7'h77 :
		TR_141 = TR_136 ;
	7'h78 :
		TR_141 = TR_136 ;
	7'h79 :
		TR_141 = TR_136 ;
	7'h7a :
		TR_141 = TR_136 ;
	7'h7b :
		TR_141 = TR_136 ;
	7'h7c :
		TR_141 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7d :
		TR_141 = TR_136 ;
	7'h7e :
		TR_141 = TR_136 ;
	7'h7f :
		TR_141 = TR_136 ;
	default :
		TR_141 = 9'hx ;
	endcase
always @ ( TR_141 or U_173 or sub8u_71ot or U_183 or RG_rl_191 or M_180 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_124_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h7c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_124_t = ( ( { 9{ M_180 } } & RG_rl_191 )
		| ( { 9{ U_173 } } & TR_141 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_124_en = ( M_180 | RG_rl_124_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_124_en )
		RG_rl_124 <= RG_rl_124_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_137 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_140 = TR_137 ;
	7'h01 :
		TR_140 = TR_137 ;
	7'h02 :
		TR_140 = TR_137 ;
	7'h03 :
		TR_140 = TR_137 ;
	7'h04 :
		TR_140 = TR_137 ;
	7'h05 :
		TR_140 = TR_137 ;
	7'h06 :
		TR_140 = TR_137 ;
	7'h07 :
		TR_140 = TR_137 ;
	7'h08 :
		TR_140 = TR_137 ;
	7'h09 :
		TR_140 = TR_137 ;
	7'h0a :
		TR_140 = TR_137 ;
	7'h0b :
		TR_140 = TR_137 ;
	7'h0c :
		TR_140 = TR_137 ;
	7'h0d :
		TR_140 = TR_137 ;
	7'h0e :
		TR_140 = TR_137 ;
	7'h0f :
		TR_140 = TR_137 ;
	7'h10 :
		TR_140 = TR_137 ;
	7'h11 :
		TR_140 = TR_137 ;
	7'h12 :
		TR_140 = TR_137 ;
	7'h13 :
		TR_140 = TR_137 ;
	7'h14 :
		TR_140 = TR_137 ;
	7'h15 :
		TR_140 = TR_137 ;
	7'h16 :
		TR_140 = TR_137 ;
	7'h17 :
		TR_140 = TR_137 ;
	7'h18 :
		TR_140 = TR_137 ;
	7'h19 :
		TR_140 = TR_137 ;
	7'h1a :
		TR_140 = TR_137 ;
	7'h1b :
		TR_140 = TR_137 ;
	7'h1c :
		TR_140 = TR_137 ;
	7'h1d :
		TR_140 = TR_137 ;
	7'h1e :
		TR_140 = TR_137 ;
	7'h1f :
		TR_140 = TR_137 ;
	7'h20 :
		TR_140 = TR_137 ;
	7'h21 :
		TR_140 = TR_137 ;
	7'h22 :
		TR_140 = TR_137 ;
	7'h23 :
		TR_140 = TR_137 ;
	7'h24 :
		TR_140 = TR_137 ;
	7'h25 :
		TR_140 = TR_137 ;
	7'h26 :
		TR_140 = TR_137 ;
	7'h27 :
		TR_140 = TR_137 ;
	7'h28 :
		TR_140 = TR_137 ;
	7'h29 :
		TR_140 = TR_137 ;
	7'h2a :
		TR_140 = TR_137 ;
	7'h2b :
		TR_140 = TR_137 ;
	7'h2c :
		TR_140 = TR_137 ;
	7'h2d :
		TR_140 = TR_137 ;
	7'h2e :
		TR_140 = TR_137 ;
	7'h2f :
		TR_140 = TR_137 ;
	7'h30 :
		TR_140 = TR_137 ;
	7'h31 :
		TR_140 = TR_137 ;
	7'h32 :
		TR_140 = TR_137 ;
	7'h33 :
		TR_140 = TR_137 ;
	7'h34 :
		TR_140 = TR_137 ;
	7'h35 :
		TR_140 = TR_137 ;
	7'h36 :
		TR_140 = TR_137 ;
	7'h37 :
		TR_140 = TR_137 ;
	7'h38 :
		TR_140 = TR_137 ;
	7'h39 :
		TR_140 = TR_137 ;
	7'h3a :
		TR_140 = TR_137 ;
	7'h3b :
		TR_140 = TR_137 ;
	7'h3c :
		TR_140 = TR_137 ;
	7'h3d :
		TR_140 = TR_137 ;
	7'h3e :
		TR_140 = TR_137 ;
	7'h3f :
		TR_140 = TR_137 ;
	7'h40 :
		TR_140 = TR_137 ;
	7'h41 :
		TR_140 = TR_137 ;
	7'h42 :
		TR_140 = TR_137 ;
	7'h43 :
		TR_140 = TR_137 ;
	7'h44 :
		TR_140 = TR_137 ;
	7'h45 :
		TR_140 = TR_137 ;
	7'h46 :
		TR_140 = TR_137 ;
	7'h47 :
		TR_140 = TR_137 ;
	7'h48 :
		TR_140 = TR_137 ;
	7'h49 :
		TR_140 = TR_137 ;
	7'h4a :
		TR_140 = TR_137 ;
	7'h4b :
		TR_140 = TR_137 ;
	7'h4c :
		TR_140 = TR_137 ;
	7'h4d :
		TR_140 = TR_137 ;
	7'h4e :
		TR_140 = TR_137 ;
	7'h4f :
		TR_140 = TR_137 ;
	7'h50 :
		TR_140 = TR_137 ;
	7'h51 :
		TR_140 = TR_137 ;
	7'h52 :
		TR_140 = TR_137 ;
	7'h53 :
		TR_140 = TR_137 ;
	7'h54 :
		TR_140 = TR_137 ;
	7'h55 :
		TR_140 = TR_137 ;
	7'h56 :
		TR_140 = TR_137 ;
	7'h57 :
		TR_140 = TR_137 ;
	7'h58 :
		TR_140 = TR_137 ;
	7'h59 :
		TR_140 = TR_137 ;
	7'h5a :
		TR_140 = TR_137 ;
	7'h5b :
		TR_140 = TR_137 ;
	7'h5c :
		TR_140 = TR_137 ;
	7'h5d :
		TR_140 = TR_137 ;
	7'h5e :
		TR_140 = TR_137 ;
	7'h5f :
		TR_140 = TR_137 ;
	7'h60 :
		TR_140 = TR_137 ;
	7'h61 :
		TR_140 = TR_137 ;
	7'h62 :
		TR_140 = TR_137 ;
	7'h63 :
		TR_140 = TR_137 ;
	7'h64 :
		TR_140 = TR_137 ;
	7'h65 :
		TR_140 = TR_137 ;
	7'h66 :
		TR_140 = TR_137 ;
	7'h67 :
		TR_140 = TR_137 ;
	7'h68 :
		TR_140 = TR_137 ;
	7'h69 :
		TR_140 = TR_137 ;
	7'h6a :
		TR_140 = TR_137 ;
	7'h6b :
		TR_140 = TR_137 ;
	7'h6c :
		TR_140 = TR_137 ;
	7'h6d :
		TR_140 = TR_137 ;
	7'h6e :
		TR_140 = TR_137 ;
	7'h6f :
		TR_140 = TR_137 ;
	7'h70 :
		TR_140 = TR_137 ;
	7'h71 :
		TR_140 = TR_137 ;
	7'h72 :
		TR_140 = TR_137 ;
	7'h73 :
		TR_140 = TR_137 ;
	7'h74 :
		TR_140 = TR_137 ;
	7'h75 :
		TR_140 = TR_137 ;
	7'h76 :
		TR_140 = TR_137 ;
	7'h77 :
		TR_140 = TR_137 ;
	7'h78 :
		TR_140 = TR_137 ;
	7'h79 :
		TR_140 = TR_137 ;
	7'h7a :
		TR_140 = TR_137 ;
	7'h7b :
		TR_140 = TR_137 ;
	7'h7c :
		TR_140 = TR_137 ;
	7'h7d :
		TR_140 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7e :
		TR_140 = TR_137 ;
	7'h7f :
		TR_140 = TR_137 ;
	default :
		TR_140 = 9'hx ;
	endcase
always @ ( TR_140 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_60 or 
	U_174 or RG_rl_191 or ST1_03d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_125_t_c1 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h7d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_125_t = ( ( { 9{ ST1_03d } } & RG_rl_191 )
		| ( { 9{ U_174 } } & RG_quantized_block_rl_60 )
		| ( { 9{ U_173 } } & TR_140 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_125_en = ( ST1_03d | U_174 | RG_rl_125_t_c1 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_125_en )
		RG_rl_125 <= RG_rl_125_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_138 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		TR_139 = TR_138 ;
	7'h01 :
		TR_139 = TR_138 ;
	7'h02 :
		TR_139 = TR_138 ;
	7'h03 :
		TR_139 = TR_138 ;
	7'h04 :
		TR_139 = TR_138 ;
	7'h05 :
		TR_139 = TR_138 ;
	7'h06 :
		TR_139 = TR_138 ;
	7'h07 :
		TR_139 = TR_138 ;
	7'h08 :
		TR_139 = TR_138 ;
	7'h09 :
		TR_139 = TR_138 ;
	7'h0a :
		TR_139 = TR_138 ;
	7'h0b :
		TR_139 = TR_138 ;
	7'h0c :
		TR_139 = TR_138 ;
	7'h0d :
		TR_139 = TR_138 ;
	7'h0e :
		TR_139 = TR_138 ;
	7'h0f :
		TR_139 = TR_138 ;
	7'h10 :
		TR_139 = TR_138 ;
	7'h11 :
		TR_139 = TR_138 ;
	7'h12 :
		TR_139 = TR_138 ;
	7'h13 :
		TR_139 = TR_138 ;
	7'h14 :
		TR_139 = TR_138 ;
	7'h15 :
		TR_139 = TR_138 ;
	7'h16 :
		TR_139 = TR_138 ;
	7'h17 :
		TR_139 = TR_138 ;
	7'h18 :
		TR_139 = TR_138 ;
	7'h19 :
		TR_139 = TR_138 ;
	7'h1a :
		TR_139 = TR_138 ;
	7'h1b :
		TR_139 = TR_138 ;
	7'h1c :
		TR_139 = TR_138 ;
	7'h1d :
		TR_139 = TR_138 ;
	7'h1e :
		TR_139 = TR_138 ;
	7'h1f :
		TR_139 = TR_138 ;
	7'h20 :
		TR_139 = TR_138 ;
	7'h21 :
		TR_139 = TR_138 ;
	7'h22 :
		TR_139 = TR_138 ;
	7'h23 :
		TR_139 = TR_138 ;
	7'h24 :
		TR_139 = TR_138 ;
	7'h25 :
		TR_139 = TR_138 ;
	7'h26 :
		TR_139 = TR_138 ;
	7'h27 :
		TR_139 = TR_138 ;
	7'h28 :
		TR_139 = TR_138 ;
	7'h29 :
		TR_139 = TR_138 ;
	7'h2a :
		TR_139 = TR_138 ;
	7'h2b :
		TR_139 = TR_138 ;
	7'h2c :
		TR_139 = TR_138 ;
	7'h2d :
		TR_139 = TR_138 ;
	7'h2e :
		TR_139 = TR_138 ;
	7'h2f :
		TR_139 = TR_138 ;
	7'h30 :
		TR_139 = TR_138 ;
	7'h31 :
		TR_139 = TR_138 ;
	7'h32 :
		TR_139 = TR_138 ;
	7'h33 :
		TR_139 = TR_138 ;
	7'h34 :
		TR_139 = TR_138 ;
	7'h35 :
		TR_139 = TR_138 ;
	7'h36 :
		TR_139 = TR_138 ;
	7'h37 :
		TR_139 = TR_138 ;
	7'h38 :
		TR_139 = TR_138 ;
	7'h39 :
		TR_139 = TR_138 ;
	7'h3a :
		TR_139 = TR_138 ;
	7'h3b :
		TR_139 = TR_138 ;
	7'h3c :
		TR_139 = TR_138 ;
	7'h3d :
		TR_139 = TR_138 ;
	7'h3e :
		TR_139 = TR_138 ;
	7'h3f :
		TR_139 = TR_138 ;
	7'h40 :
		TR_139 = TR_138 ;
	7'h41 :
		TR_139 = TR_138 ;
	7'h42 :
		TR_139 = TR_138 ;
	7'h43 :
		TR_139 = TR_138 ;
	7'h44 :
		TR_139 = TR_138 ;
	7'h45 :
		TR_139 = TR_138 ;
	7'h46 :
		TR_139 = TR_138 ;
	7'h47 :
		TR_139 = TR_138 ;
	7'h48 :
		TR_139 = TR_138 ;
	7'h49 :
		TR_139 = TR_138 ;
	7'h4a :
		TR_139 = TR_138 ;
	7'h4b :
		TR_139 = TR_138 ;
	7'h4c :
		TR_139 = TR_138 ;
	7'h4d :
		TR_139 = TR_138 ;
	7'h4e :
		TR_139 = TR_138 ;
	7'h4f :
		TR_139 = TR_138 ;
	7'h50 :
		TR_139 = TR_138 ;
	7'h51 :
		TR_139 = TR_138 ;
	7'h52 :
		TR_139 = TR_138 ;
	7'h53 :
		TR_139 = TR_138 ;
	7'h54 :
		TR_139 = TR_138 ;
	7'h55 :
		TR_139 = TR_138 ;
	7'h56 :
		TR_139 = TR_138 ;
	7'h57 :
		TR_139 = TR_138 ;
	7'h58 :
		TR_139 = TR_138 ;
	7'h59 :
		TR_139 = TR_138 ;
	7'h5a :
		TR_139 = TR_138 ;
	7'h5b :
		TR_139 = TR_138 ;
	7'h5c :
		TR_139 = TR_138 ;
	7'h5d :
		TR_139 = TR_138 ;
	7'h5e :
		TR_139 = TR_138 ;
	7'h5f :
		TR_139 = TR_138 ;
	7'h60 :
		TR_139 = TR_138 ;
	7'h61 :
		TR_139 = TR_138 ;
	7'h62 :
		TR_139 = TR_138 ;
	7'h63 :
		TR_139 = TR_138 ;
	7'h64 :
		TR_139 = TR_138 ;
	7'h65 :
		TR_139 = TR_138 ;
	7'h66 :
		TR_139 = TR_138 ;
	7'h67 :
		TR_139 = TR_138 ;
	7'h68 :
		TR_139 = TR_138 ;
	7'h69 :
		TR_139 = TR_138 ;
	7'h6a :
		TR_139 = TR_138 ;
	7'h6b :
		TR_139 = TR_138 ;
	7'h6c :
		TR_139 = TR_138 ;
	7'h6d :
		TR_139 = TR_138 ;
	7'h6e :
		TR_139 = TR_138 ;
	7'h6f :
		TR_139 = TR_138 ;
	7'h70 :
		TR_139 = TR_138 ;
	7'h71 :
		TR_139 = TR_138 ;
	7'h72 :
		TR_139 = TR_138 ;
	7'h73 :
		TR_139 = TR_138 ;
	7'h74 :
		TR_139 = TR_138 ;
	7'h75 :
		TR_139 = TR_138 ;
	7'h76 :
		TR_139 = TR_138 ;
	7'h77 :
		TR_139 = TR_138 ;
	7'h78 :
		TR_139 = TR_138 ;
	7'h79 :
		TR_139 = TR_138 ;
	7'h7a :
		TR_139 = TR_138 ;
	7'h7b :
		TR_139 = TR_138 ;
	7'h7c :
		TR_139 = TR_138 ;
	7'h7d :
		TR_139 = TR_138 ;
	7'h7e :
		TR_139 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7f :
		TR_139 = TR_138 ;
	default :
		TR_139 = 9'hx ;
	endcase
always @ ( TR_139 or U_173 or sub8u_71ot or U_183 or RG_quantized_block_rl_61 or 
	U_174 or ST1_02d )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_126_t_c1 = ( ST1_02d | U_174 ) ;
	RG_rl_126_t_c2 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h7e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_126_t = ( ( { 9{ RG_rl_126_t_c1 } } & RG_quantized_block_rl_61 )
		| ( { 9{ U_173 } } & TR_139 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_126_en = ( RG_rl_126_t_c1 | RG_rl_126_t_c2 | U_173 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_126_en )
		RG_rl_126 <= RG_rl_126_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( rl_a127_t2 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h01 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h02 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h03 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h04 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h05 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h06 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h07 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h08 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h09 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h0a :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h0b :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h0c :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h0d :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h0e :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h0f :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h10 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h11 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h12 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h13 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h14 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h15 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h16 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h17 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h18 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h19 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h1a :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h1b :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h1c :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h1d :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h1e :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h1f :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h20 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h21 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h22 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h23 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h24 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h25 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h26 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h27 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h28 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h29 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h2a :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h2b :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h2c :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h2d :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h2e :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h2f :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h30 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h31 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h32 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h33 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h34 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h35 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h36 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h37 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h38 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h39 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h3a :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h3b :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h3c :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h3d :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h3e :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h3f :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h40 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h41 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h42 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h43 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h44 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h45 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h46 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h47 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h48 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h49 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h4a :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h4b :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h4c :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h4d :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h4e :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h4f :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h50 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h51 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h52 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h53 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h54 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h55 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h56 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h57 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h58 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h59 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h5a :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h5b :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h5c :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h5d :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h5e :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h5f :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h60 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h61 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h62 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h63 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h64 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h65 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h66 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h67 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h68 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h69 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h6a :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h6b :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h6c :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h6d :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h6e :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h6f :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h70 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h71 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h72 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h73 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h74 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h75 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h76 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h77 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h78 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h79 :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h7a :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h7b :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h7c :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h7d :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h7e :
		RG_rl_127_t1 = rl_a127_t2 ;
	7'h7f :
		RG_rl_127_t1 = 9'h000 ;	// line#=../rle.cpp:80
	default :
		RG_rl_127_t1 = 9'hx ;
	endcase
always @ ( RG_rl_127_t1 or U_173 or sub8u_71ot or U_183 or RG_k_quantized_block_rl_01 or 
	U_174 or C_07 or ST1_05d or ST1_02d )	// line#=../rle.cpp:57,58,83,84,85
	begin
	RG_rl_127_t_c1 = ( ( ST1_02d | ( ST1_05d & C_07 ) ) | U_174 ) ;
	RG_rl_127_t_c2 = ( U_183 & ( ~|( sub8u_71ot ^ 7'h7f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_127_t = ( ( { 9{ RG_rl_127_t_c1 } } & RG_k_quantized_block_rl_01 )
		| ( { 9{ U_173 } } & RG_rl_127_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_127_en = ( RG_rl_127_t_c1 | RG_rl_127_t_c2 | U_173 ) ;	// line#=../rle.cpp:57,58,83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:57,58,83,84,85
	if ( RG_rl_127_en )
		RG_rl_127 <= RG_rl_127_t ;	// line#=../rle.cpp:57,58,79,80,83,84,85
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h01 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h01 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_t = ( ( { 9{ RG_zz_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_en = ( RG_zz_t_c1 | RG_zz_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_en )
		RG_zz <= RG_zz_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_1_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h02 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_1_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h02 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_1_t = ( ( { 9{ RG_zz_1_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_1_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_1_en = ( RG_zz_1_t_c1 | RG_zz_1_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_1_en )
		RG_zz_1 <= RG_zz_1_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_2_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h03 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_2_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h03 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_2_t = ( ( { 9{ RG_zz_2_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_2_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_2_en = ( RG_zz_2_t_c1 | RG_zz_2_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_2_en )
		RG_zz_2 <= RG_zz_2_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_3_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h04 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_3_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h04 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_3_t = ( ( { 9{ RG_zz_3_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_3_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_3_en = ( RG_zz_3_t_c1 | RG_zz_3_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_3_en )
		RG_zz_3 <= RG_zz_3_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_4_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h05 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_4_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h05 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_4_t = ( ( { 9{ RG_zz_4_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_4_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_4_en = ( RG_zz_4_t_c1 | RG_zz_4_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_4_en )
		RG_zz_4 <= RG_zz_4_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_5_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h06 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_5_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h06 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_5_t = ( ( { 9{ RG_zz_5_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_5_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_5_en = ( RG_zz_5_t_c1 | RG_zz_5_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_5_en )
		RG_zz_5 <= RG_zz_5_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_6_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h07 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_6_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h07 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_6_t = ( ( { 9{ RG_zz_6_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_6_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_6_en = ( RG_zz_6_t_c1 | RG_zz_6_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_6_en )
		RG_zz_6 <= RG_zz_6_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_7_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h08 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_7_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h08 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_7_t = ( ( { 9{ RG_zz_7_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_7_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_7_en = ( RG_zz_7_t_c1 | RG_zz_7_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_7_en )
		RG_zz_7 <= RG_zz_7_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_8_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h09 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_8_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h09 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_8_t = ( ( { 9{ RG_zz_8_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_8_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_8_en = ( RG_zz_8_t_c1 | RG_zz_8_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_8_en )
		RG_zz_8 <= RG_zz_8_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_9_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h0a ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_9_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h0a ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_9_t = ( ( { 9{ RG_zz_9_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_9_t_c2 } } & M_184 )	// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_9_en = ( RG_zz_9_t_c1 | RG_zz_9_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_9_en )
		RG_zz_9 <= RG_zz_9_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_10_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h0b ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_10_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h0b ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_10_t = ( ( { 9{ RG_zz_10_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_10_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_10_en = ( RG_zz_10_t_c1 | RG_zz_10_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_10_en )
		RG_zz_10 <= RG_zz_10_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_11_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h0c ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_11_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h0c ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_11_t = ( ( { 9{ RG_zz_11_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_11_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_11_en = ( RG_zz_11_t_c1 | RG_zz_11_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_11_en )
		RG_zz_11 <= RG_zz_11_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_12_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h0d ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_12_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h0d ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_12_t = ( ( { 9{ RG_zz_12_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_12_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_12_en = ( RG_zz_12_t_c1 | RG_zz_12_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_12_en )
		RG_zz_12 <= RG_zz_12_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_13_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h0e ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_13_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h0e ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_13_t = ( ( { 9{ RG_zz_13_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_13_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_13_en = ( RG_zz_13_t_c1 | RG_zz_13_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_13_en )
		RG_zz_13 <= RG_zz_13_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_14_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h0f ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_14_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h0f ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_14_t = ( ( { 9{ RG_zz_14_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_14_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_14_en = ( RG_zz_14_t_c1 | RG_zz_14_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_14_en )
		RG_zz_14 <= RG_zz_14_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_15_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h10 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_15_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h10 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_15_t = ( ( { 9{ RG_zz_15_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_15_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_15_en = ( RG_zz_15_t_c1 | RG_zz_15_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_15_en )
		RG_zz_15 <= RG_zz_15_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_16_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h11 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_16_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h11 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_16_t = ( ( { 9{ RG_zz_16_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_16_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_16_en = ( RG_zz_16_t_c1 | RG_zz_16_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_16_en )
		RG_zz_16 <= RG_zz_16_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_17_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h12 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_17_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h12 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_17_t = ( ( { 9{ RG_zz_17_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_17_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_17_en = ( RG_zz_17_t_c1 | RG_zz_17_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_17_en )
		RG_zz_17 <= RG_zz_17_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_18_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h13 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_18_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h13 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_18_t = ( ( { 9{ RG_zz_18_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_18_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_18_en = ( RG_zz_18_t_c1 | RG_zz_18_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_18_en )
		RG_zz_18 <= RG_zz_18_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_19_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h14 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_19_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h14 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_19_t = ( ( { 9{ RG_zz_19_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_19_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_19_en = ( RG_zz_19_t_c1 | RG_zz_19_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_19_en )
		RG_zz_19 <= RG_zz_19_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_20_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h15 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_20_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h15 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_20_t = ( ( { 9{ RG_zz_20_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_20_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_20_en = ( RG_zz_20_t_c1 | RG_zz_20_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_20_en )
		RG_zz_20 <= RG_zz_20_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_21_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h16 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_21_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h16 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_21_t = ( ( { 9{ RG_zz_21_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_21_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_21_en = ( RG_zz_21_t_c1 | RG_zz_21_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_21_en )
		RG_zz_21 <= RG_zz_21_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_22_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h17 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_22_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h17 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_22_t = ( ( { 9{ RG_zz_22_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_22_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_22_en = ( RG_zz_22_t_c1 | RG_zz_22_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_22_en )
		RG_zz_22 <= RG_zz_22_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_23_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h18 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_23_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h18 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_23_t = ( ( { 9{ RG_zz_23_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_23_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_23_en = ( RG_zz_23_t_c1 | RG_zz_23_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_23_en )
		RG_zz_23 <= RG_zz_23_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_24_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h19 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_24_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h19 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_24_t = ( ( { 9{ RG_zz_24_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_24_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_24_en = ( RG_zz_24_t_c1 | RG_zz_24_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_24_en )
		RG_zz_24 <= RG_zz_24_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_25_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h1a ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_25_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h1a ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_25_t = ( ( { 9{ RG_zz_25_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_25_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_25_en = ( RG_zz_25_t_c1 | RG_zz_25_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_25_en )
		RG_zz_25 <= RG_zz_25_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_26_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h1b ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_26_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h1b ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_26_t = ( ( { 9{ RG_zz_26_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_26_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_26_en = ( RG_zz_26_t_c1 | RG_zz_26_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_26_en )
		RG_zz_26 <= RG_zz_26_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_27_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h1c ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_27_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h1c ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_27_t = ( ( { 9{ RG_zz_27_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_27_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_27_en = ( RG_zz_27_t_c1 | RG_zz_27_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_27_en )
		RG_zz_27 <= RG_zz_27_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_28_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h1d ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_28_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h1d ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_28_t = ( ( { 9{ RG_zz_28_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_28_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_28_en = ( RG_zz_28_t_c1 | RG_zz_28_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_28_en )
		RG_zz_28 <= RG_zz_28_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_29_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h1e ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_29_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h1e ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_29_t = ( ( { 9{ RG_zz_29_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_29_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_29_en = ( RG_zz_29_t_c1 | RG_zz_29_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_29_en )
		RG_zz_29 <= RG_zz_29_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_30_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h1f ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_30_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h1f ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_30_t = ( ( { 9{ RG_zz_30_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_30_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_30_en = ( RG_zz_30_t_c1 | RG_zz_30_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_30_en )
		RG_zz_30 <= RG_zz_30_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_31_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h20 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_31_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h20 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_31_t = ( ( { 9{ RG_zz_31_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_31_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_31_en = ( RG_zz_31_t_c1 | RG_zz_31_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_31_en )
		RG_zz_31 <= RG_zz_31_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_32_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h21 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_32_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h21 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_32_t = ( ( { 9{ RG_zz_32_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_32_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_32_en = ( RG_zz_32_t_c1 | RG_zz_32_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_32_en )
		RG_zz_32 <= RG_zz_32_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_33_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h22 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_33_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h22 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_33_t = ( ( { 9{ RG_zz_33_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_33_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_33_en = ( RG_zz_33_t_c1 | RG_zz_33_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_33_en )
		RG_zz_33 <= RG_zz_33_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_34_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h23 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_34_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h23 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_34_t = ( ( { 9{ RG_zz_34_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_34_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_34_en = ( RG_zz_34_t_c1 | RG_zz_34_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_34_en )
		RG_zz_34 <= RG_zz_34_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_35_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h24 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_35_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h24 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_35_t = ( ( { 9{ RG_zz_35_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_35_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_35_en = ( RG_zz_35_t_c1 | RG_zz_35_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_35_en )
		RG_zz_35 <= RG_zz_35_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_36_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h25 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_36_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h25 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_36_t = ( ( { 9{ RG_zz_36_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_36_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_36_en = ( RG_zz_36_t_c1 | RG_zz_36_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_36_en )
		RG_zz_36 <= RG_zz_36_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_37_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h26 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_37_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h26 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_37_t = ( ( { 9{ RG_zz_37_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_37_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_37_en = ( RG_zz_37_t_c1 | RG_zz_37_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_37_en )
		RG_zz_37 <= RG_zz_37_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_38_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h27 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_38_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h27 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_38_t = ( ( { 9{ RG_zz_38_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_38_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_38_en = ( RG_zz_38_t_c1 | RG_zz_38_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_38_en )
		RG_zz_38 <= RG_zz_38_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_39_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h28 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_39_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h28 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_39_t = ( ( { 9{ RG_zz_39_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_39_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_39_en = ( RG_zz_39_t_c1 | RG_zz_39_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_39_en )
		RG_zz_39 <= RG_zz_39_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_40_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h29 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_40_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h29 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_40_t = ( ( { 9{ RG_zz_40_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_40_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_40_en = ( RG_zz_40_t_c1 | RG_zz_40_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_40_en )
		RG_zz_40 <= RG_zz_40_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_41_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h2a ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_41_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h2a ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_41_t = ( ( { 9{ RG_zz_41_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_41_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_41_en = ( RG_zz_41_t_c1 | RG_zz_41_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_41_en )
		RG_zz_41 <= RG_zz_41_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_42_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h2b ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_42_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h2b ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_42_t = ( ( { 9{ RG_zz_42_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_42_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_42_en = ( RG_zz_42_t_c1 | RG_zz_42_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_42_en )
		RG_zz_42 <= RG_zz_42_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_43_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h2c ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_43_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h2c ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_43_t = ( ( { 9{ RG_zz_43_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_43_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_43_en = ( RG_zz_43_t_c1 | RG_zz_43_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_43_en )
		RG_zz_43 <= RG_zz_43_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_44_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h2d ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_44_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h2d ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_44_t = ( ( { 9{ RG_zz_44_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_44_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_44_en = ( RG_zz_44_t_c1 | RG_zz_44_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_44_en )
		RG_zz_44 <= RG_zz_44_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_45_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h2e ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_45_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h2e ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_45_t = ( ( { 9{ RG_zz_45_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_45_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_45_en = ( RG_zz_45_t_c1 | RG_zz_45_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_45_en )
		RG_zz_45 <= RG_zz_45_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_46_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h2f ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_46_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h2f ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_46_t = ( ( { 9{ RG_zz_46_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_46_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_46_en = ( RG_zz_46_t_c1 | RG_zz_46_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_46_en )
		RG_zz_46 <= RG_zz_46_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_47_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h30 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_47_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h30 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_47_t = ( ( { 9{ RG_zz_47_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_47_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_47_en = ( RG_zz_47_t_c1 | RG_zz_47_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_47_en )
		RG_zz_47 <= RG_zz_47_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_48_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h31 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_48_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h31 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_48_t = ( ( { 9{ RG_zz_48_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_48_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_48_en = ( RG_zz_48_t_c1 | RG_zz_48_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_48_en )
		RG_zz_48 <= RG_zz_48_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_49_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h32 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_49_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h32 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_49_t = ( ( { 9{ RG_zz_49_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_49_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_49_en = ( RG_zz_49_t_c1 | RG_zz_49_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_49_en )
		RG_zz_49 <= RG_zz_49_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_50_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h33 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_50_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h33 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_50_t = ( ( { 9{ RG_zz_50_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_50_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_50_en = ( RG_zz_50_t_c1 | RG_zz_50_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_50_en )
		RG_zz_50 <= RG_zz_50_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_51_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h34 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_51_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h34 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_51_t = ( ( { 9{ RG_zz_51_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_51_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_51_en = ( RG_zz_51_t_c1 | RG_zz_51_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_51_en )
		RG_zz_51 <= RG_zz_51_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_52_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h35 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_52_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h35 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_52_t = ( ( { 9{ RG_zz_52_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_52_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_52_en = ( RG_zz_52_t_c1 | RG_zz_52_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_52_en )
		RG_zz_52 <= RG_zz_52_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_53_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h36 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_53_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h36 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_53_t = ( ( { 9{ RG_zz_53_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_53_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_53_en = ( RG_zz_53_t_c1 | RG_zz_53_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_53_en )
		RG_zz_53 <= RG_zz_53_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_54_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h37 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_54_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h37 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_54_t = ( ( { 9{ RG_zz_54_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_54_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_54_en = ( RG_zz_54_t_c1 | RG_zz_54_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_54_en )
		RG_zz_54 <= RG_zz_54_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_55_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h38 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_55_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h38 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_55_t = ( ( { 9{ RG_zz_55_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_55_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_55_en = ( RG_zz_55_t_c1 | RG_zz_55_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_55_en )
		RG_zz_55 <= RG_zz_55_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_56_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h39 ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_56_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h39 ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_56_t = ( ( { 9{ RG_zz_56_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_56_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_56_en = ( RG_zz_56_t_c1 | RG_zz_56_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_56_en )
		RG_zz_56 <= RG_zz_56_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_57_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h3a ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_57_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h3a ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_57_t = ( ( { 9{ RG_zz_57_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_57_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_57_en = ( RG_zz_57_t_c1 | RG_zz_57_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_57_en )
		RG_zz_57 <= RG_zz_57_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_58_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h3b ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_58_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h3b ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_58_t = ( ( { 9{ RG_zz_58_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_58_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_58_en = ( RG_zz_58_t_c1 | RG_zz_58_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_58_en )
		RG_zz_58 <= RG_zz_58_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_59_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h3c ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_59_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h3c ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_59_t = ( ( { 9{ RG_zz_59_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_59_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_59_en = ( RG_zz_59_t_c1 | RG_zz_59_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_59_en )
		RG_zz_59 <= RG_zz_59_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_60_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h3d ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_60_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h3d ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_60_t = ( ( { 9{ RG_zz_60_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_60_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_60_en = ( RG_zz_60_t_c1 | RG_zz_60_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_60_en )
		RG_zz_60 <= RG_zz_60_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_61_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h3e ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_61_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h3e ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_61_t = ( ( { 9{ RG_zz_61_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_61_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_61_en = ( RG_zz_61_t_c1 | RG_zz_61_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_61_en )
		RG_zz_61 <= RG_zz_61_t ;	// line#=../rle.cpp:111,142
always @ ( RG_k_1 or U_87 or M_184 or RG_k or U_05 )	// line#=../rle.cpp:111,142
	begin
	RG_zz_62_t_c1 = ( U_05 & ( ~|( RG_k ^ 6'h3f ) ) ) ;	// line#=../rle.cpp:111
	RG_zz_62_t_c2 = ( U_87 & ( ~|( RG_k_1 [5:0] ^ 6'h3f ) ) ) ;	// line#=../rle.cpp:142
	RG_zz_62_t = ( ( { 9{ RG_zz_62_t_c1 } } & M_184 )	// line#=../rle.cpp:111
		| ( { 9{ RG_zz_62_t_c2 } } & M_184 )		// line#=../rle.cpp:142
		) ;
	end
assign	RG_zz_62_en = ( RG_zz_62_t_c1 | RG_zz_62_t_c2 ) ;	// line#=../rle.cpp:111,142
always @ ( posedge clk )	// line#=../rle.cpp:111,142
	if ( RG_zz_62_en )
		RG_zz_62 <= RG_zz_62_t ;	// line#=../rle.cpp:111,142
always @ ( FF_j or ST1_07d or incr4s1ot or ST1_02d or ST1_01d )
	RG_j_t = ( ( { 4{ ST1_01d } } & 4'hf /*-4'h1*/ )	// line#=../rle.cpp:34
		| ( { 4{ ST1_02d } } & incr4s1ot )		// line#=../rle.cpp:34
		| ( { 4{ ST1_07d } } & { 3'h0 , FF_j } ) ) ;
always @ ( posedge clk )
	RG_j <= RG_j_t ;	// line#=../rle.cpp:34
assign	M_182 = ( ST1_02d | ST1_05d ) ;
always @ ( U_06 )
	TR_01 = ( { 3{ U_06 } } & 3'h7 )	// line#=../rle.cpp:134
		 ;	// line#=../rle.cpp:59,105
always @ ( decr32s1ot or U_165 or U_83 or incr32s2ot or ST1_06d or U_166 or U_163 or 
	U_84 or U_81 or TR_01 or U_06 or M_182 )
	begin
	RG_i_k_01_t_c1 = ( M_182 | U_06 ) ;	// line#=../rle.cpp:59,105,134
	RG_i_k_01_t_c2 = ( ( ( ( U_81 | U_84 ) | U_163 ) | U_166 ) | ST1_06d ) ;	// line#=../rle.cpp:64,119,129,150,160
	RG_i_k_01_t_c3 = ( U_83 | U_165 ) ;	// line#=../rle.cpp:124,155
	RG_i_k_01_t = ( ( { 32{ RG_i_k_01_t_c1 } } & { 29'h00000000 , TR_01 } )	// line#=../rle.cpp:59,105,134
		| ( { 32{ RG_i_k_01_t_c2 } } & incr32s2ot )			// line#=../rle.cpp:64,119,129,150,160
		| ( { 32{ RG_i_k_01_t_c3 } } & decr32s1ot )			// line#=../rle.cpp:124,155
		) ;
	end
assign	RG_i_k_01_en = ( RG_i_k_01_t_c1 | RG_i_k_01_t_c2 | RG_i_k_01_t_c3 ) ;
always @ ( posedge clk )
	if ( RG_i_k_01_en )
		RG_i_k_01 <= RG_i_k_01_t ;	// line#=../rle.cpp:59,64,105,119,124,129
						// ,134,150,155,160
always @ ( FF_i or U_88 or U_06 )
	TR_02 = ( ( { 1{ U_06 } } & 1'h1 )	// line#=../rle.cpp:135
		| ( { 1{ U_88 } } & FF_i ) ) ;	// line#=../rle.cpp:105
always @ ( decr32s2ot or U_166 or U_84 or incr32s1ot or C_08 or ST1_06d or U_318 or 
	U_165 or U_161 or U_83 or U_79 or TR_02 or U_88 or M_181 )	// line#=../rle.cpp:61,62
	begin
	RG_i_j_01_t_c1 = ( M_181 | U_88 ) ;	// line#=../rle.cpp:105,135
	RG_i_j_01_t_c2 = ( ( ( ( ( U_79 | U_83 ) | U_161 ) | U_165 ) | U_318 ) | 
		( ST1_06d & C_08 ) ) ;	// line#=../rle.cpp:61,62,63,74,114,125
					// ,145,156
	RG_i_j_01_t_c3 = ( U_84 | U_166 ) ;	// line#=../rle.cpp:130,161
	RG_i_j_01_t = ( ( { 32{ RG_i_j_01_t_c1 } } & { 31'h00000000 , TR_02 } )	// line#=../rle.cpp:105,135
		| ( { 32{ RG_i_j_01_t_c2 } } & incr32s1ot )			// line#=../rle.cpp:61,62,63,74,114,125
										// ,145,156
		| ( { 32{ RG_i_j_01_t_c3 } } & decr32s2ot )			// line#=../rle.cpp:130,161
		) ;
	end
assign	RG_i_j_01_en = ( RG_i_j_01_t_c1 | RG_i_j_01_t_c2 | RG_i_j_01_t_c3 ) ;	// line#=../rle.cpp:61,62
always @ ( posedge clk )	// line#=../rle.cpp:61,62
	if ( RG_i_j_01_en )
		RG_i_j_01 <= RG_i_j_01_t ;	// line#=../rle.cpp:61,62,63,74,105,114
						// ,125,130,135,145,156,161
always @ ( M_16_t or rl_a05_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h01 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h02 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h03 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h04 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h05 :
		RG_quantized_block_rl_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h06 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h07 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h08 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h09 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h0a :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h0b :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h0c :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h0d :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h0e :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h0f :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h10 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h11 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h12 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h13 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h14 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h15 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h16 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h17 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h18 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h19 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h1a :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h1b :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h1c :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h1d :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h1e :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h1f :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h20 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h21 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h22 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h23 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h24 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h25 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h26 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h27 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h28 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h29 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h2a :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h2b :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h2c :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h2d :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h2e :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h2f :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h30 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h31 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h32 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h33 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h34 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h35 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h36 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h37 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h38 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h39 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h3a :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h3b :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h3c :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h3d :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h3e :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h3f :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h40 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h41 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h42 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h43 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h44 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h45 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h46 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h47 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h48 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h49 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h4a :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h4b :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h4c :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h4d :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h4e :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h4f :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h50 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h51 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h52 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h53 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h54 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h55 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h56 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h57 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h58 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h59 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h5a :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h5b :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h5c :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h5d :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h5e :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h5f :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h60 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h61 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h62 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h63 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h64 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h65 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h66 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h67 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h68 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h69 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h6a :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h6b :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h6c :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h6d :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h6e :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h6f :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h70 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h71 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h72 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h73 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h74 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h75 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h76 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h77 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h78 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h79 :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h7a :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h7b :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h7c :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h7d :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h7e :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	7'h7f :
		RG_quantized_block_rl_t1 = rl_a05_t8 ;
	default :
		RG_quantized_block_rl_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_t1 or U_318 or TR_260 or U_317 or RG_rl_7 or ST1_07d or 
	RG_rl_131 or U_88 or jpeg_in_a00 or U_01 or RG_quantized_block_rl_2 or ST1_01d )
	RG_quantized_block_rl_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_2 )
		| ( { 9{ U_01 } } & jpeg_in_a00 )		// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_131 )
		| ( { 9{ ST1_07d } } & RG_rl_7 )
		| ( { 9{ U_317 } } & TR_260 )			// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_en )
		RG_quantized_block_rl <= RG_quantized_block_rl_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a07_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h01 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h02 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h03 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h04 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h05 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h06 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h07 :
		RG_quantized_block_rl_1_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h08 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h09 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h0a :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h0b :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h0c :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h0d :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h0e :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h0f :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h10 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h11 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h12 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h13 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h14 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h15 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h16 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h17 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h18 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h19 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h1a :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h1b :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h1c :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h1d :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h1e :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h1f :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h20 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h21 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h22 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h23 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h24 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h25 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h26 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h27 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h28 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h29 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h2a :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h2b :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h2c :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h2d :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h2e :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h2f :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h30 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h31 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h32 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h33 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h34 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h35 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h36 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h37 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h38 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h39 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h3a :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h3b :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h3c :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h3d :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h3e :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h3f :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h40 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h41 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h42 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h43 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h44 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h45 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h46 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h47 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h48 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h49 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h4a :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h4b :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h4c :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h4d :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h4e :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h4f :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h50 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h51 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h52 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h53 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h54 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h55 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h56 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h57 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h58 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h59 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h5a :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h5b :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h5c :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h5d :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h5e :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h5f :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h60 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h61 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h62 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h63 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h64 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h65 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h66 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h67 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h68 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h69 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h6a :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h6b :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h6c :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h6d :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h6e :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h6f :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h70 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h71 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h72 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h73 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h74 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h75 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h76 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h77 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h78 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h79 :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h7a :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h7b :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h7c :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h7d :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h7e :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	7'h7f :
		RG_quantized_block_rl_1_t1 = rl_a07_t8 ;
	default :
		RG_quantized_block_rl_1_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_1_t1 or U_318 or TR_258 or U_317 or RG_rl_9 or 
	ST1_07d or RG_rl_7 or U_88 or jpeg_in_a01 or U_01 or RG_quantized_block_rl_3 or 
	ST1_01d )
	RG_quantized_block_rl_1_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_3 )
		| ( { 9{ U_01 } } & jpeg_in_a01 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_7 )
		| ( { 9{ ST1_07d } } & RG_rl_9 )
		| ( { 9{ U_317 } } & TR_258 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_1_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_1_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_1_en )
		RG_quantized_block_rl_1 <= RG_quantized_block_rl_1_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a09_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h01 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h02 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h03 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h04 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h05 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h06 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h07 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h08 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h09 :
		RG_quantized_block_rl_2_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h0a :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h0b :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h0c :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h0d :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h0e :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h0f :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h10 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h11 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h12 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h13 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h14 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h15 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h16 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h17 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h18 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h19 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h1a :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h1b :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h1c :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h1d :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h1e :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h1f :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h20 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h21 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h22 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h23 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h24 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h25 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h26 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h27 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h28 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h29 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h2a :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h2b :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h2c :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h2d :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h2e :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h2f :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h30 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h31 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h32 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h33 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h34 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h35 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h36 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h37 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h38 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h39 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h3a :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h3b :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h3c :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h3d :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h3e :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h3f :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h40 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h41 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h42 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h43 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h44 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h45 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h46 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h47 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h48 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h49 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h4a :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h4b :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h4c :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h4d :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h4e :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h4f :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h50 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h51 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h52 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h53 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h54 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h55 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h56 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h57 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h58 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h59 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h5a :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h5b :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h5c :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h5d :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h5e :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h5f :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h60 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h61 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h62 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h63 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h64 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h65 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h66 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h67 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h68 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h69 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h6a :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h6b :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h6c :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h6d :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h6e :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h6f :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h70 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h71 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h72 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h73 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h74 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h75 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h76 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h77 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h78 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h79 :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h7a :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h7b :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h7c :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h7d :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h7e :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	7'h7f :
		RG_quantized_block_rl_2_t1 = rl_a09_t8 ;
	default :
		RG_quantized_block_rl_2_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_2_t1 or U_318 or TR_256 or U_317 or RG_rl_11 or 
	ST1_07d or RG_rl_9 or U_88 or jpeg_in_a02 or U_01 or RG_quantized_block_rl_4 or 
	ST1_01d )
	RG_quantized_block_rl_2_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_4 )
		| ( { 9{ U_01 } } & jpeg_in_a02 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_9 )
		| ( { 9{ ST1_07d } } & RG_rl_11 )
		| ( { 9{ U_317 } } & TR_256 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_2_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_2_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_2_en )
		RG_quantized_block_rl_2 <= RG_quantized_block_rl_2_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a11_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h01 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h02 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h03 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h04 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h05 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h06 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h07 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h08 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h09 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h0a :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h0b :
		RG_quantized_block_rl_3_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h0c :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h0d :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h0e :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h0f :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h10 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h11 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h12 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h13 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h14 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h15 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h16 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h17 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h18 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h19 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h1a :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h1b :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h1c :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h1d :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h1e :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h1f :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h20 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h21 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h22 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h23 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h24 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h25 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h26 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h27 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h28 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h29 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h2a :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h2b :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h2c :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h2d :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h2e :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h2f :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h30 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h31 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h32 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h33 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h34 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h35 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h36 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h37 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h38 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h39 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h3a :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h3b :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h3c :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h3d :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h3e :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h3f :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h40 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h41 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h42 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h43 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h44 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h45 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h46 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h47 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h48 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h49 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h4a :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h4b :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h4c :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h4d :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h4e :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h4f :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h50 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h51 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h52 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h53 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h54 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h55 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h56 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h57 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h58 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h59 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h5a :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h5b :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h5c :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h5d :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h5e :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h5f :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h60 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h61 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h62 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h63 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h64 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h65 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h66 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h67 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h68 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h69 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h6a :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h6b :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h6c :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h6d :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h6e :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h6f :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h70 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h71 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h72 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h73 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h74 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h75 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h76 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h77 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h78 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h79 :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h7a :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h7b :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h7c :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h7d :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h7e :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	7'h7f :
		RG_quantized_block_rl_3_t1 = rl_a11_t8 ;
	default :
		RG_quantized_block_rl_3_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_3_t1 or U_318 or TR_254 or U_317 or RG_rl_13 or 
	ST1_07d or RG_rl_11 or U_88 or jpeg_in_a03 or U_01 or RG_quantized_block_rl_5 or 
	ST1_01d )
	RG_quantized_block_rl_3_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_5 )
		| ( { 9{ U_01 } } & jpeg_in_a03 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_11 )
		| ( { 9{ ST1_07d } } & RG_rl_13 )
		| ( { 9{ U_317 } } & TR_254 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_3_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_3_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_3_en )
		RG_quantized_block_rl_3 <= RG_quantized_block_rl_3_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a13_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h01 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h02 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h03 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h04 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h05 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h06 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h07 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h08 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h09 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h0a :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h0b :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h0c :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h0d :
		RG_quantized_block_rl_4_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h0e :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h0f :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h10 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h11 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h12 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h13 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h14 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h15 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h16 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h17 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h18 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h19 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h1a :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h1b :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h1c :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h1d :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h1e :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h1f :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h20 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h21 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h22 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h23 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h24 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h25 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h26 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h27 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h28 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h29 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h2a :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h2b :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h2c :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h2d :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h2e :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h2f :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h30 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h31 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h32 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h33 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h34 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h35 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h36 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h37 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h38 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h39 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h3a :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h3b :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h3c :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h3d :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h3e :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h3f :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h40 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h41 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h42 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h43 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h44 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h45 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h46 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h47 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h48 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h49 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h4a :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h4b :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h4c :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h4d :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h4e :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h4f :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h50 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h51 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h52 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h53 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h54 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h55 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h56 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h57 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h58 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h59 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h5a :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h5b :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h5c :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h5d :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h5e :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h5f :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h60 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h61 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h62 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h63 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h64 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h65 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h66 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h67 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h68 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h69 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h6a :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h6b :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h6c :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h6d :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h6e :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h6f :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h70 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h71 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h72 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h73 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h74 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h75 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h76 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h77 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h78 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h79 :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h7a :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h7b :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h7c :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h7d :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h7e :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	7'h7f :
		RG_quantized_block_rl_4_t1 = rl_a13_t8 ;
	default :
		RG_quantized_block_rl_4_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_4_t1 or U_318 or TR_252 or U_317 or RG_rl_15 or 
	ST1_07d or RG_rl_13 or U_88 or jpeg_in_a04 or U_01 or RG_quantized_block_rl_6 or 
	ST1_01d )
	RG_quantized_block_rl_4_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_6 )
		| ( { 9{ U_01 } } & jpeg_in_a04 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_13 )
		| ( { 9{ ST1_07d } } & RG_rl_15 )
		| ( { 9{ U_317 } } & TR_252 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_4_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_4_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_4_en )
		RG_quantized_block_rl_4 <= RG_quantized_block_rl_4_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a15_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h01 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h02 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h03 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h04 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h05 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h06 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h07 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h08 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h09 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h0a :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h0b :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h0c :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h0d :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h0e :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h0f :
		RG_quantized_block_rl_5_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h10 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h11 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h12 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h13 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h14 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h15 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h16 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h17 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h18 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h19 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h1a :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h1b :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h1c :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h1d :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h1e :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h1f :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h20 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h21 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h22 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h23 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h24 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h25 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h26 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h27 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h28 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h29 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h2a :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h2b :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h2c :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h2d :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h2e :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h2f :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h30 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h31 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h32 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h33 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h34 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h35 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h36 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h37 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h38 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h39 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h3a :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h3b :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h3c :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h3d :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h3e :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h3f :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h40 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h41 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h42 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h43 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h44 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h45 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h46 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h47 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h48 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h49 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h4a :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h4b :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h4c :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h4d :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h4e :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h4f :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h50 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h51 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h52 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h53 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h54 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h55 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h56 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h57 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h58 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h59 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h5a :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h5b :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h5c :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h5d :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h5e :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h5f :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h60 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h61 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h62 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h63 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h64 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h65 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h66 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h67 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h68 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h69 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h6a :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h6b :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h6c :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h6d :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h6e :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h6f :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h70 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h71 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h72 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h73 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h74 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h75 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h76 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h77 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h78 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h79 :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h7a :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h7b :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h7c :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h7d :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h7e :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	7'h7f :
		RG_quantized_block_rl_5_t1 = rl_a15_t8 ;
	default :
		RG_quantized_block_rl_5_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_5_t1 or U_318 or TR_250 or U_317 or RG_rl_17 or 
	ST1_07d or RG_rl_15 or U_88 or jpeg_in_a05 or U_01 or RG_quantized_block_rl_7 or 
	ST1_01d )
	RG_quantized_block_rl_5_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_7 )
		| ( { 9{ U_01 } } & jpeg_in_a05 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_15 )
		| ( { 9{ ST1_07d } } & RG_rl_17 )
		| ( { 9{ U_317 } } & TR_250 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_5_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_5_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_5_en )
		RG_quantized_block_rl_5 <= RG_quantized_block_rl_5_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a17_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h01 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h02 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h03 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h04 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h05 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h06 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h07 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h08 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h09 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h0a :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h0b :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h0c :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h0d :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h0e :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h0f :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h10 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h11 :
		RG_quantized_block_rl_6_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h12 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h13 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h14 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h15 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h16 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h17 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h18 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h19 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h1a :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h1b :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h1c :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h1d :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h1e :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h1f :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h20 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h21 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h22 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h23 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h24 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h25 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h26 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h27 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h28 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h29 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h2a :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h2b :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h2c :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h2d :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h2e :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h2f :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h30 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h31 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h32 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h33 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h34 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h35 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h36 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h37 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h38 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h39 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h3a :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h3b :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h3c :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h3d :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h3e :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h3f :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h40 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h41 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h42 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h43 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h44 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h45 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h46 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h47 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h48 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h49 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h4a :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h4b :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h4c :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h4d :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h4e :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h4f :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h50 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h51 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h52 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h53 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h54 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h55 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h56 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h57 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h58 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h59 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h5a :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h5b :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h5c :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h5d :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h5e :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h5f :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h60 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h61 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h62 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h63 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h64 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h65 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h66 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h67 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h68 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h69 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h6a :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h6b :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h6c :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h6d :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h6e :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h6f :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h70 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h71 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h72 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h73 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h74 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h75 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h76 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h77 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h78 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h79 :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h7a :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h7b :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h7c :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h7d :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h7e :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	7'h7f :
		RG_quantized_block_rl_6_t1 = rl_a17_t8 ;
	default :
		RG_quantized_block_rl_6_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_6_t1 or U_318 or TR_248 or U_317 or RG_rl_19 or 
	ST1_07d or RG_rl_17 or U_88 or jpeg_in_a06 or U_01 or RG_quantized_block_rl_8 or 
	ST1_01d )
	RG_quantized_block_rl_6_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_8 )
		| ( { 9{ U_01 } } & jpeg_in_a06 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_17 )
		| ( { 9{ ST1_07d } } & RG_rl_19 )
		| ( { 9{ U_317 } } & TR_248 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_6_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_6_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_6_en )
		RG_quantized_block_rl_6 <= RG_quantized_block_rl_6_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a19_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h01 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h02 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h03 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h04 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h05 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h06 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h07 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h08 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h09 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h0a :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h0b :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h0c :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h0d :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h0e :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h0f :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h10 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h11 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h12 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h13 :
		RG_quantized_block_rl_7_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h14 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h15 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h16 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h17 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h18 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h19 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h1a :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h1b :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h1c :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h1d :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h1e :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h1f :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h20 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h21 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h22 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h23 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h24 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h25 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h26 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h27 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h28 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h29 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h2a :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h2b :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h2c :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h2d :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h2e :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h2f :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h30 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h31 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h32 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h33 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h34 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h35 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h36 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h37 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h38 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h39 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h3a :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h3b :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h3c :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h3d :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h3e :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h3f :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h40 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h41 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h42 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h43 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h44 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h45 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h46 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h47 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h48 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h49 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h4a :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h4b :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h4c :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h4d :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h4e :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h4f :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h50 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h51 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h52 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h53 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h54 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h55 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h56 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h57 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h58 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h59 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h5a :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h5b :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h5c :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h5d :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h5e :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h5f :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h60 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h61 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h62 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h63 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h64 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h65 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h66 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h67 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h68 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h69 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h6a :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h6b :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h6c :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h6d :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h6e :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h6f :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h70 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h71 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h72 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h73 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h74 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h75 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h76 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h77 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h78 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h79 :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h7a :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h7b :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h7c :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h7d :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h7e :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	7'h7f :
		RG_quantized_block_rl_7_t1 = rl_a19_t8 ;
	default :
		RG_quantized_block_rl_7_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_7_t1 or U_318 or TR_246 or U_317 or RG_rl_21 or 
	ST1_07d or RG_rl_19 or U_88 or jpeg_in_a07 or U_01 or RG_quantized_block_rl_9 or 
	ST1_01d )
	RG_quantized_block_rl_7_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_9 )
		| ( { 9{ U_01 } } & jpeg_in_a07 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_19 )
		| ( { 9{ ST1_07d } } & RG_rl_21 )
		| ( { 9{ U_317 } } & TR_246 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_7_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_7_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_7_en )
		RG_quantized_block_rl_7 <= RG_quantized_block_rl_7_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a21_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h01 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h02 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h03 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h04 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h05 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h06 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h07 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h08 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h09 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h0a :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h0b :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h0c :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h0d :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h0e :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h0f :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h10 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h11 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h12 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h13 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h14 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h15 :
		RG_quantized_block_rl_8_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h16 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h17 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h18 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h19 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h1a :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h1b :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h1c :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h1d :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h1e :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h1f :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h20 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h21 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h22 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h23 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h24 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h25 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h26 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h27 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h28 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h29 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h2a :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h2b :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h2c :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h2d :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h2e :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h2f :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h30 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h31 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h32 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h33 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h34 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h35 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h36 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h37 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h38 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h39 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h3a :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h3b :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h3c :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h3d :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h3e :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h3f :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h40 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h41 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h42 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h43 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h44 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h45 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h46 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h47 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h48 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h49 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h4a :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h4b :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h4c :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h4d :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h4e :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h4f :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h50 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h51 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h52 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h53 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h54 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h55 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h56 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h57 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h58 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h59 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h5a :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h5b :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h5c :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h5d :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h5e :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h5f :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h60 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h61 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h62 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h63 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h64 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h65 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h66 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h67 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h68 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h69 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h6a :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h6b :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h6c :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h6d :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h6e :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h6f :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h70 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h71 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h72 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h73 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h74 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h75 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h76 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h77 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h78 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h79 :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h7a :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h7b :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h7c :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h7d :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h7e :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	7'h7f :
		RG_quantized_block_rl_8_t1 = rl_a21_t8 ;
	default :
		RG_quantized_block_rl_8_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_8_t1 or U_318 or TR_244 or U_317 or RG_rl_23 or 
	ST1_07d or RG_rl_21 or U_88 or jpeg_in_a08 or U_01 or RG_quantized_block_rl_10 or 
	ST1_01d )
	RG_quantized_block_rl_8_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_10 )
		| ( { 9{ U_01 } } & jpeg_in_a08 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_21 )
		| ( { 9{ ST1_07d } } & RG_rl_23 )
		| ( { 9{ U_317 } } & TR_244 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_8_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_8_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_8_en )
		RG_quantized_block_rl_8 <= RG_quantized_block_rl_8_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a23_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h01 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h02 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h03 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h04 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h05 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h06 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h07 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h08 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h09 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h0a :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h0b :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h0c :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h0d :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h0e :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h0f :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h10 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h11 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h12 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h13 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h14 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h15 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h16 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h17 :
		RG_quantized_block_rl_9_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h18 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h19 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h1a :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h1b :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h1c :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h1d :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h1e :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h1f :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h20 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h21 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h22 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h23 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h24 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h25 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h26 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h27 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h28 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h29 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h2a :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h2b :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h2c :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h2d :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h2e :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h2f :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h30 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h31 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h32 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h33 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h34 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h35 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h36 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h37 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h38 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h39 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h3a :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h3b :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h3c :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h3d :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h3e :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h3f :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h40 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h41 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h42 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h43 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h44 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h45 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h46 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h47 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h48 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h49 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h4a :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h4b :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h4c :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h4d :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h4e :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h4f :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h50 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h51 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h52 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h53 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h54 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h55 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h56 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h57 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h58 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h59 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h5a :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h5b :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h5c :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h5d :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h5e :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h5f :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h60 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h61 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h62 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h63 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h64 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h65 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h66 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h67 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h68 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h69 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h6a :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h6b :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h6c :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h6d :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h6e :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h6f :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h70 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h71 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h72 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h73 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h74 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h75 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h76 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h77 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h78 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h79 :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h7a :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h7b :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h7c :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h7d :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h7e :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	7'h7f :
		RG_quantized_block_rl_9_t1 = rl_a23_t8 ;
	default :
		RG_quantized_block_rl_9_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_9_t1 or U_318 or TR_242 or U_317 or RG_rl_25 or 
	ST1_07d or RG_rl_23 or U_88 or jpeg_in_a09 or U_01 or RG_quantized_block_rl_11 or 
	ST1_01d )
	RG_quantized_block_rl_9_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_11 )
		| ( { 9{ U_01 } } & jpeg_in_a09 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_23 )
		| ( { 9{ ST1_07d } } & RG_rl_25 )
		| ( { 9{ U_317 } } & TR_242 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_9_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_9_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_9_en )
		RG_quantized_block_rl_9 <= RG_quantized_block_rl_9_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a25_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h01 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h02 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h03 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h04 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h05 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h06 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h07 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h08 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h09 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h0a :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h0b :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h0c :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h0d :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h0e :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h0f :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h10 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h11 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h12 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h13 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h14 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h15 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h16 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h17 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h18 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h19 :
		RG_quantized_block_rl_10_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h1a :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h1b :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h1c :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h1d :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h1e :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h1f :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h20 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h21 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h22 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h23 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h24 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h25 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h26 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h27 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h28 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h29 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h2a :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h2b :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h2c :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h2d :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h2e :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h2f :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h30 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h31 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h32 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h33 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h34 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h35 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h36 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h37 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h38 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h39 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h3a :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h3b :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h3c :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h3d :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h3e :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h3f :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h40 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h41 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h42 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h43 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h44 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h45 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h46 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h47 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h48 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h49 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h4a :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h4b :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h4c :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h4d :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h4e :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h4f :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h50 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h51 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h52 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h53 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h54 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h55 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h56 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h57 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h58 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h59 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h5a :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h5b :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h5c :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h5d :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h5e :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h5f :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h60 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h61 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h62 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h63 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h64 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h65 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h66 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h67 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h68 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h69 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h6a :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h6b :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h6c :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h6d :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h6e :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h6f :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h70 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h71 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h72 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h73 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h74 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h75 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h76 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h77 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h78 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h79 :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h7a :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h7b :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h7c :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h7d :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h7e :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	7'h7f :
		RG_quantized_block_rl_10_t1 = rl_a25_t8 ;
	default :
		RG_quantized_block_rl_10_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_10_t1 or U_318 or TR_240 or U_317 or RG_rl_27 or 
	ST1_07d or RG_rl_25 or U_88 or jpeg_in_a10 or U_01 or RG_quantized_block_rl_12 or 
	ST1_01d )
	RG_quantized_block_rl_10_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_12 )
		| ( { 9{ U_01 } } & jpeg_in_a10 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_25 )
		| ( { 9{ ST1_07d } } & RG_rl_27 )
		| ( { 9{ U_317 } } & TR_240 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_10_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_10_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_10_en )
		RG_quantized_block_rl_10 <= RG_quantized_block_rl_10_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a27_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h01 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h02 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h03 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h04 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h05 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h06 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h07 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h08 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h09 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h0a :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h0b :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h0c :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h0d :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h0e :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h0f :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h10 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h11 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h12 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h13 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h14 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h15 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h16 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h17 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h18 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h19 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h1a :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h1b :
		RG_quantized_block_rl_11_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h1c :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h1d :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h1e :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h1f :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h20 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h21 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h22 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h23 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h24 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h25 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h26 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h27 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h28 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h29 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h2a :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h2b :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h2c :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h2d :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h2e :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h2f :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h30 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h31 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h32 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h33 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h34 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h35 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h36 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h37 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h38 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h39 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h3a :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h3b :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h3c :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h3d :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h3e :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h3f :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h40 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h41 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h42 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h43 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h44 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h45 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h46 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h47 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h48 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h49 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h4a :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h4b :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h4c :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h4d :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h4e :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h4f :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h50 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h51 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h52 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h53 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h54 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h55 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h56 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h57 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h58 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h59 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h5a :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h5b :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h5c :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h5d :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h5e :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h5f :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h60 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h61 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h62 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h63 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h64 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h65 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h66 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h67 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h68 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h69 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h6a :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h6b :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h6c :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h6d :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h6e :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h6f :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h70 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h71 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h72 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h73 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h74 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h75 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h76 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h77 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h78 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h79 :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h7a :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h7b :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h7c :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h7d :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h7e :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	7'h7f :
		RG_quantized_block_rl_11_t1 = rl_a27_t8 ;
	default :
		RG_quantized_block_rl_11_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_11_t1 or U_318 or TR_238 or U_317 or RG_rl_29 or 
	ST1_07d or RG_rl_27 or U_88 or jpeg_in_a11 or U_01 or RG_quantized_block_rl_13 or 
	ST1_01d )
	RG_quantized_block_rl_11_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_13 )
		| ( { 9{ U_01 } } & jpeg_in_a11 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_27 )
		| ( { 9{ ST1_07d } } & RG_rl_29 )
		| ( { 9{ U_317 } } & TR_238 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_11_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_11_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_11_en )
		RG_quantized_block_rl_11 <= RG_quantized_block_rl_11_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a29_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h01 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h02 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h03 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h04 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h05 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h06 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h07 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h08 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h09 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h0a :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h0b :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h0c :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h0d :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h0e :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h0f :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h10 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h11 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h12 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h13 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h14 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h15 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h16 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h17 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h18 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h19 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h1a :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h1b :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h1c :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h1d :
		RG_quantized_block_rl_12_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h1e :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h1f :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h20 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h21 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h22 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h23 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h24 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h25 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h26 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h27 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h28 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h29 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h2a :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h2b :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h2c :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h2d :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h2e :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h2f :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h30 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h31 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h32 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h33 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h34 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h35 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h36 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h37 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h38 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h39 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h3a :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h3b :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h3c :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h3d :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h3e :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h3f :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h40 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h41 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h42 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h43 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h44 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h45 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h46 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h47 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h48 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h49 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h4a :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h4b :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h4c :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h4d :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h4e :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h4f :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h50 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h51 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h52 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h53 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h54 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h55 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h56 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h57 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h58 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h59 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h5a :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h5b :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h5c :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h5d :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h5e :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h5f :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h60 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h61 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h62 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h63 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h64 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h65 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h66 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h67 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h68 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h69 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h6a :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h6b :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h6c :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h6d :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h6e :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h6f :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h70 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h71 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h72 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h73 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h74 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h75 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h76 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h77 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h78 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h79 :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h7a :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h7b :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h7c :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h7d :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h7e :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	7'h7f :
		RG_quantized_block_rl_12_t1 = rl_a29_t8 ;
	default :
		RG_quantized_block_rl_12_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_12_t1 or U_318 or TR_236 or U_317 or RG_rl_31 or 
	ST1_07d or RG_rl_29 or U_88 or jpeg_in_a12 or U_01 or RG_quantized_block_rl_14 or 
	ST1_01d )
	RG_quantized_block_rl_12_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_14 )
		| ( { 9{ U_01 } } & jpeg_in_a12 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_29 )
		| ( { 9{ ST1_07d } } & RG_rl_31 )
		| ( { 9{ U_317 } } & TR_236 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_12_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_12_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_12_en )
		RG_quantized_block_rl_12 <= RG_quantized_block_rl_12_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a31_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h01 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h02 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h03 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h04 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h05 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h06 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h07 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h08 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h09 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h0a :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h0b :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h0c :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h0d :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h0e :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h0f :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h10 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h11 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h12 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h13 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h14 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h15 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h16 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h17 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h18 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h19 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h1a :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h1b :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h1c :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h1d :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h1e :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h1f :
		RG_quantized_block_rl_13_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h20 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h21 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h22 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h23 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h24 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h25 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h26 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h27 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h28 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h29 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h2a :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h2b :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h2c :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h2d :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h2e :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h2f :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h30 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h31 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h32 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h33 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h34 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h35 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h36 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h37 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h38 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h39 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h3a :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h3b :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h3c :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h3d :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h3e :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h3f :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h40 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h41 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h42 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h43 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h44 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h45 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h46 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h47 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h48 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h49 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h4a :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h4b :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h4c :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h4d :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h4e :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h4f :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h50 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h51 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h52 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h53 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h54 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h55 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h56 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h57 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h58 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h59 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h5a :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h5b :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h5c :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h5d :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h5e :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h5f :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h60 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h61 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h62 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h63 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h64 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h65 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h66 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h67 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h68 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h69 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h6a :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h6b :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h6c :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h6d :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h6e :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h6f :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h70 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h71 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h72 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h73 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h74 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h75 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h76 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h77 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h78 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h79 :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h7a :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h7b :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h7c :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h7d :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h7e :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	7'h7f :
		RG_quantized_block_rl_13_t1 = rl_a31_t8 ;
	default :
		RG_quantized_block_rl_13_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_13_t1 or U_318 or TR_234 or U_317 or RG_rl_33 or 
	ST1_07d or RG_rl_31 or U_88 or jpeg_in_a13 or U_01 or RG_quantized_block_rl_15 or 
	ST1_01d )
	RG_quantized_block_rl_13_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_15 )
		| ( { 9{ U_01 } } & jpeg_in_a13 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_31 )
		| ( { 9{ ST1_07d } } & RG_rl_33 )
		| ( { 9{ U_317 } } & TR_234 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_13_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_13_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_13_en )
		RG_quantized_block_rl_13 <= RG_quantized_block_rl_13_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a33_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h01 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h02 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h03 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h04 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h05 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h06 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h07 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h08 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h09 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h0a :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h0b :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h0c :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h0d :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h0e :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h0f :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h10 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h11 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h12 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h13 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h14 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h15 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h16 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h17 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h18 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h19 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h1a :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h1b :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h1c :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h1d :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h1e :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h1f :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h20 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h21 :
		RG_quantized_block_rl_14_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h22 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h23 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h24 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h25 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h26 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h27 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h28 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h29 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h2a :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h2b :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h2c :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h2d :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h2e :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h2f :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h30 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h31 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h32 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h33 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h34 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h35 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h36 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h37 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h38 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h39 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h3a :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h3b :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h3c :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h3d :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h3e :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h3f :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h40 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h41 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h42 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h43 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h44 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h45 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h46 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h47 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h48 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h49 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h4a :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h4b :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h4c :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h4d :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h4e :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h4f :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h50 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h51 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h52 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h53 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h54 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h55 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h56 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h57 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h58 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h59 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h5a :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h5b :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h5c :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h5d :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h5e :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h5f :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h60 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h61 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h62 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h63 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h64 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h65 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h66 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h67 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h68 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h69 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h6a :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h6b :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h6c :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h6d :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h6e :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h6f :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h70 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h71 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h72 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h73 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h74 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h75 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h76 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h77 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h78 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h79 :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h7a :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h7b :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h7c :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h7d :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h7e :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	7'h7f :
		RG_quantized_block_rl_14_t1 = rl_a33_t8 ;
	default :
		RG_quantized_block_rl_14_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_14_t1 or U_318 or TR_232 or U_317 or RG_rl_35 or 
	ST1_07d or RG_rl_33 or U_88 or jpeg_in_a14 or U_01 or RG_quantized_block_rl_16 or 
	ST1_01d )
	RG_quantized_block_rl_14_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_16 )
		| ( { 9{ U_01 } } & jpeg_in_a14 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_33 )
		| ( { 9{ ST1_07d } } & RG_rl_35 )
		| ( { 9{ U_317 } } & TR_232 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_14_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_14_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_14_en )
		RG_quantized_block_rl_14 <= RG_quantized_block_rl_14_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a35_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h01 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h02 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h03 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h04 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h05 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h06 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h07 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h08 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h09 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h0a :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h0b :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h0c :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h0d :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h0e :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h0f :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h10 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h11 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h12 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h13 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h14 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h15 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h16 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h17 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h18 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h19 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h1a :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h1b :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h1c :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h1d :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h1e :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h1f :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h20 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h21 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h22 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h23 :
		RG_quantized_block_rl_15_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h24 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h25 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h26 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h27 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h28 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h29 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h2a :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h2b :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h2c :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h2d :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h2e :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h2f :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h30 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h31 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h32 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h33 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h34 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h35 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h36 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h37 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h38 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h39 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h3a :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h3b :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h3c :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h3d :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h3e :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h3f :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h40 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h41 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h42 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h43 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h44 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h45 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h46 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h47 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h48 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h49 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h4a :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h4b :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h4c :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h4d :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h4e :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h4f :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h50 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h51 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h52 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h53 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h54 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h55 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h56 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h57 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h58 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h59 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h5a :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h5b :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h5c :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h5d :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h5e :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h5f :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h60 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h61 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h62 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h63 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h64 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h65 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h66 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h67 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h68 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h69 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h6a :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h6b :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h6c :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h6d :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h6e :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h6f :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h70 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h71 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h72 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h73 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h74 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h75 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h76 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h77 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h78 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h79 :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h7a :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h7b :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h7c :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h7d :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h7e :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	7'h7f :
		RG_quantized_block_rl_15_t1 = rl_a35_t8 ;
	default :
		RG_quantized_block_rl_15_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_15_t1 or U_318 or TR_230 or U_317 or RG_rl_37 or 
	ST1_07d or RG_rl_35 or U_88 or jpeg_in_a15 or U_01 or RG_quantized_block_rl_17 or 
	ST1_01d )
	RG_quantized_block_rl_15_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_17 )
		| ( { 9{ U_01 } } & jpeg_in_a15 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_35 )
		| ( { 9{ ST1_07d } } & RG_rl_37 )
		| ( { 9{ U_317 } } & TR_230 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_15_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_15_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_15_en )
		RG_quantized_block_rl_15 <= RG_quantized_block_rl_15_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a37_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h01 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h02 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h03 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h04 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h05 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h06 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h07 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h08 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h09 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h0a :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h0b :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h0c :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h0d :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h0e :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h0f :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h10 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h11 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h12 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h13 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h14 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h15 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h16 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h17 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h18 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h19 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h1a :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h1b :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h1c :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h1d :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h1e :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h1f :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h20 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h21 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h22 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h23 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h24 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h25 :
		RG_quantized_block_rl_16_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h26 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h27 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h28 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h29 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h2a :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h2b :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h2c :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h2d :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h2e :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h2f :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h30 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h31 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h32 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h33 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h34 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h35 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h36 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h37 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h38 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h39 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h3a :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h3b :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h3c :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h3d :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h3e :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h3f :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h40 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h41 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h42 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h43 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h44 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h45 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h46 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h47 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h48 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h49 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h4a :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h4b :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h4c :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h4d :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h4e :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h4f :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h50 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h51 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h52 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h53 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h54 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h55 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h56 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h57 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h58 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h59 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h5a :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h5b :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h5c :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h5d :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h5e :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h5f :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h60 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h61 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h62 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h63 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h64 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h65 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h66 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h67 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h68 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h69 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h6a :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h6b :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h6c :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h6d :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h6e :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h6f :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h70 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h71 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h72 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h73 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h74 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h75 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h76 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h77 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h78 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h79 :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h7a :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h7b :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h7c :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h7d :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h7e :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	7'h7f :
		RG_quantized_block_rl_16_t1 = rl_a37_t8 ;
	default :
		RG_quantized_block_rl_16_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_16_t1 or U_318 or TR_228 or U_317 or RG_rl_39 or 
	ST1_07d or RG_rl_37 or U_88 or jpeg_in_a16 or U_01 or RG_quantized_block_rl_18 or 
	ST1_01d )
	RG_quantized_block_rl_16_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_18 )
		| ( { 9{ U_01 } } & jpeg_in_a16 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_37 )
		| ( { 9{ ST1_07d } } & RG_rl_39 )
		| ( { 9{ U_317 } } & TR_228 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_16_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_16_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_16_en )
		RG_quantized_block_rl_16 <= RG_quantized_block_rl_16_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a39_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h01 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h02 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h03 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h04 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h05 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h06 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h07 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h08 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h09 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h0a :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h0b :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h0c :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h0d :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h0e :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h0f :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h10 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h11 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h12 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h13 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h14 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h15 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h16 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h17 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h18 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h19 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h1a :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h1b :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h1c :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h1d :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h1e :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h1f :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h20 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h21 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h22 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h23 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h24 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h25 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h26 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h27 :
		RG_quantized_block_rl_17_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h28 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h29 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h2a :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h2b :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h2c :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h2d :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h2e :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h2f :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h30 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h31 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h32 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h33 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h34 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h35 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h36 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h37 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h38 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h39 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h3a :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h3b :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h3c :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h3d :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h3e :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h3f :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h40 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h41 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h42 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h43 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h44 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h45 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h46 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h47 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h48 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h49 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h4a :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h4b :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h4c :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h4d :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h4e :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h4f :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h50 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h51 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h52 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h53 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h54 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h55 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h56 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h57 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h58 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h59 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h5a :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h5b :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h5c :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h5d :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h5e :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h5f :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h60 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h61 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h62 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h63 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h64 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h65 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h66 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h67 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h68 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h69 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h6a :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h6b :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h6c :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h6d :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h6e :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h6f :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h70 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h71 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h72 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h73 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h74 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h75 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h76 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h77 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h78 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h79 :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h7a :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h7b :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h7c :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h7d :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h7e :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	7'h7f :
		RG_quantized_block_rl_17_t1 = rl_a39_t8 ;
	default :
		RG_quantized_block_rl_17_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_17_t1 or U_318 or TR_226 or U_317 or RG_rl_41 or 
	ST1_07d or RG_rl_39 or U_88 or jpeg_in_a17 or U_01 or RG_quantized_block_rl_19 or 
	ST1_01d )
	RG_quantized_block_rl_17_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_19 )
		| ( { 9{ U_01 } } & jpeg_in_a17 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_39 )
		| ( { 9{ ST1_07d } } & RG_rl_41 )
		| ( { 9{ U_317 } } & TR_226 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_17_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_17_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_17_en )
		RG_quantized_block_rl_17 <= RG_quantized_block_rl_17_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a41_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h01 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h02 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h03 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h04 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h05 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h06 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h07 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h08 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h09 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h0a :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h0b :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h0c :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h0d :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h0e :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h0f :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h10 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h11 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h12 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h13 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h14 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h15 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h16 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h17 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h18 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h19 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h1a :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h1b :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h1c :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h1d :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h1e :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h1f :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h20 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h21 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h22 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h23 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h24 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h25 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h26 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h27 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h28 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h29 :
		RG_quantized_block_rl_18_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h2a :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h2b :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h2c :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h2d :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h2e :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h2f :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h30 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h31 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h32 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h33 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h34 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h35 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h36 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h37 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h38 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h39 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h3a :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h3b :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h3c :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h3d :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h3e :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h3f :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h40 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h41 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h42 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h43 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h44 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h45 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h46 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h47 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h48 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h49 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h4a :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h4b :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h4c :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h4d :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h4e :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h4f :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h50 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h51 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h52 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h53 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h54 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h55 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h56 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h57 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h58 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h59 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h5a :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h5b :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h5c :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h5d :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h5e :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h5f :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h60 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h61 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h62 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h63 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h64 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h65 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h66 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h67 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h68 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h69 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h6a :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h6b :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h6c :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h6d :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h6e :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h6f :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h70 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h71 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h72 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h73 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h74 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h75 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h76 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h77 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h78 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h79 :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h7a :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h7b :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h7c :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h7d :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h7e :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	7'h7f :
		RG_quantized_block_rl_18_t1 = rl_a41_t8 ;
	default :
		RG_quantized_block_rl_18_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_18_t1 or U_318 or TR_224 or U_317 or RG_rl_43 or 
	ST1_07d or RG_rl_41 or U_88 or jpeg_in_a18 or U_01 or RG_quantized_block_rl_20 or 
	ST1_01d )
	RG_quantized_block_rl_18_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_20 )
		| ( { 9{ U_01 } } & jpeg_in_a18 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_41 )
		| ( { 9{ ST1_07d } } & RG_rl_43 )
		| ( { 9{ U_317 } } & TR_224 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_18_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_18_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_18_en )
		RG_quantized_block_rl_18 <= RG_quantized_block_rl_18_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a43_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h01 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h02 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h03 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h04 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h05 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h06 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h07 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h08 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h09 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h0a :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h0b :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h0c :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h0d :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h0e :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h0f :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h10 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h11 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h12 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h13 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h14 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h15 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h16 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h17 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h18 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h19 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h1a :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h1b :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h1c :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h1d :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h1e :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h1f :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h20 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h21 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h22 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h23 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h24 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h25 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h26 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h27 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h28 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h29 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h2a :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h2b :
		RG_quantized_block_rl_19_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h2c :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h2d :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h2e :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h2f :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h30 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h31 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h32 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h33 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h34 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h35 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h36 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h37 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h38 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h39 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h3a :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h3b :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h3c :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h3d :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h3e :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h3f :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h40 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h41 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h42 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h43 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h44 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h45 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h46 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h47 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h48 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h49 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h4a :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h4b :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h4c :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h4d :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h4e :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h4f :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h50 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h51 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h52 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h53 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h54 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h55 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h56 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h57 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h58 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h59 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h5a :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h5b :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h5c :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h5d :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h5e :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h5f :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h60 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h61 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h62 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h63 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h64 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h65 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h66 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h67 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h68 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h69 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h6a :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h6b :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h6c :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h6d :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h6e :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h6f :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h70 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h71 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h72 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h73 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h74 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h75 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h76 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h77 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h78 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h79 :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h7a :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h7b :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h7c :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h7d :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h7e :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	7'h7f :
		RG_quantized_block_rl_19_t1 = rl_a43_t8 ;
	default :
		RG_quantized_block_rl_19_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_19_t1 or U_318 or TR_222 or U_317 or RG_rl_45 or 
	ST1_07d or RG_rl_43 or U_88 or jpeg_in_a19 or U_01 or RG_quantized_block_rl_21 or 
	ST1_01d )
	RG_quantized_block_rl_19_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_21 )
		| ( { 9{ U_01 } } & jpeg_in_a19 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_43 )
		| ( { 9{ ST1_07d } } & RG_rl_45 )
		| ( { 9{ U_317 } } & TR_222 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_19_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_19_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_19_en )
		RG_quantized_block_rl_19 <= RG_quantized_block_rl_19_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a45_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h01 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h02 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h03 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h04 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h05 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h06 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h07 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h08 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h09 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h0a :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h0b :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h0c :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h0d :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h0e :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h0f :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h10 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h11 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h12 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h13 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h14 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h15 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h16 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h17 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h18 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h19 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h1a :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h1b :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h1c :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h1d :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h1e :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h1f :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h20 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h21 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h22 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h23 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h24 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h25 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h26 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h27 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h28 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h29 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h2a :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h2b :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h2c :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h2d :
		RG_quantized_block_rl_20_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h2e :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h2f :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h30 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h31 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h32 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h33 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h34 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h35 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h36 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h37 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h38 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h39 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h3a :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h3b :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h3c :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h3d :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h3e :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h3f :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h40 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h41 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h42 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h43 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h44 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h45 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h46 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h47 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h48 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h49 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h4a :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h4b :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h4c :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h4d :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h4e :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h4f :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h50 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h51 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h52 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h53 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h54 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h55 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h56 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h57 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h58 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h59 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h5a :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h5b :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h5c :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h5d :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h5e :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h5f :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h60 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h61 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h62 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h63 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h64 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h65 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h66 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h67 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h68 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h69 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h6a :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h6b :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h6c :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h6d :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h6e :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h6f :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h70 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h71 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h72 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h73 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h74 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h75 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h76 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h77 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h78 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h79 :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h7a :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h7b :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h7c :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h7d :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h7e :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	7'h7f :
		RG_quantized_block_rl_20_t1 = rl_a45_t8 ;
	default :
		RG_quantized_block_rl_20_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_20_t1 or U_318 or TR_220 or U_317 or RG_rl_47 or 
	ST1_07d or RG_rl_45 or U_88 or jpeg_in_a20 or U_01 or RG_quantized_block_rl_22 or 
	ST1_01d )
	RG_quantized_block_rl_20_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_22 )
		| ( { 9{ U_01 } } & jpeg_in_a20 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_45 )
		| ( { 9{ ST1_07d } } & RG_rl_47 )
		| ( { 9{ U_317 } } & TR_220 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_20_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_20_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_20_en )
		RG_quantized_block_rl_20 <= RG_quantized_block_rl_20_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a47_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h01 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h02 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h03 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h04 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h05 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h06 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h07 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h08 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h09 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h0a :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h0b :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h0c :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h0d :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h0e :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h0f :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h10 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h11 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h12 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h13 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h14 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h15 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h16 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h17 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h18 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h19 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h1a :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h1b :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h1c :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h1d :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h1e :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h1f :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h20 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h21 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h22 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h23 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h24 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h25 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h26 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h27 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h28 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h29 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h2a :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h2b :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h2c :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h2d :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h2e :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h2f :
		RG_quantized_block_rl_21_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h30 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h31 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h32 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h33 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h34 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h35 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h36 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h37 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h38 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h39 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h3a :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h3b :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h3c :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h3d :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h3e :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h3f :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h40 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h41 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h42 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h43 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h44 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h45 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h46 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h47 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h48 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h49 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h4a :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h4b :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h4c :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h4d :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h4e :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h4f :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h50 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h51 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h52 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h53 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h54 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h55 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h56 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h57 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h58 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h59 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h5a :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h5b :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h5c :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h5d :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h5e :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h5f :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h60 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h61 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h62 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h63 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h64 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h65 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h66 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h67 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h68 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h69 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h6a :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h6b :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h6c :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h6d :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h6e :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h6f :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h70 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h71 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h72 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h73 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h74 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h75 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h76 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h77 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h78 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h79 :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h7a :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h7b :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h7c :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h7d :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h7e :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	7'h7f :
		RG_quantized_block_rl_21_t1 = rl_a47_t8 ;
	default :
		RG_quantized_block_rl_21_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_21_t1 or U_318 or TR_218 or U_317 or RG_rl_49 or 
	ST1_07d or RG_rl_47 or U_88 or jpeg_in_a21 or U_01 or RG_quantized_block_rl_23 or 
	ST1_01d )
	RG_quantized_block_rl_21_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_23 )
		| ( { 9{ U_01 } } & jpeg_in_a21 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_47 )
		| ( { 9{ ST1_07d } } & RG_rl_49 )
		| ( { 9{ U_317 } } & TR_218 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_21_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_21_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_21_en )
		RG_quantized_block_rl_21 <= RG_quantized_block_rl_21_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a49_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h01 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h02 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h03 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h04 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h05 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h06 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h07 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h08 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h09 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h0a :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h0b :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h0c :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h0d :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h0e :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h0f :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h10 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h11 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h12 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h13 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h14 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h15 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h16 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h17 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h18 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h19 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h1a :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h1b :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h1c :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h1d :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h1e :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h1f :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h20 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h21 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h22 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h23 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h24 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h25 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h26 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h27 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h28 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h29 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h2a :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h2b :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h2c :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h2d :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h2e :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h2f :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h30 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h31 :
		RG_quantized_block_rl_22_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h32 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h33 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h34 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h35 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h36 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h37 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h38 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h39 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h3a :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h3b :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h3c :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h3d :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h3e :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h3f :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h40 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h41 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h42 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h43 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h44 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h45 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h46 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h47 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h48 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h49 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h4a :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h4b :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h4c :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h4d :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h4e :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h4f :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h50 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h51 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h52 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h53 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h54 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h55 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h56 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h57 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h58 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h59 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h5a :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h5b :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h5c :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h5d :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h5e :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h5f :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h60 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h61 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h62 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h63 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h64 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h65 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h66 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h67 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h68 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h69 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h6a :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h6b :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h6c :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h6d :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h6e :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h6f :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h70 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h71 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h72 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h73 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h74 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h75 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h76 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h77 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h78 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h79 :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h7a :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h7b :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h7c :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h7d :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h7e :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	7'h7f :
		RG_quantized_block_rl_22_t1 = rl_a49_t8 ;
	default :
		RG_quantized_block_rl_22_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_22_t1 or U_318 or TR_216 or U_317 or RG_rl_51 or 
	ST1_07d or RG_rl_49 or U_88 or jpeg_in_a22 or U_01 or RG_quantized_block_rl_24 or 
	ST1_01d )
	RG_quantized_block_rl_22_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_24 )
		| ( { 9{ U_01 } } & jpeg_in_a22 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_49 )
		| ( { 9{ ST1_07d } } & RG_rl_51 )
		| ( { 9{ U_317 } } & TR_216 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_22_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_22_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_22_en )
		RG_quantized_block_rl_22 <= RG_quantized_block_rl_22_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a51_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h01 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h02 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h03 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h04 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h05 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h06 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h07 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h08 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h09 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h0a :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h0b :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h0c :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h0d :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h0e :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h0f :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h10 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h11 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h12 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h13 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h14 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h15 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h16 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h17 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h18 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h19 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h1a :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h1b :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h1c :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h1d :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h1e :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h1f :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h20 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h21 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h22 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h23 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h24 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h25 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h26 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h27 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h28 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h29 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h2a :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h2b :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h2c :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h2d :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h2e :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h2f :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h30 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h31 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h32 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h33 :
		RG_quantized_block_rl_23_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h34 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h35 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h36 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h37 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h38 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h39 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h3a :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h3b :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h3c :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h3d :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h3e :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h3f :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h40 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h41 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h42 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h43 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h44 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h45 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h46 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h47 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h48 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h49 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h4a :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h4b :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h4c :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h4d :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h4e :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h4f :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h50 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h51 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h52 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h53 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h54 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h55 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h56 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h57 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h58 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h59 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h5a :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h5b :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h5c :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h5d :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h5e :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h5f :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h60 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h61 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h62 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h63 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h64 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h65 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h66 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h67 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h68 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h69 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h6a :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h6b :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h6c :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h6d :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h6e :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h6f :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h70 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h71 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h72 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h73 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h74 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h75 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h76 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h77 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h78 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h79 :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h7a :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h7b :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h7c :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h7d :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h7e :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	7'h7f :
		RG_quantized_block_rl_23_t1 = rl_a51_t8 ;
	default :
		RG_quantized_block_rl_23_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_23_t1 or U_318 or TR_214 or U_317 or RG_rl_53 or 
	ST1_07d or RG_rl_51 or U_88 or jpeg_in_a23 or U_01 or RG_quantized_block_rl_25 or 
	ST1_01d )
	RG_quantized_block_rl_23_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_25 )
		| ( { 9{ U_01 } } & jpeg_in_a23 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_51 )
		| ( { 9{ ST1_07d } } & RG_rl_53 )
		| ( { 9{ U_317 } } & TR_214 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_23_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_23_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_23_en )
		RG_quantized_block_rl_23 <= RG_quantized_block_rl_23_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a53_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h01 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h02 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h03 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h04 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h05 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h06 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h07 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h08 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h09 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h0a :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h0b :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h0c :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h0d :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h0e :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h0f :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h10 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h11 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h12 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h13 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h14 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h15 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h16 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h17 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h18 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h19 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h1a :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h1b :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h1c :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h1d :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h1e :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h1f :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h20 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h21 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h22 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h23 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h24 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h25 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h26 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h27 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h28 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h29 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h2a :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h2b :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h2c :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h2d :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h2e :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h2f :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h30 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h31 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h32 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h33 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h34 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h35 :
		RG_quantized_block_rl_24_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h36 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h37 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h38 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h39 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h3a :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h3b :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h3c :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h3d :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h3e :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h3f :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h40 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h41 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h42 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h43 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h44 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h45 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h46 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h47 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h48 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h49 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h4a :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h4b :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h4c :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h4d :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h4e :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h4f :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h50 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h51 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h52 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h53 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h54 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h55 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h56 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h57 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h58 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h59 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h5a :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h5b :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h5c :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h5d :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h5e :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h5f :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h60 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h61 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h62 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h63 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h64 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h65 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h66 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h67 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h68 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h69 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h6a :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h6b :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h6c :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h6d :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h6e :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h6f :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h70 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h71 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h72 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h73 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h74 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h75 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h76 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h77 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h78 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h79 :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h7a :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h7b :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h7c :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h7d :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h7e :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	7'h7f :
		RG_quantized_block_rl_24_t1 = rl_a53_t8 ;
	default :
		RG_quantized_block_rl_24_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_24_t1 or U_318 or TR_212 or U_317 or RG_rl_55 or 
	ST1_07d or RG_rl_53 or U_88 or jpeg_in_a24 or U_01 or RG_quantized_block_rl_26 or 
	ST1_01d )
	RG_quantized_block_rl_24_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_26 )
		| ( { 9{ U_01 } } & jpeg_in_a24 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_53 )
		| ( { 9{ ST1_07d } } & RG_rl_55 )
		| ( { 9{ U_317 } } & TR_212 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_24_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_24_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_24_en )
		RG_quantized_block_rl_24 <= RG_quantized_block_rl_24_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a55_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h01 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h02 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h03 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h04 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h05 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h06 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h07 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h08 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h09 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h0a :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h0b :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h0c :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h0d :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h0e :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h0f :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h10 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h11 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h12 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h13 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h14 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h15 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h16 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h17 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h18 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h19 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h1a :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h1b :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h1c :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h1d :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h1e :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h1f :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h20 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h21 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h22 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h23 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h24 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h25 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h26 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h27 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h28 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h29 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h2a :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h2b :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h2c :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h2d :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h2e :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h2f :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h30 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h31 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h32 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h33 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h34 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h35 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h36 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h37 :
		RG_quantized_block_rl_25_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h38 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h39 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h3a :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h3b :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h3c :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h3d :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h3e :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h3f :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h40 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h41 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h42 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h43 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h44 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h45 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h46 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h47 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h48 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h49 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h4a :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h4b :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h4c :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h4d :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h4e :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h4f :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h50 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h51 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h52 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h53 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h54 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h55 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h56 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h57 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h58 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h59 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h5a :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h5b :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h5c :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h5d :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h5e :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h5f :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h60 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h61 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h62 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h63 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h64 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h65 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h66 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h67 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h68 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h69 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h6a :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h6b :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h6c :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h6d :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h6e :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h6f :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h70 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h71 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h72 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h73 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h74 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h75 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h76 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h77 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h78 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h79 :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h7a :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h7b :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h7c :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h7d :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h7e :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	7'h7f :
		RG_quantized_block_rl_25_t1 = rl_a55_t8 ;
	default :
		RG_quantized_block_rl_25_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_25_t1 or U_318 or TR_210 or U_317 or RG_rl_57 or 
	ST1_07d or RG_rl_55 or U_88 or jpeg_in_a25 or U_01 or RG_quantized_block_rl_27 or 
	ST1_01d )
	RG_quantized_block_rl_25_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_27 )
		| ( { 9{ U_01 } } & jpeg_in_a25 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_55 )
		| ( { 9{ ST1_07d } } & RG_rl_57 )
		| ( { 9{ U_317 } } & TR_210 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_25_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_25_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_25_en )
		RG_quantized_block_rl_25 <= RG_quantized_block_rl_25_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a57_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h01 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h02 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h03 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h04 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h05 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h06 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h07 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h08 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h09 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h0a :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h0b :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h0c :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h0d :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h0e :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h0f :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h10 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h11 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h12 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h13 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h14 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h15 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h16 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h17 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h18 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h19 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h1a :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h1b :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h1c :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h1d :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h1e :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h1f :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h20 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h21 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h22 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h23 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h24 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h25 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h26 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h27 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h28 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h29 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h2a :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h2b :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h2c :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h2d :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h2e :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h2f :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h30 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h31 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h32 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h33 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h34 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h35 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h36 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h37 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h38 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h39 :
		RG_quantized_block_rl_26_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h3a :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h3b :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h3c :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h3d :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h3e :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h3f :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h40 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h41 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h42 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h43 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h44 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h45 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h46 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h47 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h48 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h49 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h4a :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h4b :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h4c :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h4d :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h4e :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h4f :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h50 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h51 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h52 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h53 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h54 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h55 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h56 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h57 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h58 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h59 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h5a :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h5b :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h5c :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h5d :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h5e :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h5f :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h60 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h61 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h62 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h63 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h64 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h65 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h66 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h67 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h68 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h69 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h6a :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h6b :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h6c :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h6d :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h6e :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h6f :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h70 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h71 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h72 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h73 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h74 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h75 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h76 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h77 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h78 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h79 :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h7a :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h7b :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h7c :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h7d :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h7e :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	7'h7f :
		RG_quantized_block_rl_26_t1 = rl_a57_t8 ;
	default :
		RG_quantized_block_rl_26_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_26_t1 or U_318 or TR_208 or U_317 or RG_rl_59 or 
	ST1_07d or RG_rl_57 or U_88 or jpeg_in_a26 or U_01 or RG_quantized_block_rl_28 or 
	ST1_01d )
	RG_quantized_block_rl_26_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_28 )
		| ( { 9{ U_01 } } & jpeg_in_a26 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_57 )
		| ( { 9{ ST1_07d } } & RG_rl_59 )
		| ( { 9{ U_317 } } & TR_208 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_26_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_26_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_26_en )
		RG_quantized_block_rl_26 <= RG_quantized_block_rl_26_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a59_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h01 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h02 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h03 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h04 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h05 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h06 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h07 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h08 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h09 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h0a :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h0b :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h0c :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h0d :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h0e :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h0f :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h10 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h11 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h12 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h13 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h14 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h15 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h16 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h17 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h18 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h19 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h1a :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h1b :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h1c :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h1d :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h1e :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h1f :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h20 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h21 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h22 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h23 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h24 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h25 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h26 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h27 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h28 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h29 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h2a :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h2b :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h2c :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h2d :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h2e :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h2f :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h30 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h31 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h32 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h33 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h34 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h35 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h36 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h37 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h38 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h39 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h3a :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h3b :
		RG_quantized_block_rl_27_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h3c :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h3d :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h3e :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h3f :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h40 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h41 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h42 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h43 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h44 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h45 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h46 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h47 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h48 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h49 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h4a :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h4b :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h4c :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h4d :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h4e :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h4f :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h50 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h51 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h52 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h53 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h54 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h55 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h56 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h57 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h58 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h59 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h5a :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h5b :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h5c :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h5d :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h5e :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h5f :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h60 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h61 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h62 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h63 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h64 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h65 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h66 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h67 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h68 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h69 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h6a :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h6b :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h6c :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h6d :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h6e :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h6f :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h70 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h71 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h72 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h73 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h74 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h75 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h76 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h77 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h78 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h79 :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h7a :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h7b :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h7c :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h7d :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h7e :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	7'h7f :
		RG_quantized_block_rl_27_t1 = rl_a59_t8 ;
	default :
		RG_quantized_block_rl_27_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_27_t1 or U_318 or TR_206 or U_317 or RG_rl_61 or 
	ST1_07d or RG_rl_59 or U_88 or jpeg_in_a27 or U_01 or RG_quantized_block_rl_29 or 
	ST1_01d )
	RG_quantized_block_rl_27_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_29 )
		| ( { 9{ U_01 } } & jpeg_in_a27 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_59 )
		| ( { 9{ ST1_07d } } & RG_rl_61 )
		| ( { 9{ U_317 } } & TR_206 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_27_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_27_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_27_en )
		RG_quantized_block_rl_27 <= RG_quantized_block_rl_27_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a61_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h01 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h02 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h03 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h04 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h05 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h06 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h07 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h08 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h09 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h0a :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h0b :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h0c :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h0d :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h0e :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h0f :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h10 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h11 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h12 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h13 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h14 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h15 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h16 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h17 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h18 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h19 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h1a :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h1b :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h1c :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h1d :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h1e :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h1f :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h20 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h21 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h22 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h23 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h24 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h25 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h26 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h27 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h28 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h29 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h2a :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h2b :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h2c :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h2d :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h2e :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h2f :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h30 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h31 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h32 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h33 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h34 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h35 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h36 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h37 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h38 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h39 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h3a :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h3b :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h3c :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h3d :
		RG_quantized_block_rl_28_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h3e :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h3f :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h40 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h41 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h42 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h43 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h44 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h45 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h46 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h47 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h48 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h49 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h4a :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h4b :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h4c :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h4d :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h4e :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h4f :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h50 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h51 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h52 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h53 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h54 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h55 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h56 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h57 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h58 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h59 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h5a :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h5b :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h5c :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h5d :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h5e :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h5f :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h60 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h61 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h62 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h63 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h64 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h65 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h66 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h67 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h68 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h69 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h6a :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h6b :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h6c :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h6d :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h6e :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h6f :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h70 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h71 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h72 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h73 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h74 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h75 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h76 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h77 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h78 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h79 :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h7a :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h7b :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h7c :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h7d :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h7e :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	7'h7f :
		RG_quantized_block_rl_28_t1 = rl_a61_t8 ;
	default :
		RG_quantized_block_rl_28_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_28_t1 or U_318 or TR_204 or U_317 or RG_rl_63 or 
	ST1_07d or RG_rl_61 or U_88 or jpeg_in_a28 or U_01 or RG_quantized_block_rl_30 or 
	ST1_01d )
	RG_quantized_block_rl_28_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_30 )
		| ( { 9{ U_01 } } & jpeg_in_a28 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_61 )
		| ( { 9{ ST1_07d } } & RG_rl_63 )
		| ( { 9{ U_317 } } & TR_204 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_28_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_28_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_28_en )
		RG_quantized_block_rl_28 <= RG_quantized_block_rl_28_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a63_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h01 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h02 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h03 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h04 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h05 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h06 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h07 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h08 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h09 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h0a :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h0b :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h0c :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h0d :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h0e :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h0f :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h10 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h11 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h12 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h13 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h14 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h15 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h16 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h17 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h18 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h19 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h1a :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h1b :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h1c :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h1d :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h1e :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h1f :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h20 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h21 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h22 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h23 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h24 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h25 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h26 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h27 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h28 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h29 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h2a :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h2b :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h2c :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h2d :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h2e :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h2f :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h30 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h31 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h32 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h33 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h34 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h35 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h36 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h37 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h38 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h39 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h3a :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h3b :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h3c :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h3d :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h3e :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h3f :
		RG_quantized_block_rl_29_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h40 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h41 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h42 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h43 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h44 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h45 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h46 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h47 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h48 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h49 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h4a :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h4b :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h4c :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h4d :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h4e :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h4f :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h50 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h51 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h52 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h53 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h54 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h55 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h56 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h57 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h58 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h59 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h5a :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h5b :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h5c :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h5d :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h5e :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h5f :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h60 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h61 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h62 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h63 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h64 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h65 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h66 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h67 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h68 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h69 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h6a :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h6b :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h6c :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h6d :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h6e :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h6f :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h70 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h71 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h72 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h73 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h74 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h75 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h76 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h77 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h78 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h79 :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h7a :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h7b :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h7c :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h7d :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h7e :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	7'h7f :
		RG_quantized_block_rl_29_t1 = rl_a63_t8 ;
	default :
		RG_quantized_block_rl_29_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_29_t1 or U_318 or TR_202 or U_317 or RG_rl_65 or 
	ST1_07d or RG_rl_63 or U_88 or jpeg_in_a29 or U_01 or RG_quantized_block_rl_31 or 
	ST1_01d )
	RG_quantized_block_rl_29_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_31 )
		| ( { 9{ U_01 } } & jpeg_in_a29 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_63 )
		| ( { 9{ ST1_07d } } & RG_rl_65 )
		| ( { 9{ U_317 } } & TR_202 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_29_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_29_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_29_en )
		RG_quantized_block_rl_29 <= RG_quantized_block_rl_29_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a65_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h01 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h02 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h03 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h04 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h05 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h06 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h07 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h08 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h09 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h0a :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h0b :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h0c :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h0d :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h0e :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h0f :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h10 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h11 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h12 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h13 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h14 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h15 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h16 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h17 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h18 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h19 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h1a :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h1b :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h1c :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h1d :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h1e :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h1f :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h20 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h21 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h22 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h23 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h24 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h25 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h26 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h27 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h28 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h29 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h2a :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h2b :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h2c :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h2d :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h2e :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h2f :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h30 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h31 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h32 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h33 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h34 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h35 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h36 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h37 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h38 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h39 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h3a :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h3b :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h3c :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h3d :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h3e :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h3f :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h40 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h41 :
		RG_quantized_block_rl_30_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h42 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h43 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h44 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h45 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h46 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h47 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h48 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h49 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h4a :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h4b :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h4c :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h4d :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h4e :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h4f :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h50 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h51 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h52 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h53 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h54 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h55 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h56 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h57 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h58 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h59 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h5a :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h5b :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h5c :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h5d :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h5e :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h5f :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h60 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h61 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h62 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h63 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h64 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h65 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h66 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h67 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h68 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h69 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h6a :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h6b :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h6c :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h6d :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h6e :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h6f :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h70 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h71 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h72 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h73 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h74 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h75 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h76 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h77 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h78 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h79 :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h7a :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h7b :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h7c :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h7d :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h7e :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	7'h7f :
		RG_quantized_block_rl_30_t1 = rl_a65_t8 ;
	default :
		RG_quantized_block_rl_30_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_30_t1 or U_318 or TR_200 or U_317 or RG_rl_67 or 
	ST1_07d or RG_rl_65 or U_88 or jpeg_in_a30 or U_01 or RG_quantized_block_rl_32 or 
	ST1_01d )
	RG_quantized_block_rl_30_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_32 )
		| ( { 9{ U_01 } } & jpeg_in_a30 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_65 )
		| ( { 9{ ST1_07d } } & RG_rl_67 )
		| ( { 9{ U_317 } } & TR_200 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_30_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_30_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_30_en )
		RG_quantized_block_rl_30 <= RG_quantized_block_rl_30_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a67_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h01 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h02 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h03 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h04 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h05 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h06 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h07 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h08 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h09 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h0a :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h0b :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h0c :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h0d :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h0e :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h0f :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h10 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h11 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h12 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h13 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h14 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h15 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h16 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h17 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h18 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h19 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h1a :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h1b :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h1c :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h1d :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h1e :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h1f :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h20 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h21 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h22 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h23 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h24 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h25 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h26 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h27 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h28 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h29 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h2a :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h2b :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h2c :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h2d :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h2e :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h2f :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h30 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h31 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h32 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h33 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h34 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h35 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h36 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h37 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h38 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h39 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h3a :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h3b :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h3c :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h3d :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h3e :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h3f :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h40 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h41 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h42 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h43 :
		RG_quantized_block_rl_31_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h44 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h45 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h46 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h47 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h48 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h49 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h4a :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h4b :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h4c :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h4d :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h4e :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h4f :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h50 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h51 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h52 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h53 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h54 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h55 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h56 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h57 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h58 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h59 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h5a :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h5b :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h5c :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h5d :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h5e :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h5f :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h60 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h61 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h62 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h63 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h64 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h65 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h66 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h67 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h68 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h69 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h6a :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h6b :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h6c :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h6d :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h6e :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h6f :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h70 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h71 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h72 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h73 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h74 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h75 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h76 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h77 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h78 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h79 :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h7a :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h7b :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h7c :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h7d :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h7e :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	7'h7f :
		RG_quantized_block_rl_31_t1 = rl_a67_t8 ;
	default :
		RG_quantized_block_rl_31_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_31_t1 or U_318 or TR_198 or U_317 or RG_rl_69 or 
	ST1_07d or RG_rl_67 or U_88 or jpeg_in_a31 or U_01 or RG_quantized_block_rl_33 or 
	ST1_01d )
	RG_quantized_block_rl_31_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_33 )
		| ( { 9{ U_01 } } & jpeg_in_a31 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_67 )
		| ( { 9{ ST1_07d } } & RG_rl_69 )
		| ( { 9{ U_317 } } & TR_198 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_31_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_31_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_31_en )
		RG_quantized_block_rl_31 <= RG_quantized_block_rl_31_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a69_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h01 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h02 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h03 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h04 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h05 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h06 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h07 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h08 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h09 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h0a :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h0b :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h0c :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h0d :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h0e :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h0f :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h10 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h11 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h12 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h13 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h14 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h15 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h16 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h17 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h18 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h19 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h1a :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h1b :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h1c :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h1d :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h1e :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h1f :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h20 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h21 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h22 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h23 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h24 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h25 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h26 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h27 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h28 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h29 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h2a :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h2b :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h2c :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h2d :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h2e :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h2f :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h30 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h31 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h32 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h33 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h34 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h35 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h36 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h37 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h38 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h39 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h3a :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h3b :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h3c :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h3d :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h3e :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h3f :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h40 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h41 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h42 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h43 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h44 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h45 :
		RG_quantized_block_rl_32_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h46 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h47 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h48 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h49 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h4a :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h4b :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h4c :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h4d :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h4e :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h4f :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h50 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h51 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h52 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h53 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h54 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h55 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h56 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h57 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h58 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h59 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h5a :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h5b :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h5c :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h5d :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h5e :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h5f :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h60 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h61 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h62 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h63 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h64 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h65 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h66 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h67 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h68 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h69 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h6a :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h6b :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h6c :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h6d :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h6e :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h6f :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h70 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h71 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h72 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h73 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h74 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h75 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h76 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h77 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h78 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h79 :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h7a :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h7b :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h7c :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h7d :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h7e :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	7'h7f :
		RG_quantized_block_rl_32_t1 = rl_a69_t8 ;
	default :
		RG_quantized_block_rl_32_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_32_t1 or U_318 or TR_196 or U_317 or RG_rl_71 or 
	ST1_07d or RG_rl_69 or U_88 or jpeg_in_a32 or U_01 or RG_quantized_block_rl_34 or 
	ST1_01d )
	RG_quantized_block_rl_32_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_34 )
		| ( { 9{ U_01 } } & jpeg_in_a32 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_69 )
		| ( { 9{ ST1_07d } } & RG_rl_71 )
		| ( { 9{ U_317 } } & TR_196 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_32_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_32_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_32_en )
		RG_quantized_block_rl_32 <= RG_quantized_block_rl_32_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a71_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h01 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h02 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h03 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h04 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h05 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h06 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h07 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h08 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h09 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h0a :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h0b :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h0c :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h0d :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h0e :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h0f :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h10 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h11 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h12 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h13 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h14 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h15 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h16 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h17 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h18 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h19 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h1a :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h1b :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h1c :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h1d :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h1e :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h1f :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h20 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h21 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h22 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h23 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h24 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h25 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h26 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h27 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h28 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h29 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h2a :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h2b :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h2c :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h2d :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h2e :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h2f :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h30 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h31 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h32 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h33 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h34 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h35 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h36 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h37 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h38 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h39 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h3a :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h3b :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h3c :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h3d :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h3e :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h3f :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h40 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h41 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h42 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h43 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h44 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h45 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h46 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h47 :
		RG_quantized_block_rl_33_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h48 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h49 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h4a :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h4b :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h4c :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h4d :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h4e :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h4f :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h50 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h51 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h52 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h53 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h54 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h55 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h56 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h57 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h58 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h59 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h5a :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h5b :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h5c :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h5d :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h5e :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h5f :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h60 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h61 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h62 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h63 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h64 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h65 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h66 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h67 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h68 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h69 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h6a :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h6b :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h6c :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h6d :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h6e :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h6f :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h70 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h71 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h72 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h73 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h74 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h75 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h76 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h77 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h78 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h79 :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h7a :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h7b :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h7c :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h7d :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h7e :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	7'h7f :
		RG_quantized_block_rl_33_t1 = rl_a71_t8 ;
	default :
		RG_quantized_block_rl_33_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_33_t1 or U_318 or TR_194 or U_317 or RG_rl_73 or 
	ST1_07d or RG_rl_71 or U_88 or jpeg_in_a33 or U_01 or RG_quantized_block_rl_35 or 
	ST1_01d )
	RG_quantized_block_rl_33_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_35 )
		| ( { 9{ U_01 } } & jpeg_in_a33 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_71 )
		| ( { 9{ ST1_07d } } & RG_rl_73 )
		| ( { 9{ U_317 } } & TR_194 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_33_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_33_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_33_en )
		RG_quantized_block_rl_33 <= RG_quantized_block_rl_33_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a73_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h01 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h02 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h03 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h04 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h05 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h06 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h07 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h08 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h09 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h0a :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h0b :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h0c :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h0d :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h0e :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h0f :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h10 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h11 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h12 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h13 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h14 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h15 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h16 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h17 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h18 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h19 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h1a :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h1b :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h1c :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h1d :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h1e :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h1f :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h20 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h21 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h22 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h23 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h24 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h25 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h26 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h27 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h28 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h29 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h2a :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h2b :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h2c :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h2d :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h2e :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h2f :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h30 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h31 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h32 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h33 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h34 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h35 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h36 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h37 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h38 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h39 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h3a :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h3b :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h3c :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h3d :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h3e :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h3f :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h40 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h41 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h42 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h43 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h44 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h45 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h46 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h47 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h48 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h49 :
		RG_quantized_block_rl_34_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h4a :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h4b :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h4c :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h4d :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h4e :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h4f :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h50 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h51 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h52 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h53 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h54 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h55 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h56 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h57 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h58 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h59 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h5a :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h5b :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h5c :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h5d :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h5e :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h5f :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h60 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h61 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h62 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h63 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h64 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h65 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h66 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h67 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h68 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h69 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h6a :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h6b :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h6c :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h6d :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h6e :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h6f :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h70 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h71 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h72 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h73 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h74 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h75 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h76 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h77 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h78 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h79 :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h7a :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h7b :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h7c :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h7d :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h7e :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	7'h7f :
		RG_quantized_block_rl_34_t1 = rl_a73_t8 ;
	default :
		RG_quantized_block_rl_34_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_34_t1 or U_318 or TR_192 or U_317 or RG_rl_75 or 
	ST1_07d or RG_rl_73 or U_88 or jpeg_in_a34 or U_01 or RG_quantized_block_rl_36 or 
	ST1_01d )
	RG_quantized_block_rl_34_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_36 )
		| ( { 9{ U_01 } } & jpeg_in_a34 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_73 )
		| ( { 9{ ST1_07d } } & RG_rl_75 )
		| ( { 9{ U_317 } } & TR_192 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_34_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_34_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_34_en )
		RG_quantized_block_rl_34 <= RG_quantized_block_rl_34_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a75_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h01 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h02 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h03 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h04 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h05 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h06 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h07 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h08 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h09 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h0a :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h0b :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h0c :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h0d :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h0e :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h0f :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h10 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h11 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h12 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h13 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h14 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h15 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h16 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h17 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h18 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h19 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h1a :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h1b :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h1c :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h1d :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h1e :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h1f :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h20 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h21 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h22 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h23 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h24 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h25 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h26 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h27 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h28 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h29 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h2a :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h2b :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h2c :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h2d :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h2e :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h2f :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h30 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h31 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h32 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h33 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h34 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h35 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h36 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h37 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h38 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h39 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h3a :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h3b :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h3c :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h3d :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h3e :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h3f :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h40 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h41 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h42 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h43 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h44 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h45 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h46 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h47 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h48 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h49 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h4a :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h4b :
		RG_quantized_block_rl_35_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h4c :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h4d :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h4e :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h4f :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h50 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h51 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h52 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h53 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h54 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h55 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h56 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h57 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h58 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h59 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h5a :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h5b :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h5c :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h5d :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h5e :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h5f :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h60 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h61 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h62 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h63 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h64 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h65 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h66 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h67 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h68 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h69 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h6a :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h6b :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h6c :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h6d :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h6e :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h6f :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h70 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h71 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h72 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h73 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h74 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h75 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h76 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h77 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h78 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h79 :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h7a :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h7b :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h7c :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h7d :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h7e :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	7'h7f :
		RG_quantized_block_rl_35_t1 = rl_a75_t8 ;
	default :
		RG_quantized_block_rl_35_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_35_t1 or U_318 or TR_190 or U_317 or RG_rl_77 or 
	ST1_07d or RG_rl_75 or U_88 or jpeg_in_a35 or U_01 or RG_quantized_block_rl_37 or 
	ST1_01d )
	RG_quantized_block_rl_35_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_37 )
		| ( { 9{ U_01 } } & jpeg_in_a35 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_75 )
		| ( { 9{ ST1_07d } } & RG_rl_77 )
		| ( { 9{ U_317 } } & TR_190 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_35_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_35_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_35_en )
		RG_quantized_block_rl_35 <= RG_quantized_block_rl_35_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a77_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h01 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h02 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h03 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h04 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h05 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h06 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h07 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h08 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h09 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h0a :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h0b :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h0c :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h0d :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h0e :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h0f :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h10 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h11 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h12 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h13 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h14 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h15 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h16 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h17 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h18 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h19 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h1a :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h1b :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h1c :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h1d :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h1e :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h1f :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h20 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h21 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h22 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h23 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h24 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h25 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h26 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h27 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h28 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h29 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h2a :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h2b :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h2c :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h2d :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h2e :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h2f :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h30 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h31 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h32 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h33 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h34 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h35 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h36 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h37 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h38 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h39 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h3a :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h3b :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h3c :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h3d :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h3e :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h3f :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h40 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h41 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h42 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h43 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h44 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h45 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h46 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h47 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h48 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h49 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h4a :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h4b :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h4c :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h4d :
		RG_quantized_block_rl_36_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h4e :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h4f :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h50 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h51 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h52 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h53 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h54 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h55 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h56 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h57 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h58 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h59 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h5a :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h5b :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h5c :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h5d :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h5e :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h5f :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h60 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h61 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h62 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h63 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h64 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h65 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h66 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h67 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h68 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h69 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h6a :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h6b :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h6c :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h6d :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h6e :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h6f :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h70 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h71 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h72 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h73 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h74 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h75 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h76 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h77 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h78 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h79 :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h7a :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h7b :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h7c :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h7d :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h7e :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	7'h7f :
		RG_quantized_block_rl_36_t1 = rl_a77_t8 ;
	default :
		RG_quantized_block_rl_36_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_36_t1 or U_318 or TR_188 or U_317 or RG_rl_79 or 
	ST1_07d or RG_rl_77 or U_88 or jpeg_in_a36 or U_01 or RG_quantized_block_rl_38 or 
	ST1_01d )
	RG_quantized_block_rl_36_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_38 )
		| ( { 9{ U_01 } } & jpeg_in_a36 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_77 )
		| ( { 9{ ST1_07d } } & RG_rl_79 )
		| ( { 9{ U_317 } } & TR_188 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_36_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_36_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_36_en )
		RG_quantized_block_rl_36 <= RG_quantized_block_rl_36_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a79_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h01 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h02 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h03 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h04 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h05 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h06 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h07 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h08 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h09 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h0a :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h0b :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h0c :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h0d :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h0e :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h0f :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h10 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h11 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h12 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h13 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h14 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h15 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h16 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h17 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h18 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h19 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h1a :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h1b :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h1c :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h1d :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h1e :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h1f :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h20 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h21 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h22 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h23 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h24 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h25 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h26 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h27 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h28 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h29 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h2a :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h2b :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h2c :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h2d :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h2e :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h2f :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h30 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h31 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h32 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h33 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h34 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h35 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h36 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h37 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h38 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h39 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h3a :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h3b :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h3c :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h3d :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h3e :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h3f :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h40 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h41 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h42 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h43 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h44 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h45 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h46 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h47 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h48 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h49 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h4a :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h4b :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h4c :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h4d :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h4e :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h4f :
		RG_quantized_block_rl_37_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h50 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h51 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h52 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h53 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h54 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h55 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h56 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h57 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h58 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h59 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h5a :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h5b :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h5c :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h5d :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h5e :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h5f :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h60 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h61 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h62 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h63 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h64 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h65 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h66 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h67 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h68 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h69 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h6a :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h6b :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h6c :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h6d :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h6e :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h6f :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h70 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h71 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h72 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h73 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h74 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h75 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h76 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h77 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h78 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h79 :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h7a :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h7b :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h7c :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h7d :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h7e :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	7'h7f :
		RG_quantized_block_rl_37_t1 = rl_a79_t8 ;
	default :
		RG_quantized_block_rl_37_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_37_t1 or U_318 or TR_186 or U_317 or RG_rl_81 or 
	ST1_07d or RG_rl_79 or U_88 or jpeg_in_a37 or U_01 or RG_quantized_block_rl_39 or 
	ST1_01d )
	RG_quantized_block_rl_37_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_39 )
		| ( { 9{ U_01 } } & jpeg_in_a37 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_79 )
		| ( { 9{ ST1_07d } } & RG_rl_81 )
		| ( { 9{ U_317 } } & TR_186 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_37_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_37_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_37_en )
		RG_quantized_block_rl_37 <= RG_quantized_block_rl_37_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a81_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h01 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h02 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h03 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h04 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h05 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h06 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h07 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h08 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h09 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h0a :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h0b :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h0c :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h0d :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h0e :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h0f :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h10 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h11 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h12 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h13 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h14 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h15 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h16 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h17 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h18 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h19 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h1a :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h1b :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h1c :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h1d :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h1e :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h1f :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h20 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h21 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h22 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h23 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h24 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h25 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h26 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h27 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h28 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h29 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h2a :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h2b :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h2c :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h2d :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h2e :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h2f :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h30 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h31 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h32 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h33 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h34 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h35 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h36 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h37 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h38 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h39 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h3a :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h3b :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h3c :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h3d :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h3e :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h3f :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h40 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h41 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h42 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h43 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h44 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h45 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h46 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h47 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h48 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h49 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h4a :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h4b :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h4c :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h4d :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h4e :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h4f :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h50 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h51 :
		RG_quantized_block_rl_38_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h52 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h53 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h54 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h55 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h56 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h57 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h58 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h59 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h5a :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h5b :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h5c :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h5d :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h5e :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h5f :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h60 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h61 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h62 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h63 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h64 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h65 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h66 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h67 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h68 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h69 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h6a :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h6b :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h6c :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h6d :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h6e :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h6f :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h70 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h71 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h72 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h73 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h74 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h75 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h76 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h77 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h78 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h79 :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h7a :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h7b :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h7c :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h7d :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h7e :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	7'h7f :
		RG_quantized_block_rl_38_t1 = rl_a81_t8 ;
	default :
		RG_quantized_block_rl_38_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_38_t1 or U_318 or TR_184 or U_317 or RG_rl_83 or 
	ST1_07d or RG_rl_81 or U_88 or jpeg_in_a38 or U_01 or RG_quantized_block_rl_40 or 
	ST1_01d )
	RG_quantized_block_rl_38_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_40 )
		| ( { 9{ U_01 } } & jpeg_in_a38 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_81 )
		| ( { 9{ ST1_07d } } & RG_rl_83 )
		| ( { 9{ U_317 } } & TR_184 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_38_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_38_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_38_en )
		RG_quantized_block_rl_38 <= RG_quantized_block_rl_38_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a83_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h01 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h02 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h03 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h04 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h05 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h06 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h07 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h08 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h09 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h0a :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h0b :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h0c :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h0d :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h0e :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h0f :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h10 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h11 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h12 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h13 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h14 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h15 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h16 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h17 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h18 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h19 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h1a :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h1b :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h1c :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h1d :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h1e :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h1f :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h20 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h21 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h22 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h23 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h24 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h25 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h26 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h27 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h28 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h29 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h2a :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h2b :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h2c :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h2d :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h2e :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h2f :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h30 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h31 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h32 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h33 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h34 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h35 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h36 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h37 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h38 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h39 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h3a :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h3b :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h3c :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h3d :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h3e :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h3f :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h40 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h41 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h42 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h43 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h44 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h45 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h46 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h47 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h48 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h49 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h4a :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h4b :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h4c :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h4d :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h4e :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h4f :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h50 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h51 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h52 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h53 :
		RG_quantized_block_rl_39_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h54 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h55 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h56 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h57 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h58 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h59 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h5a :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h5b :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h5c :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h5d :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h5e :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h5f :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h60 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h61 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h62 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h63 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h64 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h65 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h66 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h67 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h68 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h69 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h6a :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h6b :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h6c :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h6d :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h6e :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h6f :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h70 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h71 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h72 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h73 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h74 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h75 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h76 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h77 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h78 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h79 :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h7a :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h7b :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h7c :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h7d :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h7e :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	7'h7f :
		RG_quantized_block_rl_39_t1 = rl_a83_t8 ;
	default :
		RG_quantized_block_rl_39_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_39_t1 or U_318 or TR_182 or U_317 or RG_rl_85 or 
	ST1_07d or RG_rl_83 or U_88 or jpeg_in_a39 or U_01 or RG_quantized_block_rl_41 or 
	ST1_01d )
	RG_quantized_block_rl_39_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_41 )
		| ( { 9{ U_01 } } & jpeg_in_a39 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_83 )
		| ( { 9{ ST1_07d } } & RG_rl_85 )
		| ( { 9{ U_317 } } & TR_182 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_39_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_39_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_39_en )
		RG_quantized_block_rl_39 <= RG_quantized_block_rl_39_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a85_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h01 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h02 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h03 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h04 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h05 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h06 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h07 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h08 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h09 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h0a :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h0b :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h0c :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h0d :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h0e :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h0f :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h10 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h11 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h12 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h13 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h14 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h15 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h16 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h17 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h18 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h19 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h1a :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h1b :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h1c :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h1d :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h1e :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h1f :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h20 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h21 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h22 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h23 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h24 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h25 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h26 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h27 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h28 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h29 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h2a :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h2b :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h2c :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h2d :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h2e :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h2f :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h30 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h31 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h32 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h33 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h34 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h35 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h36 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h37 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h38 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h39 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h3a :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h3b :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h3c :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h3d :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h3e :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h3f :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h40 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h41 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h42 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h43 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h44 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h45 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h46 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h47 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h48 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h49 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h4a :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h4b :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h4c :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h4d :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h4e :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h4f :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h50 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h51 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h52 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h53 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h54 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h55 :
		RG_quantized_block_rl_40_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h56 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h57 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h58 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h59 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h5a :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h5b :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h5c :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h5d :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h5e :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h5f :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h60 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h61 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h62 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h63 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h64 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h65 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h66 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h67 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h68 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h69 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h6a :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h6b :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h6c :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h6d :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h6e :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h6f :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h70 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h71 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h72 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h73 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h74 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h75 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h76 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h77 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h78 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h79 :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h7a :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h7b :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h7c :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h7d :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h7e :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	7'h7f :
		RG_quantized_block_rl_40_t1 = rl_a85_t8 ;
	default :
		RG_quantized_block_rl_40_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_40_t1 or U_318 or TR_180 or U_317 or RG_rl_87 or 
	ST1_07d or RG_rl_85 or U_88 or jpeg_in_a40 or U_01 or RG_quantized_block_rl_42 or 
	ST1_01d )
	RG_quantized_block_rl_40_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_42 )
		| ( { 9{ U_01 } } & jpeg_in_a40 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_85 )
		| ( { 9{ ST1_07d } } & RG_rl_87 )
		| ( { 9{ U_317 } } & TR_180 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_40_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_40_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_40_en )
		RG_quantized_block_rl_40 <= RG_quantized_block_rl_40_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a87_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h01 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h02 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h03 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h04 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h05 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h06 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h07 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h08 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h09 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h0a :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h0b :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h0c :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h0d :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h0e :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h0f :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h10 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h11 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h12 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h13 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h14 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h15 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h16 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h17 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h18 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h19 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h1a :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h1b :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h1c :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h1d :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h1e :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h1f :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h20 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h21 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h22 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h23 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h24 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h25 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h26 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h27 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h28 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h29 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h2a :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h2b :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h2c :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h2d :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h2e :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h2f :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h30 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h31 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h32 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h33 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h34 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h35 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h36 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h37 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h38 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h39 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h3a :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h3b :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h3c :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h3d :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h3e :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h3f :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h40 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h41 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h42 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h43 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h44 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h45 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h46 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h47 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h48 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h49 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h4a :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h4b :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h4c :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h4d :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h4e :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h4f :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h50 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h51 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h52 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h53 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h54 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h55 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h56 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h57 :
		RG_quantized_block_rl_41_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h58 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h59 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h5a :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h5b :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h5c :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h5d :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h5e :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h5f :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h60 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h61 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h62 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h63 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h64 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h65 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h66 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h67 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h68 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h69 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h6a :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h6b :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h6c :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h6d :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h6e :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h6f :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h70 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h71 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h72 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h73 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h74 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h75 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h76 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h77 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h78 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h79 :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h7a :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h7b :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h7c :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h7d :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h7e :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	7'h7f :
		RG_quantized_block_rl_41_t1 = rl_a87_t8 ;
	default :
		RG_quantized_block_rl_41_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_41_t1 or U_318 or TR_178 or U_317 or RG_rl_89 or 
	ST1_07d or RG_rl_87 or U_88 or jpeg_in_a41 or U_01 or RG_quantized_block_rl_43 or 
	ST1_01d )
	RG_quantized_block_rl_41_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_43 )
		| ( { 9{ U_01 } } & jpeg_in_a41 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_87 )
		| ( { 9{ ST1_07d } } & RG_rl_89 )
		| ( { 9{ U_317 } } & TR_178 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_41_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_41_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_41_en )
		RG_quantized_block_rl_41 <= RG_quantized_block_rl_41_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a89_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h01 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h02 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h03 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h04 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h05 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h06 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h07 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h08 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h09 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h0a :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h0b :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h0c :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h0d :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h0e :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h0f :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h10 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h11 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h12 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h13 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h14 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h15 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h16 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h17 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h18 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h19 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h1a :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h1b :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h1c :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h1d :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h1e :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h1f :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h20 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h21 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h22 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h23 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h24 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h25 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h26 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h27 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h28 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h29 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h2a :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h2b :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h2c :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h2d :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h2e :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h2f :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h30 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h31 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h32 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h33 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h34 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h35 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h36 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h37 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h38 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h39 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h3a :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h3b :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h3c :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h3d :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h3e :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h3f :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h40 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h41 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h42 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h43 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h44 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h45 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h46 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h47 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h48 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h49 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h4a :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h4b :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h4c :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h4d :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h4e :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h4f :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h50 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h51 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h52 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h53 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h54 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h55 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h56 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h57 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h58 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h59 :
		RG_quantized_block_rl_42_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h5a :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h5b :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h5c :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h5d :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h5e :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h5f :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h60 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h61 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h62 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h63 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h64 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h65 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h66 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h67 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h68 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h69 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h6a :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h6b :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h6c :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h6d :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h6e :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h6f :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h70 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h71 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h72 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h73 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h74 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h75 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h76 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h77 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h78 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h79 :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h7a :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h7b :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h7c :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h7d :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h7e :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	7'h7f :
		RG_quantized_block_rl_42_t1 = rl_a89_t8 ;
	default :
		RG_quantized_block_rl_42_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_42_t1 or U_318 or TR_176 or U_317 or RG_rl_91 or 
	ST1_07d or RG_rl_89 or U_88 or jpeg_in_a42 or U_01 or RG_quantized_block_rl_44 or 
	ST1_01d )
	RG_quantized_block_rl_42_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_44 )
		| ( { 9{ U_01 } } & jpeg_in_a42 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_89 )
		| ( { 9{ ST1_07d } } & RG_rl_91 )
		| ( { 9{ U_317 } } & TR_176 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_42_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_42_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_42_en )
		RG_quantized_block_rl_42 <= RG_quantized_block_rl_42_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a91_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h01 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h02 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h03 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h04 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h05 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h06 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h07 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h08 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h09 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h0a :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h0b :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h0c :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h0d :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h0e :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h0f :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h10 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h11 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h12 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h13 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h14 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h15 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h16 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h17 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h18 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h19 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h1a :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h1b :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h1c :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h1d :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h1e :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h1f :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h20 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h21 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h22 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h23 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h24 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h25 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h26 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h27 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h28 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h29 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h2a :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h2b :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h2c :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h2d :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h2e :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h2f :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h30 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h31 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h32 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h33 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h34 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h35 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h36 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h37 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h38 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h39 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h3a :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h3b :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h3c :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h3d :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h3e :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h3f :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h40 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h41 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h42 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h43 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h44 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h45 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h46 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h47 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h48 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h49 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h4a :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h4b :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h4c :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h4d :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h4e :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h4f :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h50 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h51 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h52 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h53 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h54 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h55 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h56 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h57 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h58 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h59 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h5a :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h5b :
		RG_quantized_block_rl_43_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h5c :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h5d :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h5e :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h5f :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h60 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h61 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h62 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h63 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h64 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h65 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h66 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h67 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h68 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h69 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h6a :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h6b :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h6c :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h6d :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h6e :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h6f :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h70 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h71 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h72 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h73 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h74 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h75 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h76 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h77 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h78 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h79 :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h7a :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h7b :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h7c :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h7d :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h7e :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	7'h7f :
		RG_quantized_block_rl_43_t1 = rl_a91_t8 ;
	default :
		RG_quantized_block_rl_43_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_43_t1 or U_318 or TR_174 or U_317 or RG_rl_93 or 
	ST1_07d or RG_rl_91 or U_88 or jpeg_in_a43 or U_01 or RG_quantized_block_rl_45 or 
	ST1_01d )
	RG_quantized_block_rl_43_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_45 )
		| ( { 9{ U_01 } } & jpeg_in_a43 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_91 )
		| ( { 9{ ST1_07d } } & RG_rl_93 )
		| ( { 9{ U_317 } } & TR_174 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_43_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_43_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_43_en )
		RG_quantized_block_rl_43 <= RG_quantized_block_rl_43_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a93_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h01 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h02 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h03 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h04 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h05 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h06 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h07 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h08 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h09 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h0a :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h0b :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h0c :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h0d :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h0e :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h0f :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h10 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h11 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h12 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h13 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h14 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h15 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h16 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h17 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h18 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h19 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h1a :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h1b :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h1c :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h1d :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h1e :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h1f :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h20 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h21 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h22 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h23 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h24 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h25 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h26 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h27 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h28 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h29 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h2a :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h2b :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h2c :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h2d :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h2e :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h2f :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h30 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h31 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h32 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h33 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h34 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h35 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h36 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h37 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h38 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h39 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h3a :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h3b :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h3c :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h3d :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h3e :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h3f :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h40 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h41 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h42 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h43 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h44 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h45 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h46 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h47 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h48 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h49 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h4a :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h4b :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h4c :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h4d :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h4e :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h4f :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h50 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h51 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h52 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h53 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h54 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h55 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h56 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h57 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h58 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h59 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h5a :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h5b :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h5c :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h5d :
		RG_quantized_block_rl_44_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h5e :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h5f :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h60 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h61 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h62 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h63 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h64 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h65 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h66 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h67 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h68 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h69 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h6a :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h6b :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h6c :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h6d :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h6e :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h6f :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h70 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h71 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h72 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h73 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h74 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h75 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h76 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h77 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h78 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h79 :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h7a :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h7b :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h7c :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h7d :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h7e :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	7'h7f :
		RG_quantized_block_rl_44_t1 = rl_a93_t8 ;
	default :
		RG_quantized_block_rl_44_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_44_t1 or U_318 or TR_172 or U_317 or RG_rl_95 or 
	ST1_07d or RG_rl_93 or U_88 or jpeg_in_a44 or U_01 or RG_quantized_block_rl_46 or 
	ST1_01d )
	RG_quantized_block_rl_44_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_46 )
		| ( { 9{ U_01 } } & jpeg_in_a44 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_93 )
		| ( { 9{ ST1_07d } } & RG_rl_95 )
		| ( { 9{ U_317 } } & TR_172 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_44_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_44_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_44_en )
		RG_quantized_block_rl_44 <= RG_quantized_block_rl_44_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a95_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h01 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h02 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h03 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h04 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h05 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h06 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h07 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h08 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h09 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h0a :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h0b :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h0c :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h0d :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h0e :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h0f :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h10 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h11 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h12 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h13 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h14 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h15 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h16 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h17 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h18 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h19 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h1a :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h1b :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h1c :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h1d :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h1e :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h1f :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h20 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h21 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h22 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h23 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h24 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h25 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h26 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h27 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h28 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h29 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h2a :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h2b :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h2c :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h2d :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h2e :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h2f :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h30 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h31 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h32 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h33 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h34 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h35 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h36 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h37 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h38 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h39 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h3a :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h3b :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h3c :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h3d :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h3e :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h3f :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h40 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h41 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h42 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h43 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h44 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h45 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h46 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h47 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h48 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h49 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h4a :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h4b :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h4c :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h4d :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h4e :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h4f :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h50 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h51 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h52 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h53 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h54 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h55 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h56 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h57 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h58 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h59 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h5a :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h5b :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h5c :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h5d :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h5e :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h5f :
		RG_quantized_block_rl_45_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h60 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h61 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h62 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h63 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h64 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h65 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h66 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h67 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h68 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h69 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h6a :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h6b :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h6c :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h6d :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h6e :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h6f :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h70 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h71 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h72 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h73 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h74 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h75 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h76 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h77 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h78 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h79 :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h7a :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h7b :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h7c :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h7d :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h7e :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	7'h7f :
		RG_quantized_block_rl_45_t1 = rl_a95_t8 ;
	default :
		RG_quantized_block_rl_45_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_45_t1 or U_318 or TR_170 or U_317 or RG_rl_97 or 
	ST1_07d or RG_rl_95 or U_88 or jpeg_in_a45 or U_01 or RG_quantized_block_rl_47 or 
	ST1_01d )
	RG_quantized_block_rl_45_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_47 )
		| ( { 9{ U_01 } } & jpeg_in_a45 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_95 )
		| ( { 9{ ST1_07d } } & RG_rl_97 )
		| ( { 9{ U_317 } } & TR_170 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_45_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_45_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_45_en )
		RG_quantized_block_rl_45 <= RG_quantized_block_rl_45_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a97_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h01 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h02 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h03 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h04 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h05 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h06 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h07 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h08 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h09 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h0a :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h0b :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h0c :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h0d :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h0e :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h0f :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h10 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h11 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h12 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h13 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h14 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h15 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h16 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h17 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h18 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h19 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h1a :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h1b :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h1c :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h1d :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h1e :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h1f :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h20 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h21 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h22 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h23 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h24 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h25 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h26 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h27 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h28 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h29 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h2a :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h2b :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h2c :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h2d :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h2e :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h2f :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h30 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h31 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h32 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h33 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h34 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h35 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h36 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h37 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h38 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h39 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h3a :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h3b :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h3c :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h3d :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h3e :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h3f :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h40 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h41 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h42 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h43 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h44 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h45 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h46 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h47 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h48 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h49 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h4a :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h4b :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h4c :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h4d :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h4e :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h4f :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h50 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h51 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h52 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h53 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h54 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h55 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h56 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h57 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h58 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h59 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h5a :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h5b :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h5c :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h5d :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h5e :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h5f :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h60 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h61 :
		RG_quantized_block_rl_46_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h62 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h63 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h64 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h65 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h66 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h67 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h68 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h69 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h6a :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h6b :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h6c :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h6d :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h6e :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h6f :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h70 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h71 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h72 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h73 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h74 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h75 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h76 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h77 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h78 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h79 :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h7a :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h7b :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h7c :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h7d :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h7e :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	7'h7f :
		RG_quantized_block_rl_46_t1 = rl_a97_t8 ;
	default :
		RG_quantized_block_rl_46_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_46_t1 or U_318 or TR_168 or U_317 or RG_rl_99 or 
	ST1_07d or RG_rl_97 or U_88 or jpeg_in_a46 or U_01 or RG_quantized_block_rl_48 or 
	ST1_01d )
	RG_quantized_block_rl_46_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_48 )
		| ( { 9{ U_01 } } & jpeg_in_a46 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_97 )
		| ( { 9{ ST1_07d } } & RG_rl_99 )
		| ( { 9{ U_317 } } & TR_168 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_46_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_46_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_46_en )
		RG_quantized_block_rl_46 <= RG_quantized_block_rl_46_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a99_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h01 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h02 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h03 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h04 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h05 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h06 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h07 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h08 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h09 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h0a :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h0b :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h0c :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h0d :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h0e :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h0f :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h10 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h11 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h12 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h13 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h14 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h15 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h16 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h17 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h18 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h19 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h1a :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h1b :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h1c :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h1d :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h1e :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h1f :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h20 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h21 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h22 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h23 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h24 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h25 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h26 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h27 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h28 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h29 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h2a :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h2b :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h2c :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h2d :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h2e :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h2f :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h30 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h31 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h32 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h33 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h34 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h35 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h36 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h37 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h38 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h39 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h3a :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h3b :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h3c :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h3d :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h3e :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h3f :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h40 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h41 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h42 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h43 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h44 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h45 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h46 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h47 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h48 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h49 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h4a :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h4b :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h4c :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h4d :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h4e :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h4f :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h50 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h51 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h52 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h53 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h54 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h55 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h56 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h57 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h58 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h59 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h5a :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h5b :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h5c :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h5d :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h5e :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h5f :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h60 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h61 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h62 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h63 :
		RG_quantized_block_rl_47_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h64 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h65 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h66 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h67 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h68 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h69 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h6a :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h6b :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h6c :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h6d :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h6e :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h6f :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h70 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h71 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h72 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h73 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h74 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h75 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h76 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h77 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h78 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h79 :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h7a :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h7b :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h7c :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h7d :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h7e :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	7'h7f :
		RG_quantized_block_rl_47_t1 = rl_a99_t8 ;
	default :
		RG_quantized_block_rl_47_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_47_t1 or U_318 or TR_166 or U_317 or RG_rl_101 or 
	ST1_07d or RG_rl_99 or U_88 or jpeg_in_a47 or U_01 or RG_quantized_block_rl_49 or 
	ST1_01d )
	RG_quantized_block_rl_47_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_49 )
		| ( { 9{ U_01 } } & jpeg_in_a47 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_99 )
		| ( { 9{ ST1_07d } } & RG_rl_101 )
		| ( { 9{ U_317 } } & TR_166 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_47_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_47_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_47_en )
		RG_quantized_block_rl_47 <= RG_quantized_block_rl_47_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a101_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h01 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h02 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h03 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h04 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h05 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h06 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h07 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h08 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h09 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h0a :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h0b :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h0c :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h0d :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h0e :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h0f :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h10 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h11 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h12 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h13 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h14 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h15 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h16 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h17 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h18 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h19 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h1a :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h1b :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h1c :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h1d :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h1e :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h1f :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h20 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h21 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h22 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h23 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h24 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h25 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h26 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h27 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h28 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h29 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h2a :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h2b :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h2c :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h2d :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h2e :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h2f :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h30 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h31 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h32 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h33 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h34 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h35 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h36 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h37 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h38 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h39 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h3a :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h3b :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h3c :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h3d :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h3e :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h3f :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h40 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h41 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h42 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h43 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h44 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h45 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h46 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h47 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h48 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h49 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h4a :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h4b :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h4c :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h4d :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h4e :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h4f :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h50 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h51 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h52 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h53 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h54 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h55 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h56 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h57 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h58 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h59 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h5a :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h5b :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h5c :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h5d :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h5e :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h5f :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h60 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h61 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h62 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h63 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h64 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h65 :
		RG_quantized_block_rl_48_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h66 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h67 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h68 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h69 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h6a :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h6b :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h6c :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h6d :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h6e :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h6f :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h70 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h71 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h72 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h73 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h74 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h75 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h76 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h77 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h78 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h79 :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h7a :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h7b :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h7c :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h7d :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h7e :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	7'h7f :
		RG_quantized_block_rl_48_t1 = rl_a101_t8 ;
	default :
		RG_quantized_block_rl_48_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_48_t1 or U_318 or TR_164 or U_317 or RG_rl_103 or 
	ST1_07d or RG_rl_101 or U_88 or jpeg_in_a48 or U_01 or RG_quantized_block_rl_50 or 
	ST1_01d )
	RG_quantized_block_rl_48_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_50 )
		| ( { 9{ U_01 } } & jpeg_in_a48 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_101 )
		| ( { 9{ ST1_07d } } & RG_rl_103 )
		| ( { 9{ U_317 } } & TR_164 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_48_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_48_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_48_en )
		RG_quantized_block_rl_48 <= RG_quantized_block_rl_48_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a103_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h01 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h02 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h03 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h04 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h05 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h06 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h07 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h08 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h09 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h0a :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h0b :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h0c :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h0d :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h0e :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h0f :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h10 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h11 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h12 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h13 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h14 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h15 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h16 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h17 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h18 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h19 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h1a :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h1b :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h1c :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h1d :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h1e :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h1f :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h20 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h21 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h22 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h23 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h24 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h25 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h26 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h27 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h28 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h29 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h2a :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h2b :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h2c :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h2d :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h2e :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h2f :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h30 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h31 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h32 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h33 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h34 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h35 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h36 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h37 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h38 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h39 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h3a :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h3b :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h3c :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h3d :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h3e :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h3f :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h40 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h41 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h42 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h43 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h44 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h45 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h46 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h47 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h48 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h49 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h4a :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h4b :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h4c :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h4d :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h4e :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h4f :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h50 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h51 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h52 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h53 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h54 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h55 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h56 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h57 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h58 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h59 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h5a :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h5b :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h5c :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h5d :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h5e :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h5f :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h60 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h61 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h62 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h63 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h64 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h65 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h66 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h67 :
		RG_quantized_block_rl_49_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h68 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h69 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h6a :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h6b :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h6c :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h6d :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h6e :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h6f :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h70 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h71 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h72 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h73 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h74 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h75 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h76 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h77 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h78 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h79 :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h7a :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h7b :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h7c :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h7d :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h7e :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	7'h7f :
		RG_quantized_block_rl_49_t1 = rl_a103_t8 ;
	default :
		RG_quantized_block_rl_49_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_49_t1 or U_318 or TR_162 or U_317 or RG_rl_105 or 
	ST1_07d or RG_rl_103 or U_88 or jpeg_in_a49 or U_01 or RG_quantized_block_rl_51 or 
	ST1_01d )
	RG_quantized_block_rl_49_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_51 )
		| ( { 9{ U_01 } } & jpeg_in_a49 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_103 )
		| ( { 9{ ST1_07d } } & RG_rl_105 )
		| ( { 9{ U_317 } } & TR_162 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_49_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_49_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_49_en )
		RG_quantized_block_rl_49 <= RG_quantized_block_rl_49_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a105_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h01 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h02 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h03 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h04 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h05 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h06 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h07 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h08 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h09 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h0a :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h0b :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h0c :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h0d :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h0e :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h0f :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h10 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h11 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h12 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h13 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h14 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h15 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h16 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h17 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h18 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h19 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h1a :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h1b :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h1c :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h1d :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h1e :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h1f :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h20 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h21 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h22 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h23 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h24 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h25 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h26 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h27 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h28 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h29 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h2a :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h2b :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h2c :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h2d :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h2e :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h2f :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h30 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h31 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h32 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h33 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h34 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h35 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h36 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h37 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h38 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h39 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h3a :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h3b :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h3c :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h3d :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h3e :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h3f :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h40 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h41 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h42 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h43 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h44 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h45 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h46 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h47 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h48 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h49 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h4a :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h4b :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h4c :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h4d :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h4e :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h4f :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h50 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h51 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h52 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h53 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h54 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h55 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h56 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h57 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h58 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h59 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h5a :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h5b :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h5c :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h5d :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h5e :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h5f :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h60 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h61 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h62 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h63 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h64 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h65 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h66 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h67 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h68 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h69 :
		RG_quantized_block_rl_50_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h6a :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h6b :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h6c :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h6d :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h6e :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h6f :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h70 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h71 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h72 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h73 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h74 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h75 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h76 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h77 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h78 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h79 :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h7a :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h7b :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h7c :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h7d :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h7e :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	7'h7f :
		RG_quantized_block_rl_50_t1 = rl_a105_t8 ;
	default :
		RG_quantized_block_rl_50_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_50_t1 or U_318 or TR_160 or U_317 or RG_rl_107 or 
	ST1_07d or RG_rl_105 or U_88 or jpeg_in_a50 or U_01 or RG_quantized_block_rl_52 or 
	ST1_01d )
	RG_quantized_block_rl_50_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_52 )
		| ( { 9{ U_01 } } & jpeg_in_a50 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_105 )
		| ( { 9{ ST1_07d } } & RG_rl_107 )
		| ( { 9{ U_317 } } & TR_160 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_50_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_50_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_50_en )
		RG_quantized_block_rl_50 <= RG_quantized_block_rl_50_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a107_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h01 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h02 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h03 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h04 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h05 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h06 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h07 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h08 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h09 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h0a :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h0b :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h0c :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h0d :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h0e :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h0f :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h10 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h11 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h12 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h13 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h14 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h15 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h16 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h17 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h18 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h19 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h1a :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h1b :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h1c :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h1d :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h1e :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h1f :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h20 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h21 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h22 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h23 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h24 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h25 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h26 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h27 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h28 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h29 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h2a :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h2b :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h2c :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h2d :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h2e :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h2f :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h30 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h31 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h32 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h33 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h34 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h35 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h36 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h37 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h38 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h39 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h3a :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h3b :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h3c :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h3d :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h3e :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h3f :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h40 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h41 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h42 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h43 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h44 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h45 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h46 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h47 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h48 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h49 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h4a :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h4b :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h4c :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h4d :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h4e :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h4f :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h50 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h51 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h52 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h53 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h54 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h55 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h56 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h57 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h58 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h59 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h5a :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h5b :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h5c :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h5d :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h5e :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h5f :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h60 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h61 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h62 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h63 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h64 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h65 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h66 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h67 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h68 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h69 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h6a :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h6b :
		RG_quantized_block_rl_51_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h6c :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h6d :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h6e :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h6f :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h70 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h71 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h72 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h73 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h74 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h75 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h76 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h77 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h78 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h79 :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h7a :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h7b :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h7c :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h7d :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h7e :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	7'h7f :
		RG_quantized_block_rl_51_t1 = rl_a107_t8 ;
	default :
		RG_quantized_block_rl_51_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_51_t1 or U_318 or TR_158 or U_317 or RG_rl_109 or 
	ST1_07d or RG_rl_107 or U_88 or jpeg_in_a51 or U_01 or RG_quantized_block_rl_53 or 
	ST1_01d )
	RG_quantized_block_rl_51_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_53 )
		| ( { 9{ U_01 } } & jpeg_in_a51 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_107 )
		| ( { 9{ ST1_07d } } & RG_rl_109 )
		| ( { 9{ U_317 } } & TR_158 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_51_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_51_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_51_en )
		RG_quantized_block_rl_51 <= RG_quantized_block_rl_51_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a109_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h01 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h02 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h03 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h04 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h05 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h06 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h07 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h08 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h09 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h0a :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h0b :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h0c :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h0d :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h0e :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h0f :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h10 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h11 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h12 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h13 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h14 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h15 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h16 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h17 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h18 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h19 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h1a :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h1b :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h1c :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h1d :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h1e :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h1f :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h20 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h21 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h22 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h23 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h24 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h25 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h26 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h27 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h28 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h29 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h2a :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h2b :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h2c :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h2d :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h2e :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h2f :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h30 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h31 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h32 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h33 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h34 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h35 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h36 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h37 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h38 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h39 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h3a :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h3b :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h3c :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h3d :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h3e :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h3f :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h40 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h41 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h42 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h43 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h44 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h45 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h46 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h47 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h48 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h49 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h4a :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h4b :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h4c :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h4d :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h4e :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h4f :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h50 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h51 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h52 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h53 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h54 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h55 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h56 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h57 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h58 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h59 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h5a :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h5b :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h5c :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h5d :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h5e :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h5f :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h60 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h61 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h62 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h63 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h64 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h65 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h66 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h67 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h68 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h69 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h6a :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h6b :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h6c :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h6d :
		RG_quantized_block_rl_52_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h6e :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h6f :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h70 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h71 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h72 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h73 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h74 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h75 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h76 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h77 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h78 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h79 :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h7a :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h7b :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h7c :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h7d :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h7e :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	7'h7f :
		RG_quantized_block_rl_52_t1 = rl_a109_t8 ;
	default :
		RG_quantized_block_rl_52_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_52_t1 or U_318 or TR_156 or U_317 or RG_rl_111 or 
	ST1_07d or RG_rl_109 or U_88 or jpeg_in_a52 or U_01 or RG_quantized_block_rl_54 or 
	ST1_01d )
	RG_quantized_block_rl_52_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_54 )
		| ( { 9{ U_01 } } & jpeg_in_a52 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_109 )
		| ( { 9{ ST1_07d } } & RG_rl_111 )
		| ( { 9{ U_317 } } & TR_156 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_52_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_52_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_52_en )
		RG_quantized_block_rl_52 <= RG_quantized_block_rl_52_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a111_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h01 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h02 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h03 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h04 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h05 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h06 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h07 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h08 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h09 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h0a :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h0b :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h0c :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h0d :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h0e :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h0f :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h10 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h11 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h12 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h13 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h14 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h15 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h16 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h17 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h18 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h19 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h1a :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h1b :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h1c :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h1d :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h1e :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h1f :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h20 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h21 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h22 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h23 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h24 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h25 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h26 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h27 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h28 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h29 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h2a :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h2b :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h2c :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h2d :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h2e :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h2f :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h30 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h31 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h32 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h33 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h34 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h35 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h36 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h37 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h38 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h39 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h3a :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h3b :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h3c :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h3d :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h3e :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h3f :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h40 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h41 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h42 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h43 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h44 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h45 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h46 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h47 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h48 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h49 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h4a :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h4b :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h4c :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h4d :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h4e :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h4f :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h50 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h51 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h52 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h53 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h54 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h55 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h56 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h57 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h58 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h59 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h5a :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h5b :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h5c :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h5d :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h5e :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h5f :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h60 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h61 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h62 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h63 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h64 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h65 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h66 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h67 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h68 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h69 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h6a :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h6b :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h6c :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h6d :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h6e :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h6f :
		RG_quantized_block_rl_53_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h70 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h71 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h72 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h73 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h74 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h75 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h76 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h77 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h78 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h79 :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h7a :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h7b :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h7c :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h7d :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h7e :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	7'h7f :
		RG_quantized_block_rl_53_t1 = rl_a111_t8 ;
	default :
		RG_quantized_block_rl_53_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_53_t1 or U_318 or TR_154 or U_317 or RG_rl_113 or 
	ST1_07d or RG_rl_111 or U_88 or jpeg_in_a53 or U_01 or RG_quantized_block_rl_55 or 
	ST1_01d )
	RG_quantized_block_rl_53_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_55 )
		| ( { 9{ U_01 } } & jpeg_in_a53 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_111 )
		| ( { 9{ ST1_07d } } & RG_rl_113 )
		| ( { 9{ U_317 } } & TR_154 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_53_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_53_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_53_en )
		RG_quantized_block_rl_53 <= RG_quantized_block_rl_53_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a113_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h01 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h02 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h03 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h04 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h05 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h06 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h07 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h08 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h09 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h0a :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h0b :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h0c :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h0d :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h0e :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h0f :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h10 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h11 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h12 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h13 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h14 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h15 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h16 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h17 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h18 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h19 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h1a :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h1b :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h1c :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h1d :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h1e :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h1f :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h20 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h21 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h22 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h23 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h24 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h25 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h26 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h27 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h28 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h29 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h2a :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h2b :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h2c :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h2d :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h2e :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h2f :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h30 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h31 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h32 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h33 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h34 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h35 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h36 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h37 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h38 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h39 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h3a :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h3b :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h3c :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h3d :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h3e :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h3f :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h40 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h41 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h42 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h43 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h44 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h45 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h46 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h47 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h48 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h49 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h4a :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h4b :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h4c :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h4d :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h4e :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h4f :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h50 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h51 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h52 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h53 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h54 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h55 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h56 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h57 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h58 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h59 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h5a :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h5b :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h5c :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h5d :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h5e :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h5f :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h60 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h61 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h62 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h63 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h64 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h65 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h66 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h67 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h68 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h69 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h6a :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h6b :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h6c :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h6d :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h6e :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h6f :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h70 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h71 :
		RG_quantized_block_rl_54_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h72 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h73 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h74 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h75 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h76 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h77 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h78 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h79 :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h7a :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h7b :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h7c :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h7d :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h7e :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	7'h7f :
		RG_quantized_block_rl_54_t1 = rl_a113_t8 ;
	default :
		RG_quantized_block_rl_54_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_54_t1 or U_318 or TR_152 or U_317 or RG_rl_115 or 
	ST1_07d or RG_rl_113 or U_88 or jpeg_in_a54 or U_01 or RG_quantized_block_rl_56 or 
	ST1_01d )
	RG_quantized_block_rl_54_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_56 )
		| ( { 9{ U_01 } } & jpeg_in_a54 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_113 )
		| ( { 9{ ST1_07d } } & RG_rl_115 )
		| ( { 9{ U_317 } } & TR_152 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_54_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_54_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_54_en )
		RG_quantized_block_rl_54 <= RG_quantized_block_rl_54_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a115_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h01 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h02 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h03 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h04 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h05 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h06 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h07 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h08 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h09 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h0a :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h0b :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h0c :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h0d :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h0e :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h0f :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h10 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h11 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h12 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h13 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h14 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h15 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h16 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h17 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h18 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h19 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h1a :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h1b :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h1c :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h1d :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h1e :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h1f :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h20 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h21 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h22 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h23 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h24 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h25 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h26 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h27 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h28 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h29 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h2a :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h2b :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h2c :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h2d :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h2e :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h2f :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h30 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h31 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h32 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h33 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h34 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h35 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h36 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h37 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h38 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h39 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h3a :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h3b :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h3c :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h3d :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h3e :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h3f :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h40 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h41 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h42 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h43 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h44 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h45 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h46 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h47 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h48 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h49 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h4a :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h4b :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h4c :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h4d :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h4e :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h4f :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h50 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h51 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h52 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h53 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h54 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h55 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h56 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h57 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h58 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h59 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h5a :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h5b :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h5c :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h5d :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h5e :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h5f :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h60 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h61 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h62 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h63 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h64 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h65 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h66 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h67 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h68 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h69 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h6a :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h6b :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h6c :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h6d :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h6e :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h6f :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h70 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h71 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h72 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h73 :
		RG_quantized_block_rl_55_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h74 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h75 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h76 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h77 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h78 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h79 :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h7a :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h7b :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h7c :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h7d :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h7e :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	7'h7f :
		RG_quantized_block_rl_55_t1 = rl_a115_t8 ;
	default :
		RG_quantized_block_rl_55_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_55_t1 or U_318 or TR_150 or U_317 or RG_rl_117 or 
	ST1_07d or RG_rl_115 or U_88 or jpeg_in_a55 or U_01 or RG_quantized_block_rl_57 or 
	ST1_01d )
	RG_quantized_block_rl_55_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_57 )
		| ( { 9{ U_01 } } & jpeg_in_a55 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_115 )
		| ( { 9{ ST1_07d } } & RG_rl_117 )
		| ( { 9{ U_317 } } & TR_150 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_55_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_55_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_55_en )
		RG_quantized_block_rl_55 <= RG_quantized_block_rl_55_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a117_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h01 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h02 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h03 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h04 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h05 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h06 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h07 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h08 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h09 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h0a :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h0b :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h0c :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h0d :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h0e :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h0f :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h10 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h11 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h12 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h13 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h14 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h15 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h16 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h17 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h18 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h19 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h1a :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h1b :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h1c :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h1d :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h1e :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h1f :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h20 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h21 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h22 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h23 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h24 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h25 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h26 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h27 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h28 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h29 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h2a :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h2b :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h2c :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h2d :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h2e :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h2f :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h30 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h31 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h32 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h33 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h34 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h35 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h36 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h37 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h38 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h39 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h3a :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h3b :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h3c :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h3d :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h3e :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h3f :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h40 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h41 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h42 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h43 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h44 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h45 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h46 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h47 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h48 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h49 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h4a :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h4b :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h4c :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h4d :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h4e :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h4f :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h50 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h51 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h52 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h53 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h54 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h55 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h56 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h57 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h58 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h59 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h5a :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h5b :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h5c :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h5d :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h5e :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h5f :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h60 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h61 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h62 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h63 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h64 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h65 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h66 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h67 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h68 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h69 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h6a :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h6b :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h6c :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h6d :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h6e :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h6f :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h70 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h71 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h72 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h73 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h74 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h75 :
		RG_quantized_block_rl_56_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h76 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h77 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h78 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h79 :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h7a :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h7b :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h7c :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h7d :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h7e :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	7'h7f :
		RG_quantized_block_rl_56_t1 = rl_a117_t8 ;
	default :
		RG_quantized_block_rl_56_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_56_t1 or U_318 or TR_148 or U_317 or RG_rl_119 or 
	ST1_07d or RG_rl_117 or U_88 or jpeg_in_a56 or U_01 or RG_quantized_block_rl_58 or 
	ST1_01d )
	RG_quantized_block_rl_56_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_58 )
		| ( { 9{ U_01 } } & jpeg_in_a56 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_117 )
		| ( { 9{ ST1_07d } } & RG_rl_119 )
		| ( { 9{ U_317 } } & TR_148 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_56_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_56_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_56_en )
		RG_quantized_block_rl_56 <= RG_quantized_block_rl_56_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a119_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h01 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h02 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h03 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h04 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h05 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h06 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h07 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h08 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h09 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h0a :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h0b :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h0c :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h0d :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h0e :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h0f :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h10 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h11 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h12 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h13 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h14 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h15 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h16 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h17 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h18 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h19 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h1a :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h1b :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h1c :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h1d :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h1e :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h1f :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h20 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h21 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h22 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h23 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h24 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h25 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h26 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h27 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h28 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h29 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h2a :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h2b :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h2c :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h2d :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h2e :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h2f :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h30 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h31 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h32 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h33 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h34 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h35 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h36 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h37 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h38 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h39 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h3a :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h3b :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h3c :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h3d :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h3e :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h3f :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h40 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h41 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h42 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h43 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h44 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h45 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h46 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h47 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h48 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h49 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h4a :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h4b :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h4c :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h4d :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h4e :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h4f :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h50 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h51 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h52 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h53 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h54 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h55 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h56 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h57 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h58 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h59 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h5a :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h5b :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h5c :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h5d :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h5e :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h5f :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h60 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h61 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h62 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h63 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h64 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h65 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h66 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h67 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h68 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h69 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h6a :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h6b :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h6c :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h6d :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h6e :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h6f :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h70 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h71 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h72 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h73 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h74 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h75 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h76 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h77 :
		RG_quantized_block_rl_57_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h78 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h79 :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h7a :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h7b :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h7c :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h7d :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h7e :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	7'h7f :
		RG_quantized_block_rl_57_t1 = rl_a119_t8 ;
	default :
		RG_quantized_block_rl_57_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_57_t1 or U_318 or TR_146 or U_317 or RG_rl_121 or 
	ST1_07d or RG_rl_119 or U_88 or jpeg_in_a57 or U_01 or RG_quantized_block_rl_59 or 
	ST1_01d )
	RG_quantized_block_rl_57_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_59 )
		| ( { 9{ U_01 } } & jpeg_in_a57 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_119 )
		| ( { 9{ ST1_07d } } & RG_rl_121 )
		| ( { 9{ U_317 } } & TR_146 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_57_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_57_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_57_en )
		RG_quantized_block_rl_57 <= RG_quantized_block_rl_57_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a121_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h01 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h02 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h03 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h04 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h05 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h06 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h07 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h08 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h09 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h0a :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h0b :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h0c :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h0d :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h0e :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h0f :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h10 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h11 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h12 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h13 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h14 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h15 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h16 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h17 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h18 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h19 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h1a :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h1b :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h1c :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h1d :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h1e :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h1f :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h20 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h21 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h22 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h23 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h24 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h25 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h26 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h27 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h28 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h29 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h2a :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h2b :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h2c :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h2d :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h2e :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h2f :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h30 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h31 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h32 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h33 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h34 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h35 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h36 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h37 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h38 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h39 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h3a :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h3b :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h3c :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h3d :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h3e :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h3f :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h40 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h41 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h42 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h43 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h44 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h45 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h46 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h47 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h48 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h49 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h4a :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h4b :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h4c :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h4d :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h4e :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h4f :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h50 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h51 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h52 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h53 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h54 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h55 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h56 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h57 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h58 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h59 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h5a :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h5b :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h5c :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h5d :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h5e :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h5f :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h60 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h61 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h62 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h63 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h64 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h65 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h66 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h67 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h68 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h69 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h6a :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h6b :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h6c :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h6d :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h6e :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h6f :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h70 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h71 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h72 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h73 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h74 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h75 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h76 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h77 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h78 :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h79 :
		RG_quantized_block_rl_58_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h7a :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h7b :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h7c :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h7d :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h7e :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	7'h7f :
		RG_quantized_block_rl_58_t1 = rl_a121_t8 ;
	default :
		RG_quantized_block_rl_58_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_58_t1 or U_318 or TR_144 or U_317 or RG_rl_123 or 
	ST1_07d or RG_rl_121 or U_88 or jpeg_in_a58 or U_01 or RG_quantized_block_rl_60 or 
	ST1_01d )
	RG_quantized_block_rl_58_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_60 )
		| ( { 9{ U_01 } } & jpeg_in_a58 )			// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_121 )
		| ( { 9{ ST1_07d } } & RG_rl_123 )
		| ( { 9{ U_317 } } & TR_144 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_58_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_58_en = ( ST1_01d | U_01 | U_88 | ST1_07d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_58_en )
		RG_quantized_block_rl_58 <= RG_quantized_block_rl_58_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a123_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h01 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h02 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h03 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h04 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h05 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h06 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h07 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h08 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h09 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h0a :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h0b :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h0c :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h0d :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h0e :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h0f :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h10 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h11 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h12 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h13 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h14 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h15 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h16 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h17 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h18 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h19 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h1a :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h1b :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h1c :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h1d :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h1e :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h1f :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h20 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h21 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h22 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h23 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h24 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h25 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h26 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h27 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h28 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h29 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h2a :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h2b :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h2c :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h2d :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h2e :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h2f :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h30 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h31 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h32 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h33 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h34 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h35 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h36 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h37 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h38 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h39 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h3a :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h3b :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h3c :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h3d :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h3e :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h3f :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h40 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h41 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h42 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h43 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h44 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h45 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h46 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h47 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h48 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h49 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h4a :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h4b :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h4c :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h4d :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h4e :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h4f :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h50 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h51 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h52 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h53 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h54 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h55 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h56 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h57 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h58 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h59 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h5a :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h5b :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h5c :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h5d :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h5e :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h5f :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h60 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h61 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h62 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h63 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h64 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h65 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h66 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h67 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h68 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h69 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h6a :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h6b :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h6c :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h6d :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h6e :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h6f :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h70 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h71 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h72 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h73 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h74 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h75 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h76 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h77 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h78 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h79 :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h7a :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h7b :
		RG_quantized_block_rl_59_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h7c :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h7d :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h7e :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	7'h7f :
		RG_quantized_block_rl_59_t1 = rl_a123_t8 ;
	default :
		RG_quantized_block_rl_59_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_59_t1 or U_318 or TR_142 or U_317 or RG_rl_123 or 
	U_88 or jpeg_in_a59 or ST1_02d )
	RG_quantized_block_rl_59_t = ( ( { 9{ ST1_02d } } & jpeg_in_a59 )	// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_123 )
		| ( { 9{ U_317 } } & TR_142 )					// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_59_t1 )		// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_59_en = ( ST1_02d | U_88 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_59_en )
		RG_quantized_block_rl_59 <= RG_quantized_block_rl_59_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a125_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h01 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h02 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h03 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h04 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h05 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h06 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h07 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h08 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h09 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h0a :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h0b :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h0c :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h0d :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h0e :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h0f :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h10 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h11 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h12 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h13 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h14 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h15 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h16 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h17 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h18 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h19 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h1a :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h1b :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h1c :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h1d :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h1e :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h1f :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h20 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h21 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h22 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h23 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h24 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h25 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h26 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h27 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h28 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h29 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h2a :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h2b :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h2c :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h2d :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h2e :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h2f :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h30 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h31 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h32 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h33 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h34 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h35 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h36 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h37 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h38 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h39 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h3a :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h3b :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h3c :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h3d :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h3e :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h3f :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h40 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h41 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h42 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h43 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h44 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h45 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h46 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h47 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h48 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h49 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h4a :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h4b :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h4c :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h4d :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h4e :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h4f :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h50 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h51 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h52 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h53 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h54 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h55 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h56 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h57 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h58 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h59 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h5a :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h5b :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h5c :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h5d :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h5e :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h5f :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h60 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h61 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h62 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h63 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h64 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h65 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h66 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h67 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h68 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h69 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h6a :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h6b :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h6c :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h6d :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h6e :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h6f :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h70 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h71 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h72 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h73 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h74 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h75 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h76 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h77 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h78 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h79 :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h7a :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h7b :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h7c :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h7d :
		RG_quantized_block_rl_60_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h7e :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	7'h7f :
		RG_quantized_block_rl_60_t1 = rl_a125_t8 ;
	default :
		RG_quantized_block_rl_60_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_60_t1 or U_318 or TR_140 or U_317 or RG_rl_125 or 
	U_88 or jpeg_in_a60 or ST1_02d )
	RG_quantized_block_rl_60_t = ( ( { 9{ ST1_02d } } & jpeg_in_a60 )	// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_rl_125 )
		| ( { 9{ U_317 } } & TR_140 )					// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_60_t1 )		// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_60_en = ( ST1_02d | U_88 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_60_en )
		RG_quantized_block_rl_60 <= RG_quantized_block_rl_60_t ;	// line#=../rle.cpp:45,68,69,73,74
always @ ( M_16_t or rl_a126_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h01 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h02 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h03 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h04 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h05 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h06 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h07 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h08 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h09 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h0a :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h0b :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h0c :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h0d :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h0e :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h0f :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h10 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h11 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h12 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h13 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h14 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h15 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h16 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h17 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h18 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h19 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h1a :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h1b :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h1c :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h1d :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h1e :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h1f :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h20 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h21 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h22 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h23 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h24 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h25 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h26 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h27 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h28 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h29 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h2a :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h2b :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h2c :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h2d :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h2e :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h2f :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h30 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h31 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h32 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h33 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h34 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h35 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h36 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h37 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h38 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h39 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h3a :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h3b :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h3c :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h3d :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h3e :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h3f :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h40 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h41 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h42 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h43 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h44 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h45 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h46 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h47 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h48 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h49 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h4a :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h4b :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h4c :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h4d :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h4e :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h4f :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h50 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h51 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h52 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h53 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h54 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h55 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h56 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h57 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h58 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h59 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h5a :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h5b :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h5c :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h5d :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h5e :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h5f :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h60 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h61 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h62 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h63 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h64 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h65 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h66 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h67 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h68 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h69 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h6a :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h6b :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h6c :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h6d :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h6e :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h6f :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h70 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h71 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h72 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h73 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h74 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h75 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h76 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h77 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h78 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h79 :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h7a :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h7b :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h7c :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h7d :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	7'h7e :
		RG_quantized_block_rl_61_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h7f :
		RG_quantized_block_rl_61_t1 = rl_a126_t8 ;
	default :
		RG_quantized_block_rl_61_t1 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_61_t1 or U_318 or TR_139 or U_317 or RG_rl_126 or 
	M_183 or jpeg_in_a61 or U_01 or RG_k_quantized_block_rl_01 or ST1_01d )
	RG_quantized_block_rl_61_t = ( ( { 9{ ST1_01d } } & RG_k_quantized_block_rl_01 )
		| ( { 9{ U_01 } } & jpeg_in_a61 )			// line#=../rle.cpp:45
		| ( { 9{ M_183 } } & RG_rl_126 )
		| ( { 9{ U_317 } } & TR_139 )				// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_quantized_block_rl_61_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_quantized_block_rl_61_en = ( ST1_01d | U_01 | M_183 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_61_en )
		RG_quantized_block_rl_61 <= RG_quantized_block_rl_61_t ;	// line#=../rle.cpp:45,68,69,73,74
assign	M_183 = ( U_88 | ST1_07d ) ;
always @ ( rl_a127_t7 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h01 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h02 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h03 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h04 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h05 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h06 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h07 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h08 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h09 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h0a :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h0b :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h0c :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h0d :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h0e :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h0f :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h10 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h11 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h12 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h13 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h14 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h15 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h16 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h17 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h18 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h19 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h1a :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h1b :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h1c :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h1d :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h1e :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h1f :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h20 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h21 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h22 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h23 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h24 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h25 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h26 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h27 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h28 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h29 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h2a :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h2b :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h2c :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h2d :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h2e :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h2f :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h30 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h31 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h32 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h33 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h34 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h35 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h36 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h37 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h38 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h39 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h3a :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h3b :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h3c :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h3d :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h3e :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h3f :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h40 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h41 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h42 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h43 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h44 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h45 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h46 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h47 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h48 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h49 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h4a :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h4b :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h4c :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h4d :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h4e :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h4f :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h50 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h51 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h52 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h53 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h54 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h55 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h56 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h57 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h58 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h59 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h5a :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h5b :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h5c :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h5d :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h5e :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h5f :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h60 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h61 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h62 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h63 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h64 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h65 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h66 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h67 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h68 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h69 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h6a :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h6b :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h6c :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h6d :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h6e :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h6f :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h70 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h71 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h72 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h73 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h74 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h75 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h76 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h77 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h78 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h79 :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h7a :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h7b :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h7c :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h7d :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h7e :
		RG_k_quantized_block_rl_01_t1 = rl_a127_t7 ;
	7'h7f :
		RG_k_quantized_block_rl_01_t1 = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_k_quantized_block_rl_01_t1 = 9'hx ;
	endcase
always @ ( M_16_t or rl_a127_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h01 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h02 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h03 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h04 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h05 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h06 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h07 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h08 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h09 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h0a :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h0b :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h0c :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h0d :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h0e :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h0f :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h10 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h11 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h12 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h13 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h14 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h15 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h16 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h17 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h18 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h19 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h1a :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h1b :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h1c :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h1d :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h1e :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h1f :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h20 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h21 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h22 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h23 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h24 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h25 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h26 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h27 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h28 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h29 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h2a :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h2b :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h2c :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h2d :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h2e :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h2f :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h30 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h31 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h32 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h33 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h34 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h35 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h36 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h37 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h38 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h39 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h3a :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h3b :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h3c :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h3d :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h3e :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h3f :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h40 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h41 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h42 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h43 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h44 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h45 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h46 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h47 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h48 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h49 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h4a :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h4b :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h4c :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h4d :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h4e :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h4f :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h50 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h51 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h52 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h53 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h54 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h55 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h56 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h57 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h58 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h59 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h5a :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h5b :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h5c :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h5d :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h5e :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h5f :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h60 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h61 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h62 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h63 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h64 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h65 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h66 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h67 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h68 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h69 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h6a :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h6b :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h6c :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h6d :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h6e :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h6f :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h70 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h71 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h72 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h73 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h74 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h75 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h76 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h77 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h78 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h79 :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h7a :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h7b :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h7c :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h7d :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h7e :
		RG_k_quantized_block_rl_01_t2 = rl_a127_t8 ;
	7'h7f :
		RG_k_quantized_block_rl_01_t2 = M_16_t ;	// line#=../rle.cpp:74
	default :
		RG_k_quantized_block_rl_01_t2 = 9'hx ;
	endcase
always @ ( RG_k_quantized_block_rl_01_t2 or U_318 or RG_k_quantized_block_rl_01_t1 or 
	U_317 or RG_i_k_01 or ST1_06d or RG_rl_127 or M_183 or jpeg_in_a62 or U_01 or 
	RG_quantized_block_rl_zz or ST1_01d )
	RG_k_quantized_block_rl_01_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_zz )
		| ( { 9{ U_01 } } & jpeg_in_a62 )			// line#=../rle.cpp:45
		| ( { 9{ M_183 } } & RG_rl_127 )
		| ( { 9{ ST1_06d } } & RG_i_k_01 [8:0] )		// line#=../rle.cpp:61,62
		| ( { 9{ U_317 } } & RG_k_quantized_block_rl_01_t1 )	// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_k_quantized_block_rl_01_t2 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_k_quantized_block_rl_01_en = ( ST1_01d | U_01 | M_183 | ST1_06d | U_317 | 
	U_318 ) ;
always @ ( posedge clk )
	if ( RG_k_quantized_block_rl_01_en )
		RG_k_quantized_block_rl_01 <= RG_k_quantized_block_rl_01_t ;	// line#=../rle.cpp:45,61,62,68,69,73,74
always @ ( RG_rl_125 or U_184 or RG_previous_dc_zz or U_88 or jpeg_in_a63 or U_01 or 
	RG_quantized_block_rl_61 or ST1_01d )
	RG_quantized_block_rl_zz_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_61 )
		| ( { 9{ U_01 } } & jpeg_in_a63 )	// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & RG_previous_dc_zz )
		| ( { 9{ U_184 } } & RG_rl_125 ) ) ;
assign	RG_quantized_block_rl_zz_en = ( ST1_01d | U_01 | U_88 | U_184 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_zz_en )
		RG_quantized_block_rl_zz <= RG_quantized_block_rl_zz_t ;	// line#=../rle.cpp:45
always @ ( incr8u3ot or ST1_03d )
	RG_k_t = ( { 6{ ST1_03d } } & incr8u3ot [5:0] )	// line#=../rle.cpp:111
		 ;	// line#=../rle.cpp:105
always @ ( posedge clk )
	RG_k <= RG_k_t ;	// line#=../rle.cpp:105,111
assign	M_181 = ( ST1_02d | U_06 ) ;
always @ ( U_163 or U_79 or U_161 or U_81 or M_181 )
	begin
	FF_d_t_c1 = ( ( M_181 | U_81 ) | U_161 ) ;	// line#=../rle.cpp:105,120,136,146
	FF_d_t_c2 = ( U_79 | U_163 ) ;	// line#=../rle.cpp:115,151
	FF_d_t = ( { 1{ FF_d_t_c2 } } & 1'h1 )	// line#=../rle.cpp:115,151
		 ;	// line#=../rle.cpp:105,120,136,146
	end
assign	FF_d_en = ( FF_d_t_c1 | FF_d_t_c2 ) ;
always @ ( posedge clk )
	if ( FF_d_en )
		FF_d <= FF_d_t ;	// line#=../rle.cpp:105,115,120,136,146
					// ,151
assign	FF_j_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:36
	if ( FF_j_en )
		FF_j <= 1'h0 ;
assign	FF_i_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:37,39
	if ( FF_i_en )
		FF_i <= 1'h1 ;
always @ ( rl_a00_t8 or M_16_t or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_previous_dc_rl_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h01 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h02 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h03 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h04 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h05 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h06 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h07 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h08 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h09 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h0a :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h0b :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h0c :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h0d :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h0e :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h0f :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h10 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h11 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h12 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h13 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h14 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h15 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h16 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h17 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h18 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h19 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h1a :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h1b :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h1c :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h1d :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h1e :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h1f :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h20 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h21 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h22 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h23 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h24 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h25 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h26 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h27 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h28 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h29 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h2a :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h2b :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h2c :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h2d :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h2e :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h2f :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h30 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h31 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h32 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h33 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h34 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h35 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h36 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h37 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h38 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h39 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h3a :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h3b :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h3c :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h3d :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h3e :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h3f :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h40 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h41 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h42 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h43 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h44 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h45 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h46 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h47 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h48 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h49 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h4a :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h4b :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h4c :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h4d :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h4e :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h4f :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h50 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h51 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h52 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h53 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h54 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h55 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h56 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h57 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h58 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h59 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h5a :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h5b :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h5c :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h5d :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h5e :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h5f :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h60 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h61 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h62 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h63 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h64 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h65 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h66 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h67 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h68 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h69 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h6a :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h6b :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h6c :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h6d :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h6e :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h6f :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h70 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h71 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h72 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h73 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h74 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h75 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h76 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h77 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h78 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h79 :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h7a :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h7b :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h7c :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h7d :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h7e :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	7'h7f :
		RG_previous_dc_rl_t1 = rl_a00_t8 ;
	default :
		RG_previous_dc_rl_t1 = 9'hx ;
	endcase
always @ ( RG_previous_dc_rl_t1 or U_318 or TR_265 or U_317 or RG_previous_dc_zz or 
	ST1_07d or sub12s_91ot or U_88 )
	RG_previous_dc_rl_t = ( ( { 9{ U_88 } } & sub12s_91ot )	// line#=../rle.cpp:52
		| ( { 9{ ST1_07d } } & RG_previous_dc_zz )
		| ( { 9{ U_317 } } & TR_265 )			// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_previous_dc_rl_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_previous_dc_rl_en = ( U_88 | ST1_07d | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( !rst )
		RG_previous_dc_rl <= 9'h000 ;
	else if ( RG_previous_dc_rl_en )
		RG_previous_dc_rl <= RG_previous_dc_rl_t ;	// line#=../rle.cpp:52,68,69,73,74
always @ ( M_16_t or rl_a01_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h01 :
		RG_rl_128_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h02 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h03 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h04 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h05 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h06 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h07 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h08 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h09 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h0a :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h0b :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h0c :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h0d :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h0e :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h0f :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h10 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h11 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h12 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h13 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h14 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h15 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h16 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h17 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h18 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h19 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h1a :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h1b :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h1c :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h1d :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h1e :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h1f :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h20 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h21 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h22 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h23 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h24 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h25 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h26 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h27 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h28 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h29 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h2a :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h2b :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h2c :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h2d :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h2e :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h2f :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h30 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h31 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h32 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h33 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h34 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h35 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h36 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h37 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h38 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h39 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h3a :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h3b :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h3c :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h3d :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h3e :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h3f :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h40 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h41 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h42 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h43 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h44 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h45 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h46 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h47 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h48 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h49 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h4a :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h4b :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h4c :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h4d :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h4e :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h4f :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h50 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h51 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h52 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h53 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h54 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h55 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h56 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h57 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h58 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h59 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h5a :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h5b :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h5c :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h5d :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h5e :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h5f :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h60 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h61 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h62 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h63 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h64 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h65 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h66 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h67 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h68 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h69 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h6a :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h6b :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h6c :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h6d :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h6e :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h6f :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h70 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h71 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h72 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h73 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h74 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h75 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h76 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h77 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h78 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h79 :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h7a :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h7b :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h7c :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h7d :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h7e :
		RG_rl_128_t1 = rl_a01_t8 ;
	7'h7f :
		RG_rl_128_t1 = rl_a01_t8 ;
	default :
		RG_rl_128_t1 = 9'hx ;
	endcase
always @ ( RG_rl_128_t1 or U_318 or TR_264 or U_317 or RG_rl_1 or ST1_03d )
	RG_rl_128_t = ( ( { 9{ ST1_03d } } & RG_rl_1 )
		| ( { 9{ U_317 } } & TR_264 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_128_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_128_en = ( ST1_03d | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_128_en )
		RG_rl_128 <= RG_rl_128_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a02_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h01 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h02 :
		RG_rl_129_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h03 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h04 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h05 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h06 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h07 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h08 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h09 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h0a :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h0b :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h0c :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h0d :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h0e :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h0f :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h10 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h11 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h12 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h13 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h14 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h15 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h16 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h17 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h18 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h19 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h1a :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h1b :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h1c :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h1d :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h1e :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h1f :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h20 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h21 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h22 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h23 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h24 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h25 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h26 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h27 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h28 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h29 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h2a :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h2b :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h2c :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h2d :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h2e :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h2f :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h30 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h31 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h32 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h33 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h34 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h35 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h36 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h37 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h38 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h39 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h3a :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h3b :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h3c :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h3d :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h3e :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h3f :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h40 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h41 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h42 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h43 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h44 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h45 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h46 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h47 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h48 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h49 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h4a :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h4b :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h4c :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h4d :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h4e :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h4f :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h50 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h51 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h52 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h53 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h54 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h55 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h56 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h57 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h58 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h59 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h5a :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h5b :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h5c :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h5d :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h5e :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h5f :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h60 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h61 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h62 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h63 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h64 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h65 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h66 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h67 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h68 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h69 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h6a :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h6b :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h6c :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h6d :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h6e :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h6f :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h70 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h71 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h72 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h73 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h74 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h75 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h76 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h77 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h78 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h79 :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h7a :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h7b :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h7c :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h7d :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h7e :
		RG_rl_129_t1 = rl_a02_t8 ;
	7'h7f :
		RG_rl_129_t1 = rl_a02_t8 ;
	default :
		RG_rl_129_t1 = 9'hx ;
	endcase
always @ ( RG_rl_129_t1 or U_318 or TR_263 or U_317 or RG_rl_2 or ST1_03d )
	RG_rl_129_t = ( ( { 9{ ST1_03d } } & RG_rl_2 )
		| ( { 9{ U_317 } } & TR_263 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_129_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_129_en = ( ST1_03d | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_129_en )
		RG_rl_129 <= RG_rl_129_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a03_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h01 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h02 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h03 :
		RG_rl_130_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h04 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h05 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h06 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h07 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h08 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h09 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h0a :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h0b :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h0c :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h0d :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h0e :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h0f :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h10 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h11 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h12 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h13 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h14 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h15 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h16 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h17 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h18 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h19 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h1a :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h1b :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h1c :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h1d :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h1e :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h1f :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h20 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h21 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h22 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h23 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h24 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h25 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h26 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h27 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h28 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h29 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h2a :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h2b :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h2c :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h2d :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h2e :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h2f :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h30 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h31 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h32 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h33 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h34 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h35 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h36 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h37 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h38 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h39 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h3a :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h3b :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h3c :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h3d :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h3e :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h3f :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h40 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h41 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h42 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h43 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h44 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h45 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h46 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h47 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h48 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h49 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h4a :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h4b :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h4c :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h4d :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h4e :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h4f :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h50 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h51 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h52 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h53 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h54 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h55 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h56 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h57 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h58 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h59 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h5a :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h5b :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h5c :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h5d :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h5e :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h5f :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h60 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h61 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h62 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h63 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h64 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h65 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h66 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h67 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h68 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h69 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h6a :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h6b :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h6c :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h6d :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h6e :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h6f :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h70 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h71 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h72 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h73 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h74 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h75 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h76 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h77 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h78 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h79 :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h7a :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h7b :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h7c :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h7d :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h7e :
		RG_rl_130_t1 = rl_a03_t8 ;
	7'h7f :
		RG_rl_130_t1 = rl_a03_t8 ;
	default :
		RG_rl_130_t1 = 9'hx ;
	endcase
always @ ( RG_rl_130_t1 or U_318 or TR_262 or U_317 or RG_rl_3 or ST1_03d )
	RG_rl_130_t = ( ( { 9{ ST1_03d } } & RG_rl_3 )
		| ( { 9{ U_317 } } & TR_262 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_130_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_130_en = ( ST1_03d | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_130_en )
		RG_rl_130 <= RG_rl_130_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a04_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h01 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h02 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h03 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h04 :
		RG_rl_131_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h05 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h06 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h07 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h08 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h09 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h0a :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h0b :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h0c :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h0d :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h0e :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h0f :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h10 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h11 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h12 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h13 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h14 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h15 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h16 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h17 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h18 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h19 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h1a :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h1b :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h1c :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h1d :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h1e :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h1f :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h20 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h21 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h22 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h23 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h24 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h25 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h26 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h27 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h28 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h29 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h2a :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h2b :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h2c :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h2d :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h2e :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h2f :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h30 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h31 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h32 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h33 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h34 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h35 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h36 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h37 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h38 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h39 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h3a :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h3b :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h3c :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h3d :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h3e :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h3f :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h40 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h41 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h42 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h43 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h44 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h45 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h46 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h47 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h48 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h49 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h4a :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h4b :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h4c :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h4d :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h4e :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h4f :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h50 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h51 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h52 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h53 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h54 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h55 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h56 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h57 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h58 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h59 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h5a :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h5b :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h5c :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h5d :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h5e :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h5f :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h60 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h61 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h62 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h63 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h64 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h65 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h66 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h67 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h68 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h69 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h6a :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h6b :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h6c :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h6d :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h6e :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h6f :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h70 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h71 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h72 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h73 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h74 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h75 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h76 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h77 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h78 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h79 :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h7a :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h7b :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h7c :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h7d :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h7e :
		RG_rl_131_t1 = rl_a04_t8 ;
	7'h7f :
		RG_rl_131_t1 = rl_a04_t8 ;
	default :
		RG_rl_131_t1 = 9'hx ;
	endcase
always @ ( RG_rl_131_t1 or U_318 or TR_261 or U_317 or RG_rl_5 or ST1_07d or RG_rl_4 or 
	U_88 or RG_quantized_block_rl_1 or ST1_01d )
	RG_rl_131_t = ( ( { 9{ ST1_01d } } & RG_quantized_block_rl_1 )
		| ( { 9{ U_88 } } & RG_rl_4 )
		| ( { 9{ ST1_07d } } & RG_rl_5 )
		| ( { 9{ U_317 } } & TR_261 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_131_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_131_en = ( ST1_01d | U_88 | ST1_07d | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_131_en )
		RG_rl_131 <= RG_rl_131_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a06_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h01 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h02 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h03 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h04 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h05 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h06 :
		RG_rl_132_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h07 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h08 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h09 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h0a :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h0b :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h0c :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h0d :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h0e :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h0f :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h10 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h11 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h12 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h13 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h14 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h15 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h16 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h17 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h18 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h19 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h1a :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h1b :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h1c :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h1d :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h1e :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h1f :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h20 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h21 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h22 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h23 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h24 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h25 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h26 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h27 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h28 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h29 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h2a :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h2b :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h2c :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h2d :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h2e :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h2f :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h30 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h31 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h32 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h33 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h34 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h35 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h36 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h37 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h38 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h39 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h3a :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h3b :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h3c :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h3d :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h3e :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h3f :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h40 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h41 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h42 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h43 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h44 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h45 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h46 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h47 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h48 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h49 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h4a :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h4b :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h4c :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h4d :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h4e :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h4f :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h50 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h51 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h52 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h53 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h54 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h55 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h56 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h57 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h58 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h59 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h5a :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h5b :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h5c :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h5d :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h5e :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h5f :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h60 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h61 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h62 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h63 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h64 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h65 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h66 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h67 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h68 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h69 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h6a :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h6b :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h6c :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h6d :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h6e :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h6f :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h70 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h71 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h72 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h73 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h74 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h75 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h76 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h77 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h78 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h79 :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h7a :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h7b :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h7c :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h7d :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h7e :
		RG_rl_132_t1 = rl_a06_t8 ;
	7'h7f :
		RG_rl_132_t1 = rl_a06_t8 ;
	default :
		RG_rl_132_t1 = 9'hx ;
	endcase
always @ ( RG_rl_132_t1 or U_318 or TR_259 or U_317 or RG_rl_6 or U_06 or RG_quantized_block_rl or 
	ST1_02d )
	RG_rl_132_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl )
		| ( { 9{ U_06 } } & RG_rl_6 )
		| ( { 9{ U_317 } } & TR_259 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_132_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_132_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_132_en )
		RG_rl_132 <= RG_rl_132_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a08_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h01 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h02 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h03 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h04 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h05 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h06 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h07 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h08 :
		RG_rl_133_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h09 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h0a :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h0b :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h0c :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h0d :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h0e :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h0f :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h10 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h11 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h12 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h13 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h14 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h15 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h16 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h17 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h18 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h19 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h1a :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h1b :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h1c :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h1d :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h1e :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h1f :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h20 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h21 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h22 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h23 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h24 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h25 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h26 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h27 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h28 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h29 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h2a :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h2b :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h2c :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h2d :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h2e :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h2f :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h30 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h31 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h32 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h33 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h34 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h35 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h36 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h37 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h38 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h39 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h3a :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h3b :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h3c :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h3d :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h3e :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h3f :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h40 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h41 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h42 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h43 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h44 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h45 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h46 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h47 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h48 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h49 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h4a :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h4b :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h4c :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h4d :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h4e :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h4f :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h50 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h51 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h52 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h53 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h54 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h55 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h56 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h57 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h58 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h59 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h5a :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h5b :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h5c :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h5d :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h5e :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h5f :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h60 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h61 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h62 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h63 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h64 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h65 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h66 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h67 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h68 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h69 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h6a :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h6b :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h6c :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h6d :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h6e :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h6f :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h70 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h71 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h72 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h73 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h74 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h75 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h76 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h77 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h78 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h79 :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h7a :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h7b :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h7c :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h7d :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h7e :
		RG_rl_133_t1 = rl_a08_t8 ;
	7'h7f :
		RG_rl_133_t1 = rl_a08_t8 ;
	default :
		RG_rl_133_t1 = 9'hx ;
	endcase
always @ ( RG_rl_133_t1 or U_318 or TR_257 or U_317 or RG_rl_8 or U_06 or RG_quantized_block_rl_1 or 
	ST1_02d )
	RG_rl_133_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_1 )
		| ( { 9{ U_06 } } & RG_rl_8 )
		| ( { 9{ U_317 } } & TR_257 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_133_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_133_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_133_en )
		RG_rl_133 <= RG_rl_133_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a10_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h01 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h02 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h03 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h04 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h05 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h06 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h07 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h08 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h09 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h0a :
		RG_rl_134_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h0b :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h0c :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h0d :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h0e :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h0f :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h10 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h11 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h12 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h13 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h14 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h15 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h16 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h17 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h18 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h19 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h1a :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h1b :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h1c :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h1d :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h1e :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h1f :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h20 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h21 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h22 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h23 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h24 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h25 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h26 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h27 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h28 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h29 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h2a :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h2b :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h2c :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h2d :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h2e :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h2f :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h30 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h31 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h32 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h33 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h34 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h35 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h36 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h37 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h38 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h39 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h3a :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h3b :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h3c :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h3d :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h3e :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h3f :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h40 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h41 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h42 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h43 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h44 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h45 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h46 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h47 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h48 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h49 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h4a :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h4b :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h4c :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h4d :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h4e :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h4f :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h50 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h51 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h52 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h53 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h54 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h55 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h56 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h57 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h58 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h59 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h5a :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h5b :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h5c :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h5d :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h5e :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h5f :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h60 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h61 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h62 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h63 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h64 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h65 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h66 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h67 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h68 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h69 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h6a :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h6b :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h6c :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h6d :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h6e :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h6f :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h70 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h71 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h72 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h73 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h74 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h75 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h76 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h77 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h78 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h79 :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h7a :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h7b :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h7c :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h7d :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h7e :
		RG_rl_134_t1 = rl_a10_t8 ;
	7'h7f :
		RG_rl_134_t1 = rl_a10_t8 ;
	default :
		RG_rl_134_t1 = 9'hx ;
	endcase
always @ ( RG_rl_134_t1 or U_318 or TR_255 or U_317 or RG_rl_10 or U_06 or RG_quantized_block_rl_2 or 
	ST1_02d )
	RG_rl_134_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_2 )
		| ( { 9{ U_06 } } & RG_rl_10 )
		| ( { 9{ U_317 } } & TR_255 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_134_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_134_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_134_en )
		RG_rl_134 <= RG_rl_134_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a12_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h01 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h02 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h03 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h04 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h05 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h06 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h07 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h08 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h09 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h0a :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h0b :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h0c :
		RG_rl_135_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h0d :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h0e :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h0f :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h10 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h11 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h12 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h13 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h14 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h15 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h16 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h17 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h18 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h19 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h1a :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h1b :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h1c :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h1d :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h1e :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h1f :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h20 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h21 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h22 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h23 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h24 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h25 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h26 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h27 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h28 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h29 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h2a :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h2b :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h2c :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h2d :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h2e :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h2f :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h30 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h31 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h32 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h33 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h34 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h35 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h36 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h37 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h38 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h39 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h3a :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h3b :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h3c :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h3d :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h3e :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h3f :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h40 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h41 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h42 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h43 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h44 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h45 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h46 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h47 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h48 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h49 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h4a :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h4b :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h4c :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h4d :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h4e :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h4f :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h50 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h51 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h52 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h53 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h54 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h55 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h56 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h57 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h58 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h59 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h5a :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h5b :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h5c :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h5d :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h5e :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h5f :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h60 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h61 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h62 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h63 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h64 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h65 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h66 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h67 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h68 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h69 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h6a :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h6b :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h6c :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h6d :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h6e :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h6f :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h70 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h71 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h72 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h73 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h74 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h75 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h76 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h77 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h78 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h79 :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h7a :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h7b :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h7c :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h7d :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h7e :
		RG_rl_135_t1 = rl_a12_t8 ;
	7'h7f :
		RG_rl_135_t1 = rl_a12_t8 ;
	default :
		RG_rl_135_t1 = 9'hx ;
	endcase
always @ ( RG_rl_135_t1 or U_318 or TR_253 or U_317 or RG_rl_12 or U_06 or RG_quantized_block_rl_3 or 
	ST1_02d )
	RG_rl_135_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_3 )
		| ( { 9{ U_06 } } & RG_rl_12 )
		| ( { 9{ U_317 } } & TR_253 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_135_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_135_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_135_en )
		RG_rl_135 <= RG_rl_135_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a14_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h01 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h02 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h03 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h04 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h05 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h06 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h07 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h08 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h09 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h0a :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h0b :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h0c :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h0d :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h0e :
		RG_rl_136_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h0f :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h10 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h11 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h12 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h13 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h14 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h15 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h16 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h17 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h18 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h19 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h1a :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h1b :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h1c :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h1d :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h1e :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h1f :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h20 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h21 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h22 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h23 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h24 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h25 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h26 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h27 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h28 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h29 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h2a :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h2b :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h2c :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h2d :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h2e :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h2f :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h30 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h31 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h32 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h33 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h34 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h35 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h36 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h37 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h38 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h39 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h3a :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h3b :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h3c :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h3d :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h3e :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h3f :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h40 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h41 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h42 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h43 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h44 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h45 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h46 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h47 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h48 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h49 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h4a :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h4b :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h4c :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h4d :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h4e :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h4f :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h50 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h51 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h52 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h53 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h54 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h55 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h56 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h57 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h58 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h59 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h5a :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h5b :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h5c :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h5d :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h5e :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h5f :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h60 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h61 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h62 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h63 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h64 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h65 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h66 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h67 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h68 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h69 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h6a :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h6b :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h6c :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h6d :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h6e :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h6f :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h70 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h71 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h72 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h73 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h74 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h75 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h76 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h77 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h78 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h79 :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h7a :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h7b :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h7c :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h7d :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h7e :
		RG_rl_136_t1 = rl_a14_t8 ;
	7'h7f :
		RG_rl_136_t1 = rl_a14_t8 ;
	default :
		RG_rl_136_t1 = 9'hx ;
	endcase
always @ ( RG_rl_136_t1 or U_318 or TR_251 or U_317 or RG_rl_14 or U_06 or RG_quantized_block_rl_4 or 
	ST1_02d )
	RG_rl_136_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_4 )
		| ( { 9{ U_06 } } & RG_rl_14 )
		| ( { 9{ U_317 } } & TR_251 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_136_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_136_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_136_en )
		RG_rl_136 <= RG_rl_136_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a16_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h01 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h02 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h03 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h04 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h05 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h06 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h07 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h08 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h09 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h0a :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h0b :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h0c :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h0d :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h0e :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h0f :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h10 :
		RG_rl_137_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h11 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h12 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h13 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h14 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h15 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h16 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h17 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h18 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h19 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h1a :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h1b :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h1c :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h1d :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h1e :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h1f :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h20 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h21 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h22 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h23 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h24 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h25 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h26 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h27 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h28 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h29 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h2a :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h2b :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h2c :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h2d :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h2e :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h2f :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h30 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h31 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h32 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h33 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h34 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h35 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h36 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h37 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h38 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h39 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h3a :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h3b :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h3c :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h3d :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h3e :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h3f :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h40 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h41 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h42 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h43 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h44 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h45 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h46 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h47 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h48 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h49 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h4a :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h4b :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h4c :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h4d :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h4e :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h4f :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h50 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h51 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h52 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h53 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h54 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h55 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h56 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h57 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h58 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h59 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h5a :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h5b :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h5c :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h5d :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h5e :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h5f :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h60 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h61 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h62 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h63 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h64 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h65 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h66 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h67 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h68 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h69 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h6a :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h6b :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h6c :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h6d :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h6e :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h6f :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h70 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h71 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h72 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h73 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h74 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h75 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h76 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h77 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h78 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h79 :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h7a :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h7b :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h7c :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h7d :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h7e :
		RG_rl_137_t1 = rl_a16_t8 ;
	7'h7f :
		RG_rl_137_t1 = rl_a16_t8 ;
	default :
		RG_rl_137_t1 = 9'hx ;
	endcase
always @ ( RG_rl_137_t1 or U_318 or TR_249 or U_317 or RG_rl_16 or U_06 or RG_quantized_block_rl_5 or 
	ST1_02d )
	RG_rl_137_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_5 )
		| ( { 9{ U_06 } } & RG_rl_16 )
		| ( { 9{ U_317 } } & TR_249 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_137_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_137_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_137_en )
		RG_rl_137 <= RG_rl_137_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a18_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h01 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h02 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h03 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h04 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h05 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h06 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h07 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h08 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h09 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h0a :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h0b :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h0c :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h0d :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h0e :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h0f :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h10 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h11 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h12 :
		RG_rl_138_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h13 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h14 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h15 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h16 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h17 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h18 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h19 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h1a :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h1b :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h1c :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h1d :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h1e :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h1f :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h20 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h21 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h22 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h23 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h24 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h25 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h26 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h27 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h28 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h29 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h2a :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h2b :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h2c :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h2d :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h2e :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h2f :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h30 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h31 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h32 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h33 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h34 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h35 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h36 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h37 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h38 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h39 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h3a :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h3b :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h3c :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h3d :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h3e :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h3f :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h40 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h41 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h42 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h43 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h44 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h45 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h46 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h47 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h48 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h49 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h4a :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h4b :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h4c :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h4d :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h4e :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h4f :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h50 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h51 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h52 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h53 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h54 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h55 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h56 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h57 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h58 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h59 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h5a :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h5b :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h5c :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h5d :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h5e :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h5f :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h60 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h61 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h62 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h63 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h64 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h65 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h66 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h67 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h68 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h69 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h6a :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h6b :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h6c :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h6d :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h6e :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h6f :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h70 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h71 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h72 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h73 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h74 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h75 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h76 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h77 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h78 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h79 :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h7a :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h7b :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h7c :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h7d :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h7e :
		RG_rl_138_t1 = rl_a18_t8 ;
	7'h7f :
		RG_rl_138_t1 = rl_a18_t8 ;
	default :
		RG_rl_138_t1 = 9'hx ;
	endcase
always @ ( RG_rl_138_t1 or U_318 or TR_247 or U_317 or RG_rl_18 or U_06 or RG_quantized_block_rl_6 or 
	ST1_02d )
	RG_rl_138_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_6 )
		| ( { 9{ U_06 } } & RG_rl_18 )
		| ( { 9{ U_317 } } & TR_247 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_138_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_138_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_138_en )
		RG_rl_138 <= RG_rl_138_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a20_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h01 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h02 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h03 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h04 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h05 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h06 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h07 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h08 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h09 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h0a :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h0b :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h0c :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h0d :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h0e :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h0f :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h10 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h11 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h12 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h13 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h14 :
		RG_rl_139_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h15 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h16 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h17 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h18 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h19 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h1a :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h1b :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h1c :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h1d :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h1e :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h1f :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h20 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h21 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h22 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h23 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h24 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h25 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h26 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h27 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h28 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h29 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h2a :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h2b :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h2c :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h2d :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h2e :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h2f :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h30 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h31 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h32 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h33 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h34 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h35 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h36 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h37 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h38 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h39 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h3a :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h3b :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h3c :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h3d :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h3e :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h3f :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h40 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h41 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h42 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h43 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h44 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h45 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h46 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h47 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h48 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h49 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h4a :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h4b :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h4c :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h4d :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h4e :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h4f :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h50 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h51 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h52 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h53 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h54 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h55 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h56 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h57 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h58 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h59 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h5a :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h5b :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h5c :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h5d :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h5e :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h5f :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h60 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h61 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h62 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h63 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h64 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h65 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h66 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h67 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h68 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h69 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h6a :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h6b :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h6c :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h6d :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h6e :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h6f :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h70 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h71 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h72 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h73 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h74 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h75 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h76 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h77 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h78 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h79 :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h7a :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h7b :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h7c :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h7d :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h7e :
		RG_rl_139_t1 = rl_a20_t8 ;
	7'h7f :
		RG_rl_139_t1 = rl_a20_t8 ;
	default :
		RG_rl_139_t1 = 9'hx ;
	endcase
always @ ( RG_rl_139_t1 or U_318 or TR_245 or U_317 or RG_rl_20 or U_06 or RG_quantized_block_rl_7 or 
	ST1_02d )
	RG_rl_139_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_7 )
		| ( { 9{ U_06 } } & RG_rl_20 )
		| ( { 9{ U_317 } } & TR_245 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_139_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_139_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_139_en )
		RG_rl_139 <= RG_rl_139_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a22_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h01 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h02 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h03 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h04 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h05 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h06 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h07 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h08 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h09 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h0a :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h0b :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h0c :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h0d :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h0e :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h0f :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h10 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h11 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h12 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h13 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h14 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h15 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h16 :
		RG_rl_140_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h17 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h18 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h19 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h1a :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h1b :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h1c :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h1d :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h1e :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h1f :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h20 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h21 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h22 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h23 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h24 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h25 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h26 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h27 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h28 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h29 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h2a :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h2b :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h2c :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h2d :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h2e :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h2f :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h30 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h31 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h32 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h33 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h34 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h35 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h36 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h37 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h38 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h39 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h3a :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h3b :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h3c :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h3d :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h3e :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h3f :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h40 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h41 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h42 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h43 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h44 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h45 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h46 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h47 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h48 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h49 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h4a :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h4b :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h4c :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h4d :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h4e :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h4f :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h50 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h51 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h52 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h53 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h54 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h55 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h56 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h57 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h58 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h59 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h5a :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h5b :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h5c :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h5d :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h5e :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h5f :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h60 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h61 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h62 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h63 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h64 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h65 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h66 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h67 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h68 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h69 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h6a :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h6b :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h6c :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h6d :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h6e :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h6f :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h70 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h71 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h72 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h73 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h74 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h75 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h76 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h77 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h78 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h79 :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h7a :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h7b :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h7c :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h7d :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h7e :
		RG_rl_140_t1 = rl_a22_t8 ;
	7'h7f :
		RG_rl_140_t1 = rl_a22_t8 ;
	default :
		RG_rl_140_t1 = 9'hx ;
	endcase
always @ ( RG_rl_140_t1 or U_318 or TR_243 or U_317 or RG_rl_22 or U_06 or RG_quantized_block_rl_8 or 
	ST1_02d )
	RG_rl_140_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_8 )
		| ( { 9{ U_06 } } & RG_rl_22 )
		| ( { 9{ U_317 } } & TR_243 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_140_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_140_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_140_en )
		RG_rl_140 <= RG_rl_140_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a24_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h01 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h02 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h03 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h04 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h05 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h06 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h07 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h08 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h09 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h0a :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h0b :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h0c :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h0d :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h0e :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h0f :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h10 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h11 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h12 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h13 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h14 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h15 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h16 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h17 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h18 :
		RG_rl_141_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h19 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h1a :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h1b :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h1c :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h1d :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h1e :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h1f :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h20 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h21 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h22 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h23 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h24 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h25 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h26 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h27 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h28 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h29 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h2a :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h2b :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h2c :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h2d :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h2e :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h2f :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h30 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h31 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h32 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h33 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h34 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h35 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h36 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h37 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h38 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h39 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h3a :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h3b :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h3c :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h3d :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h3e :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h3f :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h40 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h41 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h42 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h43 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h44 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h45 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h46 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h47 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h48 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h49 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h4a :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h4b :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h4c :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h4d :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h4e :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h4f :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h50 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h51 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h52 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h53 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h54 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h55 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h56 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h57 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h58 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h59 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h5a :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h5b :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h5c :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h5d :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h5e :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h5f :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h60 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h61 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h62 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h63 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h64 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h65 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h66 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h67 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h68 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h69 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h6a :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h6b :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h6c :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h6d :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h6e :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h6f :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h70 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h71 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h72 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h73 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h74 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h75 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h76 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h77 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h78 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h79 :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h7a :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h7b :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h7c :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h7d :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h7e :
		RG_rl_141_t1 = rl_a24_t8 ;
	7'h7f :
		RG_rl_141_t1 = rl_a24_t8 ;
	default :
		RG_rl_141_t1 = 9'hx ;
	endcase
always @ ( RG_rl_141_t1 or U_318 or TR_241 or U_317 or RG_rl_24 or U_06 or RG_quantized_block_rl_9 or 
	ST1_02d )
	RG_rl_141_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_9 )
		| ( { 9{ U_06 } } & RG_rl_24 )
		| ( { 9{ U_317 } } & TR_241 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_141_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_141_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_141_en )
		RG_rl_141 <= RG_rl_141_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a26_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h01 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h02 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h03 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h04 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h05 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h06 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h07 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h08 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h09 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h0a :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h0b :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h0c :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h0d :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h0e :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h0f :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h10 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h11 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h12 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h13 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h14 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h15 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h16 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h17 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h18 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h19 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h1a :
		RG_rl_142_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h1b :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h1c :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h1d :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h1e :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h1f :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h20 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h21 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h22 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h23 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h24 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h25 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h26 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h27 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h28 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h29 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h2a :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h2b :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h2c :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h2d :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h2e :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h2f :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h30 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h31 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h32 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h33 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h34 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h35 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h36 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h37 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h38 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h39 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h3a :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h3b :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h3c :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h3d :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h3e :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h3f :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h40 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h41 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h42 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h43 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h44 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h45 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h46 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h47 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h48 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h49 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h4a :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h4b :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h4c :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h4d :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h4e :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h4f :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h50 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h51 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h52 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h53 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h54 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h55 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h56 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h57 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h58 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h59 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h5a :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h5b :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h5c :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h5d :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h5e :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h5f :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h60 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h61 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h62 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h63 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h64 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h65 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h66 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h67 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h68 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h69 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h6a :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h6b :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h6c :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h6d :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h6e :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h6f :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h70 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h71 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h72 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h73 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h74 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h75 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h76 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h77 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h78 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h79 :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h7a :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h7b :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h7c :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h7d :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h7e :
		RG_rl_142_t1 = rl_a26_t8 ;
	7'h7f :
		RG_rl_142_t1 = rl_a26_t8 ;
	default :
		RG_rl_142_t1 = 9'hx ;
	endcase
always @ ( RG_rl_142_t1 or U_318 or TR_239 or U_317 or RG_rl_26 or U_06 or RG_quantized_block_rl_10 or 
	ST1_02d )
	RG_rl_142_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_10 )
		| ( { 9{ U_06 } } & RG_rl_26 )
		| ( { 9{ U_317 } } & TR_239 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_142_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_142_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_142_en )
		RG_rl_142 <= RG_rl_142_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a28_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h01 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h02 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h03 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h04 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h05 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h06 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h07 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h08 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h09 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h0a :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h0b :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h0c :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h0d :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h0e :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h0f :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h10 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h11 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h12 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h13 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h14 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h15 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h16 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h17 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h18 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h19 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h1a :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h1b :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h1c :
		RG_rl_143_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h1d :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h1e :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h1f :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h20 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h21 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h22 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h23 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h24 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h25 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h26 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h27 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h28 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h29 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h2a :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h2b :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h2c :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h2d :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h2e :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h2f :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h30 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h31 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h32 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h33 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h34 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h35 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h36 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h37 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h38 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h39 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h3a :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h3b :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h3c :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h3d :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h3e :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h3f :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h40 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h41 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h42 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h43 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h44 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h45 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h46 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h47 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h48 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h49 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h4a :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h4b :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h4c :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h4d :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h4e :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h4f :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h50 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h51 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h52 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h53 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h54 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h55 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h56 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h57 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h58 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h59 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h5a :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h5b :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h5c :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h5d :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h5e :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h5f :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h60 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h61 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h62 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h63 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h64 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h65 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h66 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h67 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h68 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h69 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h6a :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h6b :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h6c :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h6d :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h6e :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h6f :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h70 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h71 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h72 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h73 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h74 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h75 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h76 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h77 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h78 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h79 :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h7a :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h7b :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h7c :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h7d :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h7e :
		RG_rl_143_t1 = rl_a28_t8 ;
	7'h7f :
		RG_rl_143_t1 = rl_a28_t8 ;
	default :
		RG_rl_143_t1 = 9'hx ;
	endcase
always @ ( RG_rl_143_t1 or U_318 or TR_237 or U_317 or RG_rl_28 or U_06 or RG_quantized_block_rl_11 or 
	ST1_02d )
	RG_rl_143_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_11 )
		| ( { 9{ U_06 } } & RG_rl_28 )
		| ( { 9{ U_317 } } & TR_237 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_143_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_143_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_143_en )
		RG_rl_143 <= RG_rl_143_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a30_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h01 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h02 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h03 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h04 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h05 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h06 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h07 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h08 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h09 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h0a :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h0b :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h0c :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h0d :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h0e :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h0f :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h10 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h11 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h12 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h13 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h14 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h15 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h16 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h17 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h18 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h19 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h1a :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h1b :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h1c :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h1d :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h1e :
		RG_rl_144_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h1f :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h20 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h21 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h22 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h23 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h24 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h25 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h26 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h27 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h28 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h29 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h2a :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h2b :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h2c :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h2d :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h2e :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h2f :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h30 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h31 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h32 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h33 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h34 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h35 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h36 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h37 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h38 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h39 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h3a :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h3b :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h3c :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h3d :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h3e :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h3f :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h40 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h41 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h42 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h43 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h44 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h45 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h46 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h47 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h48 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h49 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h4a :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h4b :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h4c :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h4d :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h4e :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h4f :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h50 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h51 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h52 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h53 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h54 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h55 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h56 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h57 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h58 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h59 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h5a :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h5b :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h5c :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h5d :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h5e :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h5f :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h60 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h61 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h62 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h63 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h64 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h65 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h66 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h67 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h68 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h69 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h6a :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h6b :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h6c :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h6d :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h6e :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h6f :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h70 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h71 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h72 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h73 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h74 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h75 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h76 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h77 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h78 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h79 :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h7a :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h7b :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h7c :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h7d :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h7e :
		RG_rl_144_t1 = rl_a30_t8 ;
	7'h7f :
		RG_rl_144_t1 = rl_a30_t8 ;
	default :
		RG_rl_144_t1 = 9'hx ;
	endcase
always @ ( RG_rl_144_t1 or U_318 or TR_235 or U_317 or RG_rl_30 or U_06 or RG_quantized_block_rl_12 or 
	ST1_02d )
	RG_rl_144_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_12 )
		| ( { 9{ U_06 } } & RG_rl_30 )
		| ( { 9{ U_317 } } & TR_235 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_144_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_144_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_144_en )
		RG_rl_144 <= RG_rl_144_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a32_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h01 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h02 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h03 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h04 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h05 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h06 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h07 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h08 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h09 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h0a :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h0b :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h0c :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h0d :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h0e :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h0f :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h10 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h11 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h12 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h13 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h14 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h15 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h16 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h17 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h18 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h19 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h1a :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h1b :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h1c :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h1d :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h1e :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h1f :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h20 :
		RG_rl_145_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h21 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h22 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h23 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h24 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h25 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h26 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h27 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h28 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h29 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h2a :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h2b :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h2c :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h2d :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h2e :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h2f :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h30 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h31 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h32 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h33 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h34 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h35 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h36 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h37 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h38 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h39 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h3a :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h3b :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h3c :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h3d :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h3e :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h3f :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h40 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h41 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h42 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h43 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h44 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h45 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h46 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h47 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h48 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h49 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h4a :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h4b :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h4c :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h4d :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h4e :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h4f :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h50 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h51 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h52 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h53 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h54 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h55 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h56 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h57 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h58 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h59 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h5a :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h5b :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h5c :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h5d :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h5e :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h5f :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h60 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h61 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h62 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h63 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h64 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h65 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h66 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h67 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h68 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h69 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h6a :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h6b :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h6c :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h6d :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h6e :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h6f :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h70 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h71 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h72 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h73 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h74 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h75 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h76 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h77 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h78 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h79 :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h7a :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h7b :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h7c :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h7d :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h7e :
		RG_rl_145_t1 = rl_a32_t8 ;
	7'h7f :
		RG_rl_145_t1 = rl_a32_t8 ;
	default :
		RG_rl_145_t1 = 9'hx ;
	endcase
always @ ( RG_rl_145_t1 or U_318 or TR_233 or U_317 or RG_rl_32 or U_06 or RG_quantized_block_rl_13 or 
	ST1_02d )
	RG_rl_145_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_13 )
		| ( { 9{ U_06 } } & RG_rl_32 )
		| ( { 9{ U_317 } } & TR_233 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_145_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_145_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_145_en )
		RG_rl_145 <= RG_rl_145_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a34_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h01 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h02 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h03 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h04 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h05 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h06 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h07 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h08 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h09 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h0a :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h0b :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h0c :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h0d :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h0e :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h0f :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h10 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h11 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h12 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h13 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h14 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h15 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h16 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h17 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h18 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h19 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h1a :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h1b :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h1c :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h1d :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h1e :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h1f :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h20 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h21 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h22 :
		RG_rl_146_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h23 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h24 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h25 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h26 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h27 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h28 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h29 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h2a :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h2b :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h2c :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h2d :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h2e :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h2f :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h30 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h31 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h32 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h33 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h34 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h35 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h36 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h37 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h38 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h39 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h3a :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h3b :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h3c :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h3d :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h3e :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h3f :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h40 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h41 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h42 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h43 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h44 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h45 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h46 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h47 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h48 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h49 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h4a :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h4b :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h4c :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h4d :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h4e :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h4f :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h50 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h51 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h52 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h53 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h54 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h55 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h56 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h57 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h58 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h59 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h5a :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h5b :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h5c :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h5d :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h5e :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h5f :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h60 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h61 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h62 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h63 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h64 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h65 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h66 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h67 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h68 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h69 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h6a :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h6b :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h6c :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h6d :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h6e :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h6f :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h70 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h71 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h72 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h73 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h74 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h75 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h76 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h77 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h78 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h79 :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h7a :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h7b :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h7c :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h7d :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h7e :
		RG_rl_146_t1 = rl_a34_t8 ;
	7'h7f :
		RG_rl_146_t1 = rl_a34_t8 ;
	default :
		RG_rl_146_t1 = 9'hx ;
	endcase
always @ ( RG_rl_146_t1 or U_318 or TR_231 or U_317 or RG_rl_34 or U_06 or RG_quantized_block_rl_14 or 
	ST1_02d )
	RG_rl_146_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_14 )
		| ( { 9{ U_06 } } & RG_rl_34 )
		| ( { 9{ U_317 } } & TR_231 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_146_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_146_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_146_en )
		RG_rl_146 <= RG_rl_146_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a36_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h01 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h02 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h03 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h04 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h05 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h06 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h07 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h08 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h09 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h0a :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h0b :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h0c :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h0d :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h0e :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h0f :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h10 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h11 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h12 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h13 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h14 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h15 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h16 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h17 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h18 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h19 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h1a :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h1b :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h1c :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h1d :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h1e :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h1f :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h20 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h21 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h22 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h23 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h24 :
		RG_rl_147_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h25 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h26 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h27 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h28 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h29 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h2a :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h2b :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h2c :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h2d :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h2e :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h2f :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h30 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h31 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h32 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h33 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h34 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h35 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h36 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h37 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h38 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h39 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h3a :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h3b :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h3c :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h3d :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h3e :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h3f :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h40 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h41 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h42 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h43 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h44 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h45 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h46 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h47 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h48 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h49 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h4a :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h4b :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h4c :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h4d :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h4e :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h4f :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h50 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h51 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h52 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h53 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h54 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h55 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h56 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h57 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h58 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h59 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h5a :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h5b :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h5c :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h5d :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h5e :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h5f :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h60 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h61 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h62 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h63 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h64 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h65 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h66 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h67 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h68 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h69 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h6a :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h6b :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h6c :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h6d :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h6e :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h6f :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h70 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h71 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h72 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h73 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h74 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h75 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h76 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h77 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h78 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h79 :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h7a :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h7b :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h7c :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h7d :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h7e :
		RG_rl_147_t1 = rl_a36_t8 ;
	7'h7f :
		RG_rl_147_t1 = rl_a36_t8 ;
	default :
		RG_rl_147_t1 = 9'hx ;
	endcase
always @ ( RG_rl_147_t1 or U_318 or TR_229 or U_317 or RG_rl_36 or U_06 or RG_quantized_block_rl_15 or 
	ST1_02d )
	RG_rl_147_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_15 )
		| ( { 9{ U_06 } } & RG_rl_36 )
		| ( { 9{ U_317 } } & TR_229 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_147_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_147_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_147_en )
		RG_rl_147 <= RG_rl_147_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a38_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h01 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h02 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h03 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h04 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h05 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h06 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h07 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h08 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h09 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h0a :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h0b :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h0c :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h0d :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h0e :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h0f :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h10 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h11 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h12 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h13 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h14 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h15 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h16 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h17 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h18 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h19 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h1a :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h1b :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h1c :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h1d :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h1e :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h1f :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h20 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h21 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h22 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h23 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h24 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h25 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h26 :
		RG_rl_148_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h27 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h28 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h29 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h2a :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h2b :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h2c :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h2d :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h2e :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h2f :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h30 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h31 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h32 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h33 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h34 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h35 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h36 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h37 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h38 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h39 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h3a :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h3b :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h3c :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h3d :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h3e :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h3f :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h40 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h41 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h42 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h43 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h44 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h45 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h46 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h47 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h48 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h49 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h4a :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h4b :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h4c :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h4d :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h4e :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h4f :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h50 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h51 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h52 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h53 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h54 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h55 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h56 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h57 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h58 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h59 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h5a :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h5b :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h5c :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h5d :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h5e :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h5f :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h60 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h61 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h62 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h63 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h64 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h65 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h66 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h67 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h68 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h69 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h6a :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h6b :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h6c :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h6d :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h6e :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h6f :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h70 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h71 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h72 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h73 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h74 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h75 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h76 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h77 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h78 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h79 :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h7a :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h7b :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h7c :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h7d :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h7e :
		RG_rl_148_t1 = rl_a38_t8 ;
	7'h7f :
		RG_rl_148_t1 = rl_a38_t8 ;
	default :
		RG_rl_148_t1 = 9'hx ;
	endcase
always @ ( RG_rl_148_t1 or U_318 or TR_227 or U_317 or RG_rl_38 or U_06 or RG_quantized_block_rl_16 or 
	ST1_02d )
	RG_rl_148_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_16 )
		| ( { 9{ U_06 } } & RG_rl_38 )
		| ( { 9{ U_317 } } & TR_227 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_148_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_148_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_148_en )
		RG_rl_148 <= RG_rl_148_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a40_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h01 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h02 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h03 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h04 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h05 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h06 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h07 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h08 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h09 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h0a :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h0b :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h0c :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h0d :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h0e :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h0f :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h10 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h11 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h12 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h13 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h14 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h15 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h16 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h17 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h18 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h19 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h1a :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h1b :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h1c :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h1d :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h1e :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h1f :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h20 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h21 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h22 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h23 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h24 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h25 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h26 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h27 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h28 :
		RG_rl_149_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h29 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h2a :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h2b :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h2c :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h2d :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h2e :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h2f :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h30 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h31 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h32 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h33 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h34 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h35 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h36 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h37 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h38 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h39 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h3a :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h3b :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h3c :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h3d :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h3e :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h3f :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h40 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h41 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h42 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h43 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h44 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h45 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h46 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h47 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h48 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h49 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h4a :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h4b :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h4c :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h4d :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h4e :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h4f :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h50 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h51 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h52 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h53 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h54 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h55 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h56 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h57 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h58 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h59 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h5a :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h5b :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h5c :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h5d :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h5e :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h5f :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h60 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h61 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h62 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h63 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h64 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h65 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h66 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h67 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h68 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h69 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h6a :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h6b :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h6c :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h6d :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h6e :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h6f :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h70 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h71 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h72 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h73 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h74 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h75 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h76 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h77 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h78 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h79 :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h7a :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h7b :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h7c :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h7d :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h7e :
		RG_rl_149_t1 = rl_a40_t8 ;
	7'h7f :
		RG_rl_149_t1 = rl_a40_t8 ;
	default :
		RG_rl_149_t1 = 9'hx ;
	endcase
always @ ( RG_rl_149_t1 or U_318 or TR_225 or U_317 or RG_rl_40 or U_06 or RG_quantized_block_rl_17 or 
	ST1_02d )
	RG_rl_149_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_17 )
		| ( { 9{ U_06 } } & RG_rl_40 )
		| ( { 9{ U_317 } } & TR_225 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_149_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_149_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_149_en )
		RG_rl_149 <= RG_rl_149_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a42_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h01 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h02 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h03 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h04 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h05 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h06 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h07 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h08 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h09 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h0a :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h0b :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h0c :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h0d :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h0e :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h0f :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h10 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h11 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h12 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h13 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h14 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h15 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h16 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h17 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h18 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h19 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h1a :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h1b :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h1c :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h1d :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h1e :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h1f :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h20 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h21 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h22 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h23 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h24 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h25 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h26 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h27 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h28 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h29 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h2a :
		RG_rl_150_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h2b :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h2c :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h2d :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h2e :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h2f :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h30 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h31 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h32 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h33 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h34 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h35 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h36 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h37 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h38 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h39 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h3a :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h3b :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h3c :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h3d :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h3e :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h3f :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h40 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h41 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h42 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h43 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h44 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h45 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h46 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h47 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h48 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h49 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h4a :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h4b :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h4c :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h4d :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h4e :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h4f :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h50 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h51 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h52 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h53 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h54 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h55 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h56 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h57 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h58 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h59 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h5a :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h5b :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h5c :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h5d :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h5e :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h5f :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h60 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h61 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h62 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h63 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h64 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h65 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h66 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h67 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h68 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h69 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h6a :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h6b :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h6c :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h6d :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h6e :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h6f :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h70 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h71 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h72 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h73 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h74 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h75 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h76 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h77 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h78 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h79 :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h7a :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h7b :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h7c :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h7d :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h7e :
		RG_rl_150_t1 = rl_a42_t8 ;
	7'h7f :
		RG_rl_150_t1 = rl_a42_t8 ;
	default :
		RG_rl_150_t1 = 9'hx ;
	endcase
always @ ( RG_rl_150_t1 or U_318 or TR_223 or U_317 or RG_rl_42 or U_06 or RG_quantized_block_rl_18 or 
	ST1_02d )
	RG_rl_150_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_18 )
		| ( { 9{ U_06 } } & RG_rl_42 )
		| ( { 9{ U_317 } } & TR_223 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_150_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_150_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_150_en )
		RG_rl_150 <= RG_rl_150_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a44_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h01 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h02 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h03 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h04 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h05 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h06 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h07 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h08 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h09 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h0a :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h0b :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h0c :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h0d :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h0e :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h0f :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h10 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h11 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h12 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h13 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h14 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h15 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h16 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h17 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h18 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h19 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h1a :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h1b :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h1c :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h1d :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h1e :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h1f :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h20 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h21 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h22 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h23 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h24 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h25 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h26 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h27 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h28 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h29 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h2a :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h2b :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h2c :
		RG_rl_151_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h2d :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h2e :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h2f :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h30 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h31 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h32 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h33 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h34 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h35 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h36 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h37 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h38 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h39 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h3a :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h3b :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h3c :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h3d :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h3e :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h3f :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h40 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h41 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h42 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h43 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h44 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h45 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h46 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h47 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h48 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h49 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h4a :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h4b :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h4c :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h4d :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h4e :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h4f :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h50 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h51 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h52 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h53 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h54 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h55 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h56 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h57 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h58 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h59 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h5a :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h5b :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h5c :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h5d :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h5e :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h5f :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h60 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h61 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h62 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h63 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h64 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h65 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h66 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h67 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h68 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h69 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h6a :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h6b :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h6c :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h6d :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h6e :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h6f :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h70 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h71 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h72 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h73 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h74 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h75 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h76 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h77 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h78 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h79 :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h7a :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h7b :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h7c :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h7d :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h7e :
		RG_rl_151_t1 = rl_a44_t8 ;
	7'h7f :
		RG_rl_151_t1 = rl_a44_t8 ;
	default :
		RG_rl_151_t1 = 9'hx ;
	endcase
always @ ( RG_rl_151_t1 or U_318 or TR_221 or U_317 or RG_rl_44 or U_06 or RG_quantized_block_rl_19 or 
	ST1_02d )
	RG_rl_151_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_19 )
		| ( { 9{ U_06 } } & RG_rl_44 )
		| ( { 9{ U_317 } } & TR_221 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_151_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_151_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_151_en )
		RG_rl_151 <= RG_rl_151_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a46_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h01 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h02 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h03 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h04 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h05 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h06 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h07 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h08 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h09 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h0a :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h0b :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h0c :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h0d :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h0e :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h0f :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h10 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h11 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h12 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h13 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h14 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h15 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h16 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h17 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h18 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h19 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h1a :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h1b :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h1c :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h1d :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h1e :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h1f :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h20 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h21 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h22 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h23 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h24 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h25 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h26 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h27 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h28 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h29 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h2a :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h2b :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h2c :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h2d :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h2e :
		RG_rl_152_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h2f :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h30 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h31 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h32 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h33 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h34 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h35 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h36 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h37 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h38 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h39 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h3a :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h3b :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h3c :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h3d :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h3e :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h3f :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h40 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h41 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h42 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h43 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h44 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h45 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h46 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h47 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h48 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h49 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h4a :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h4b :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h4c :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h4d :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h4e :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h4f :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h50 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h51 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h52 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h53 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h54 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h55 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h56 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h57 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h58 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h59 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h5a :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h5b :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h5c :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h5d :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h5e :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h5f :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h60 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h61 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h62 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h63 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h64 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h65 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h66 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h67 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h68 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h69 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h6a :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h6b :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h6c :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h6d :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h6e :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h6f :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h70 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h71 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h72 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h73 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h74 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h75 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h76 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h77 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h78 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h79 :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h7a :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h7b :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h7c :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h7d :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h7e :
		RG_rl_152_t1 = rl_a46_t8 ;
	7'h7f :
		RG_rl_152_t1 = rl_a46_t8 ;
	default :
		RG_rl_152_t1 = 9'hx ;
	endcase
always @ ( RG_rl_152_t1 or U_318 or TR_219 or U_317 or RG_rl_46 or U_06 or RG_quantized_block_rl_20 or 
	ST1_02d )
	RG_rl_152_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_20 )
		| ( { 9{ U_06 } } & RG_rl_46 )
		| ( { 9{ U_317 } } & TR_219 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_152_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_152_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_152_en )
		RG_rl_152 <= RG_rl_152_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a48_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h01 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h02 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h03 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h04 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h05 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h06 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h07 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h08 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h09 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h0a :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h0b :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h0c :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h0d :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h0e :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h0f :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h10 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h11 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h12 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h13 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h14 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h15 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h16 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h17 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h18 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h19 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h1a :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h1b :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h1c :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h1d :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h1e :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h1f :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h20 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h21 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h22 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h23 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h24 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h25 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h26 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h27 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h28 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h29 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h2a :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h2b :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h2c :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h2d :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h2e :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h2f :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h30 :
		RG_rl_153_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h31 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h32 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h33 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h34 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h35 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h36 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h37 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h38 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h39 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h3a :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h3b :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h3c :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h3d :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h3e :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h3f :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h40 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h41 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h42 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h43 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h44 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h45 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h46 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h47 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h48 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h49 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h4a :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h4b :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h4c :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h4d :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h4e :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h4f :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h50 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h51 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h52 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h53 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h54 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h55 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h56 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h57 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h58 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h59 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h5a :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h5b :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h5c :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h5d :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h5e :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h5f :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h60 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h61 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h62 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h63 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h64 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h65 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h66 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h67 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h68 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h69 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h6a :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h6b :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h6c :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h6d :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h6e :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h6f :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h70 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h71 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h72 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h73 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h74 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h75 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h76 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h77 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h78 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h79 :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h7a :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h7b :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h7c :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h7d :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h7e :
		RG_rl_153_t1 = rl_a48_t8 ;
	7'h7f :
		RG_rl_153_t1 = rl_a48_t8 ;
	default :
		RG_rl_153_t1 = 9'hx ;
	endcase
always @ ( RG_rl_153_t1 or U_318 or TR_217 or U_317 or RG_rl_48 or U_06 or RG_quantized_block_rl_21 or 
	ST1_02d )
	RG_rl_153_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_21 )
		| ( { 9{ U_06 } } & RG_rl_48 )
		| ( { 9{ U_317 } } & TR_217 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_153_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_153_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_153_en )
		RG_rl_153 <= RG_rl_153_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a50_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h01 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h02 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h03 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h04 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h05 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h06 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h07 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h08 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h09 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h0a :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h0b :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h0c :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h0d :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h0e :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h0f :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h10 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h11 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h12 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h13 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h14 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h15 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h16 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h17 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h18 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h19 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h1a :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h1b :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h1c :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h1d :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h1e :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h1f :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h20 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h21 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h22 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h23 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h24 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h25 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h26 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h27 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h28 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h29 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h2a :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h2b :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h2c :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h2d :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h2e :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h2f :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h30 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h31 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h32 :
		RG_rl_154_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h33 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h34 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h35 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h36 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h37 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h38 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h39 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h3a :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h3b :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h3c :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h3d :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h3e :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h3f :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h40 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h41 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h42 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h43 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h44 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h45 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h46 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h47 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h48 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h49 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h4a :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h4b :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h4c :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h4d :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h4e :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h4f :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h50 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h51 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h52 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h53 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h54 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h55 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h56 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h57 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h58 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h59 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h5a :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h5b :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h5c :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h5d :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h5e :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h5f :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h60 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h61 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h62 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h63 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h64 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h65 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h66 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h67 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h68 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h69 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h6a :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h6b :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h6c :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h6d :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h6e :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h6f :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h70 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h71 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h72 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h73 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h74 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h75 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h76 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h77 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h78 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h79 :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h7a :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h7b :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h7c :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h7d :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h7e :
		RG_rl_154_t1 = rl_a50_t8 ;
	7'h7f :
		RG_rl_154_t1 = rl_a50_t8 ;
	default :
		RG_rl_154_t1 = 9'hx ;
	endcase
always @ ( RG_rl_154_t1 or U_318 or TR_215 or U_317 or RG_rl_50 or U_06 or RG_quantized_block_rl_22 or 
	ST1_02d )
	RG_rl_154_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_22 )
		| ( { 9{ U_06 } } & RG_rl_50 )
		| ( { 9{ U_317 } } & TR_215 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_154_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_154_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_154_en )
		RG_rl_154 <= RG_rl_154_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a52_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h01 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h02 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h03 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h04 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h05 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h06 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h07 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h08 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h09 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h0a :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h0b :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h0c :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h0d :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h0e :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h0f :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h10 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h11 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h12 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h13 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h14 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h15 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h16 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h17 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h18 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h19 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h1a :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h1b :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h1c :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h1d :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h1e :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h1f :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h20 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h21 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h22 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h23 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h24 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h25 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h26 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h27 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h28 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h29 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h2a :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h2b :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h2c :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h2d :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h2e :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h2f :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h30 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h31 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h32 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h33 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h34 :
		RG_rl_155_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h35 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h36 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h37 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h38 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h39 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h3a :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h3b :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h3c :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h3d :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h3e :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h3f :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h40 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h41 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h42 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h43 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h44 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h45 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h46 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h47 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h48 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h49 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h4a :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h4b :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h4c :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h4d :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h4e :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h4f :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h50 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h51 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h52 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h53 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h54 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h55 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h56 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h57 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h58 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h59 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h5a :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h5b :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h5c :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h5d :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h5e :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h5f :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h60 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h61 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h62 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h63 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h64 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h65 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h66 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h67 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h68 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h69 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h6a :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h6b :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h6c :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h6d :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h6e :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h6f :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h70 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h71 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h72 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h73 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h74 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h75 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h76 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h77 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h78 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h79 :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h7a :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h7b :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h7c :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h7d :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h7e :
		RG_rl_155_t1 = rl_a52_t8 ;
	7'h7f :
		RG_rl_155_t1 = rl_a52_t8 ;
	default :
		RG_rl_155_t1 = 9'hx ;
	endcase
always @ ( RG_rl_155_t1 or U_318 or TR_213 or U_317 or RG_rl_52 or U_06 or RG_quantized_block_rl_23 or 
	ST1_02d )
	RG_rl_155_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_23 )
		| ( { 9{ U_06 } } & RG_rl_52 )
		| ( { 9{ U_317 } } & TR_213 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_155_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_155_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_155_en )
		RG_rl_155 <= RG_rl_155_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a54_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h01 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h02 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h03 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h04 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h05 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h06 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h07 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h08 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h09 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h0a :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h0b :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h0c :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h0d :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h0e :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h0f :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h10 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h11 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h12 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h13 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h14 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h15 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h16 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h17 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h18 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h19 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h1a :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h1b :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h1c :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h1d :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h1e :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h1f :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h20 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h21 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h22 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h23 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h24 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h25 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h26 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h27 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h28 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h29 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h2a :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h2b :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h2c :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h2d :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h2e :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h2f :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h30 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h31 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h32 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h33 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h34 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h35 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h36 :
		RG_rl_156_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h37 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h38 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h39 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h3a :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h3b :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h3c :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h3d :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h3e :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h3f :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h40 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h41 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h42 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h43 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h44 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h45 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h46 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h47 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h48 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h49 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h4a :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h4b :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h4c :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h4d :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h4e :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h4f :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h50 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h51 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h52 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h53 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h54 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h55 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h56 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h57 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h58 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h59 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h5a :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h5b :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h5c :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h5d :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h5e :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h5f :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h60 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h61 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h62 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h63 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h64 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h65 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h66 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h67 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h68 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h69 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h6a :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h6b :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h6c :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h6d :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h6e :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h6f :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h70 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h71 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h72 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h73 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h74 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h75 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h76 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h77 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h78 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h79 :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h7a :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h7b :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h7c :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h7d :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h7e :
		RG_rl_156_t1 = rl_a54_t8 ;
	7'h7f :
		RG_rl_156_t1 = rl_a54_t8 ;
	default :
		RG_rl_156_t1 = 9'hx ;
	endcase
always @ ( RG_rl_156_t1 or U_318 or TR_211 or U_317 or RG_rl_54 or U_06 or RG_quantized_block_rl_24 or 
	ST1_02d )
	RG_rl_156_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_24 )
		| ( { 9{ U_06 } } & RG_rl_54 )
		| ( { 9{ U_317 } } & TR_211 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_156_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_156_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_156_en )
		RG_rl_156 <= RG_rl_156_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a56_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h01 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h02 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h03 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h04 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h05 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h06 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h07 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h08 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h09 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h0a :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h0b :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h0c :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h0d :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h0e :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h0f :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h10 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h11 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h12 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h13 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h14 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h15 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h16 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h17 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h18 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h19 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h1a :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h1b :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h1c :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h1d :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h1e :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h1f :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h20 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h21 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h22 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h23 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h24 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h25 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h26 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h27 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h28 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h29 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h2a :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h2b :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h2c :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h2d :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h2e :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h2f :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h30 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h31 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h32 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h33 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h34 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h35 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h36 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h37 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h38 :
		RG_rl_157_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h39 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h3a :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h3b :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h3c :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h3d :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h3e :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h3f :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h40 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h41 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h42 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h43 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h44 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h45 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h46 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h47 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h48 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h49 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h4a :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h4b :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h4c :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h4d :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h4e :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h4f :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h50 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h51 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h52 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h53 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h54 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h55 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h56 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h57 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h58 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h59 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h5a :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h5b :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h5c :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h5d :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h5e :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h5f :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h60 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h61 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h62 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h63 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h64 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h65 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h66 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h67 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h68 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h69 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h6a :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h6b :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h6c :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h6d :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h6e :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h6f :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h70 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h71 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h72 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h73 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h74 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h75 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h76 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h77 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h78 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h79 :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h7a :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h7b :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h7c :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h7d :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h7e :
		RG_rl_157_t1 = rl_a56_t8 ;
	7'h7f :
		RG_rl_157_t1 = rl_a56_t8 ;
	default :
		RG_rl_157_t1 = 9'hx ;
	endcase
always @ ( RG_rl_157_t1 or U_318 or TR_209 or U_317 or RG_rl_56 or U_06 or RG_quantized_block_rl_25 or 
	ST1_02d )
	RG_rl_157_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_25 )
		| ( { 9{ U_06 } } & RG_rl_56 )
		| ( { 9{ U_317 } } & TR_209 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_157_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_157_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_157_en )
		RG_rl_157 <= RG_rl_157_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a58_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h01 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h02 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h03 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h04 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h05 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h06 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h07 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h08 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h09 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h0a :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h0b :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h0c :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h0d :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h0e :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h0f :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h10 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h11 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h12 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h13 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h14 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h15 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h16 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h17 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h18 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h19 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h1a :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h1b :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h1c :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h1d :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h1e :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h1f :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h20 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h21 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h22 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h23 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h24 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h25 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h26 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h27 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h28 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h29 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h2a :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h2b :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h2c :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h2d :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h2e :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h2f :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h30 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h31 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h32 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h33 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h34 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h35 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h36 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h37 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h38 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h39 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h3a :
		RG_rl_158_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h3b :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h3c :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h3d :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h3e :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h3f :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h40 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h41 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h42 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h43 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h44 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h45 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h46 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h47 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h48 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h49 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h4a :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h4b :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h4c :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h4d :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h4e :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h4f :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h50 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h51 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h52 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h53 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h54 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h55 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h56 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h57 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h58 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h59 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h5a :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h5b :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h5c :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h5d :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h5e :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h5f :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h60 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h61 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h62 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h63 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h64 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h65 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h66 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h67 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h68 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h69 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h6a :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h6b :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h6c :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h6d :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h6e :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h6f :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h70 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h71 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h72 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h73 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h74 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h75 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h76 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h77 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h78 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h79 :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h7a :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h7b :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h7c :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h7d :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h7e :
		RG_rl_158_t1 = rl_a58_t8 ;
	7'h7f :
		RG_rl_158_t1 = rl_a58_t8 ;
	default :
		RG_rl_158_t1 = 9'hx ;
	endcase
always @ ( RG_rl_158_t1 or U_318 or TR_207 or U_317 or RG_rl_58 or U_06 or RG_quantized_block_rl_26 or 
	ST1_02d )
	RG_rl_158_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_26 )
		| ( { 9{ U_06 } } & RG_rl_58 )
		| ( { 9{ U_317 } } & TR_207 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_158_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_158_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_158_en )
		RG_rl_158 <= RG_rl_158_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a60_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h01 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h02 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h03 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h04 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h05 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h06 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h07 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h08 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h09 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h0a :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h0b :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h0c :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h0d :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h0e :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h0f :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h10 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h11 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h12 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h13 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h14 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h15 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h16 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h17 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h18 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h19 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h1a :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h1b :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h1c :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h1d :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h1e :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h1f :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h20 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h21 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h22 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h23 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h24 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h25 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h26 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h27 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h28 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h29 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h2a :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h2b :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h2c :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h2d :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h2e :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h2f :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h30 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h31 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h32 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h33 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h34 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h35 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h36 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h37 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h38 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h39 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h3a :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h3b :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h3c :
		RG_rl_159_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h3d :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h3e :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h3f :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h40 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h41 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h42 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h43 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h44 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h45 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h46 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h47 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h48 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h49 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h4a :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h4b :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h4c :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h4d :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h4e :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h4f :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h50 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h51 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h52 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h53 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h54 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h55 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h56 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h57 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h58 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h59 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h5a :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h5b :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h5c :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h5d :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h5e :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h5f :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h60 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h61 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h62 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h63 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h64 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h65 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h66 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h67 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h68 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h69 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h6a :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h6b :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h6c :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h6d :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h6e :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h6f :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h70 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h71 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h72 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h73 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h74 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h75 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h76 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h77 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h78 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h79 :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h7a :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h7b :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h7c :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h7d :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h7e :
		RG_rl_159_t1 = rl_a60_t8 ;
	7'h7f :
		RG_rl_159_t1 = rl_a60_t8 ;
	default :
		RG_rl_159_t1 = 9'hx ;
	endcase
always @ ( RG_rl_159_t1 or U_318 or TR_205 or U_317 or RG_rl_60 or U_06 or RG_quantized_block_rl_27 or 
	ST1_02d )
	RG_rl_159_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_27 )
		| ( { 9{ U_06 } } & RG_rl_60 )
		| ( { 9{ U_317 } } & TR_205 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_159_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_159_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_159_en )
		RG_rl_159 <= RG_rl_159_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a62_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h01 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h02 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h03 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h04 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h05 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h06 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h07 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h08 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h09 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h0a :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h0b :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h0c :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h0d :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h0e :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h0f :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h10 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h11 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h12 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h13 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h14 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h15 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h16 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h17 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h18 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h19 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h1a :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h1b :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h1c :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h1d :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h1e :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h1f :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h20 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h21 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h22 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h23 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h24 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h25 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h26 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h27 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h28 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h29 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h2a :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h2b :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h2c :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h2d :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h2e :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h2f :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h30 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h31 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h32 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h33 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h34 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h35 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h36 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h37 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h38 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h39 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h3a :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h3b :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h3c :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h3d :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h3e :
		RG_rl_160_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h3f :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h40 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h41 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h42 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h43 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h44 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h45 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h46 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h47 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h48 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h49 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h4a :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h4b :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h4c :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h4d :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h4e :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h4f :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h50 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h51 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h52 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h53 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h54 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h55 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h56 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h57 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h58 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h59 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h5a :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h5b :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h5c :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h5d :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h5e :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h5f :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h60 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h61 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h62 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h63 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h64 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h65 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h66 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h67 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h68 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h69 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h6a :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h6b :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h6c :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h6d :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h6e :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h6f :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h70 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h71 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h72 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h73 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h74 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h75 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h76 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h77 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h78 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h79 :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h7a :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h7b :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h7c :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h7d :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h7e :
		RG_rl_160_t1 = rl_a62_t8 ;
	7'h7f :
		RG_rl_160_t1 = rl_a62_t8 ;
	default :
		RG_rl_160_t1 = 9'hx ;
	endcase
always @ ( RG_rl_160_t1 or U_318 or TR_203 or U_317 or RG_rl_62 or U_06 or RG_quantized_block_rl_28 or 
	ST1_02d )
	RG_rl_160_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_28 )
		| ( { 9{ U_06 } } & RG_rl_62 )
		| ( { 9{ U_317 } } & TR_203 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_160_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_160_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_160_en )
		RG_rl_160 <= RG_rl_160_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a64_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h01 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h02 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h03 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h04 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h05 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h06 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h07 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h08 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h09 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h0a :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h0b :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h0c :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h0d :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h0e :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h0f :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h10 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h11 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h12 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h13 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h14 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h15 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h16 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h17 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h18 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h19 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h1a :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h1b :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h1c :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h1d :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h1e :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h1f :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h20 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h21 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h22 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h23 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h24 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h25 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h26 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h27 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h28 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h29 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h2a :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h2b :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h2c :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h2d :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h2e :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h2f :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h30 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h31 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h32 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h33 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h34 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h35 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h36 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h37 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h38 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h39 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h3a :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h3b :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h3c :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h3d :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h3e :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h3f :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h40 :
		RG_rl_161_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h41 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h42 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h43 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h44 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h45 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h46 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h47 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h48 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h49 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h4a :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h4b :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h4c :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h4d :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h4e :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h4f :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h50 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h51 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h52 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h53 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h54 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h55 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h56 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h57 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h58 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h59 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h5a :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h5b :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h5c :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h5d :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h5e :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h5f :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h60 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h61 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h62 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h63 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h64 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h65 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h66 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h67 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h68 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h69 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h6a :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h6b :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h6c :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h6d :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h6e :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h6f :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h70 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h71 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h72 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h73 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h74 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h75 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h76 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h77 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h78 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h79 :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h7a :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h7b :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h7c :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h7d :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h7e :
		RG_rl_161_t1 = rl_a64_t8 ;
	7'h7f :
		RG_rl_161_t1 = rl_a64_t8 ;
	default :
		RG_rl_161_t1 = 9'hx ;
	endcase
always @ ( RG_rl_161_t1 or U_318 or TR_201 or U_317 or RG_rl_64 or U_06 or RG_quantized_block_rl_29 or 
	ST1_02d )
	RG_rl_161_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_29 )
		| ( { 9{ U_06 } } & RG_rl_64 )
		| ( { 9{ U_317 } } & TR_201 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_161_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_161_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_161_en )
		RG_rl_161 <= RG_rl_161_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a66_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h01 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h02 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h03 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h04 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h05 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h06 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h07 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h08 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h09 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h0a :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h0b :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h0c :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h0d :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h0e :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h0f :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h10 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h11 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h12 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h13 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h14 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h15 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h16 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h17 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h18 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h19 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h1a :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h1b :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h1c :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h1d :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h1e :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h1f :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h20 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h21 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h22 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h23 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h24 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h25 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h26 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h27 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h28 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h29 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h2a :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h2b :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h2c :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h2d :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h2e :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h2f :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h30 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h31 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h32 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h33 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h34 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h35 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h36 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h37 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h38 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h39 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h3a :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h3b :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h3c :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h3d :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h3e :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h3f :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h40 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h41 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h42 :
		RG_rl_162_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h43 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h44 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h45 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h46 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h47 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h48 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h49 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h4a :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h4b :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h4c :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h4d :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h4e :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h4f :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h50 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h51 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h52 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h53 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h54 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h55 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h56 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h57 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h58 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h59 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h5a :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h5b :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h5c :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h5d :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h5e :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h5f :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h60 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h61 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h62 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h63 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h64 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h65 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h66 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h67 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h68 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h69 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h6a :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h6b :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h6c :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h6d :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h6e :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h6f :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h70 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h71 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h72 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h73 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h74 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h75 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h76 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h77 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h78 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h79 :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h7a :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h7b :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h7c :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h7d :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h7e :
		RG_rl_162_t1 = rl_a66_t8 ;
	7'h7f :
		RG_rl_162_t1 = rl_a66_t8 ;
	default :
		RG_rl_162_t1 = 9'hx ;
	endcase
always @ ( RG_rl_162_t1 or U_318 or TR_199 or U_317 or RG_rl_66 or U_06 or RG_quantized_block_rl_30 or 
	ST1_02d )
	RG_rl_162_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_30 )
		| ( { 9{ U_06 } } & RG_rl_66 )
		| ( { 9{ U_317 } } & TR_199 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_162_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_162_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_162_en )
		RG_rl_162 <= RG_rl_162_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a68_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h01 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h02 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h03 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h04 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h05 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h06 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h07 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h08 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h09 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h0a :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h0b :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h0c :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h0d :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h0e :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h0f :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h10 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h11 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h12 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h13 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h14 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h15 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h16 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h17 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h18 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h19 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h1a :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h1b :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h1c :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h1d :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h1e :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h1f :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h20 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h21 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h22 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h23 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h24 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h25 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h26 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h27 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h28 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h29 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h2a :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h2b :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h2c :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h2d :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h2e :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h2f :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h30 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h31 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h32 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h33 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h34 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h35 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h36 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h37 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h38 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h39 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h3a :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h3b :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h3c :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h3d :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h3e :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h3f :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h40 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h41 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h42 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h43 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h44 :
		RG_rl_163_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h45 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h46 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h47 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h48 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h49 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h4a :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h4b :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h4c :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h4d :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h4e :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h4f :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h50 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h51 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h52 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h53 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h54 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h55 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h56 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h57 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h58 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h59 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h5a :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h5b :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h5c :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h5d :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h5e :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h5f :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h60 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h61 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h62 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h63 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h64 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h65 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h66 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h67 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h68 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h69 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h6a :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h6b :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h6c :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h6d :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h6e :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h6f :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h70 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h71 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h72 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h73 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h74 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h75 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h76 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h77 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h78 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h79 :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h7a :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h7b :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h7c :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h7d :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h7e :
		RG_rl_163_t1 = rl_a68_t8 ;
	7'h7f :
		RG_rl_163_t1 = rl_a68_t8 ;
	default :
		RG_rl_163_t1 = 9'hx ;
	endcase
always @ ( RG_rl_163_t1 or U_318 or TR_197 or U_317 or RG_rl_68 or U_06 or RG_quantized_block_rl_31 or 
	ST1_02d )
	RG_rl_163_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_31 )
		| ( { 9{ U_06 } } & RG_rl_68 )
		| ( { 9{ U_317 } } & TR_197 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_163_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_163_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_163_en )
		RG_rl_163 <= RG_rl_163_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a70_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h01 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h02 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h03 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h04 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h05 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h06 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h07 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h08 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h09 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h0a :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h0b :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h0c :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h0d :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h0e :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h0f :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h10 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h11 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h12 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h13 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h14 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h15 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h16 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h17 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h18 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h19 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h1a :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h1b :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h1c :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h1d :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h1e :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h1f :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h20 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h21 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h22 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h23 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h24 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h25 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h26 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h27 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h28 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h29 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h2a :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h2b :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h2c :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h2d :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h2e :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h2f :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h30 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h31 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h32 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h33 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h34 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h35 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h36 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h37 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h38 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h39 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h3a :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h3b :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h3c :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h3d :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h3e :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h3f :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h40 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h41 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h42 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h43 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h44 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h45 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h46 :
		RG_rl_164_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h47 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h48 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h49 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h4a :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h4b :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h4c :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h4d :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h4e :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h4f :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h50 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h51 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h52 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h53 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h54 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h55 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h56 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h57 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h58 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h59 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h5a :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h5b :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h5c :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h5d :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h5e :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h5f :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h60 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h61 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h62 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h63 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h64 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h65 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h66 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h67 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h68 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h69 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h6a :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h6b :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h6c :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h6d :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h6e :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h6f :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h70 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h71 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h72 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h73 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h74 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h75 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h76 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h77 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h78 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h79 :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h7a :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h7b :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h7c :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h7d :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h7e :
		RG_rl_164_t1 = rl_a70_t8 ;
	7'h7f :
		RG_rl_164_t1 = rl_a70_t8 ;
	default :
		RG_rl_164_t1 = 9'hx ;
	endcase
always @ ( RG_rl_164_t1 or U_318 or TR_195 or U_317 or RG_rl_70 or U_06 or RG_quantized_block_rl_32 or 
	ST1_02d )
	RG_rl_164_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_32 )
		| ( { 9{ U_06 } } & RG_rl_70 )
		| ( { 9{ U_317 } } & TR_195 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_164_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_164_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_164_en )
		RG_rl_164 <= RG_rl_164_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a72_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h01 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h02 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h03 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h04 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h05 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h06 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h07 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h08 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h09 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h0a :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h0b :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h0c :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h0d :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h0e :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h0f :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h10 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h11 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h12 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h13 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h14 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h15 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h16 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h17 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h18 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h19 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h1a :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h1b :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h1c :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h1d :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h1e :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h1f :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h20 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h21 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h22 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h23 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h24 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h25 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h26 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h27 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h28 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h29 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h2a :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h2b :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h2c :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h2d :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h2e :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h2f :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h30 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h31 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h32 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h33 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h34 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h35 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h36 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h37 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h38 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h39 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h3a :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h3b :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h3c :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h3d :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h3e :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h3f :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h40 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h41 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h42 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h43 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h44 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h45 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h46 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h47 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h48 :
		RG_rl_165_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h49 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h4a :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h4b :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h4c :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h4d :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h4e :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h4f :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h50 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h51 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h52 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h53 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h54 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h55 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h56 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h57 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h58 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h59 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h5a :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h5b :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h5c :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h5d :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h5e :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h5f :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h60 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h61 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h62 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h63 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h64 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h65 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h66 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h67 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h68 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h69 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h6a :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h6b :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h6c :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h6d :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h6e :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h6f :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h70 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h71 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h72 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h73 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h74 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h75 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h76 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h77 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h78 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h79 :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h7a :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h7b :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h7c :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h7d :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h7e :
		RG_rl_165_t1 = rl_a72_t8 ;
	7'h7f :
		RG_rl_165_t1 = rl_a72_t8 ;
	default :
		RG_rl_165_t1 = 9'hx ;
	endcase
always @ ( RG_rl_165_t1 or U_318 or TR_193 or U_317 or RG_rl_72 or U_06 or RG_quantized_block_rl_33 or 
	ST1_02d )
	RG_rl_165_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_33 )
		| ( { 9{ U_06 } } & RG_rl_72 )
		| ( { 9{ U_317 } } & TR_193 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_165_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_165_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_165_en )
		RG_rl_165 <= RG_rl_165_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a74_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h01 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h02 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h03 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h04 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h05 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h06 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h07 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h08 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h09 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h0a :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h0b :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h0c :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h0d :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h0e :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h0f :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h10 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h11 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h12 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h13 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h14 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h15 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h16 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h17 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h18 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h19 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h1a :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h1b :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h1c :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h1d :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h1e :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h1f :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h20 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h21 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h22 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h23 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h24 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h25 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h26 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h27 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h28 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h29 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h2a :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h2b :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h2c :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h2d :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h2e :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h2f :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h30 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h31 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h32 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h33 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h34 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h35 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h36 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h37 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h38 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h39 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h3a :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h3b :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h3c :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h3d :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h3e :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h3f :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h40 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h41 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h42 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h43 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h44 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h45 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h46 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h47 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h48 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h49 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h4a :
		RG_rl_166_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h4b :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h4c :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h4d :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h4e :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h4f :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h50 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h51 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h52 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h53 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h54 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h55 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h56 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h57 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h58 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h59 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h5a :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h5b :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h5c :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h5d :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h5e :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h5f :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h60 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h61 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h62 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h63 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h64 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h65 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h66 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h67 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h68 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h69 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h6a :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h6b :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h6c :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h6d :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h6e :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h6f :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h70 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h71 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h72 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h73 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h74 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h75 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h76 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h77 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h78 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h79 :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h7a :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h7b :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h7c :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h7d :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h7e :
		RG_rl_166_t1 = rl_a74_t8 ;
	7'h7f :
		RG_rl_166_t1 = rl_a74_t8 ;
	default :
		RG_rl_166_t1 = 9'hx ;
	endcase
always @ ( RG_rl_166_t1 or U_318 or TR_191 or U_317 or RG_rl_74 or U_06 or RG_quantized_block_rl_34 or 
	ST1_02d )
	RG_rl_166_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_34 )
		| ( { 9{ U_06 } } & RG_rl_74 )
		| ( { 9{ U_317 } } & TR_191 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_166_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_166_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_166_en )
		RG_rl_166 <= RG_rl_166_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a76_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h01 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h02 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h03 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h04 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h05 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h06 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h07 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h08 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h09 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h0a :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h0b :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h0c :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h0d :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h0e :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h0f :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h10 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h11 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h12 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h13 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h14 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h15 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h16 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h17 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h18 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h19 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h1a :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h1b :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h1c :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h1d :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h1e :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h1f :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h20 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h21 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h22 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h23 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h24 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h25 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h26 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h27 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h28 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h29 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h2a :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h2b :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h2c :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h2d :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h2e :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h2f :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h30 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h31 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h32 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h33 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h34 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h35 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h36 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h37 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h38 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h39 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h3a :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h3b :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h3c :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h3d :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h3e :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h3f :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h40 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h41 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h42 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h43 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h44 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h45 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h46 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h47 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h48 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h49 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h4a :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h4b :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h4c :
		RG_rl_167_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h4d :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h4e :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h4f :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h50 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h51 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h52 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h53 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h54 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h55 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h56 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h57 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h58 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h59 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h5a :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h5b :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h5c :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h5d :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h5e :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h5f :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h60 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h61 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h62 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h63 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h64 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h65 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h66 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h67 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h68 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h69 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h6a :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h6b :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h6c :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h6d :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h6e :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h6f :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h70 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h71 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h72 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h73 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h74 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h75 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h76 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h77 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h78 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h79 :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h7a :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h7b :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h7c :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h7d :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h7e :
		RG_rl_167_t1 = rl_a76_t8 ;
	7'h7f :
		RG_rl_167_t1 = rl_a76_t8 ;
	default :
		RG_rl_167_t1 = 9'hx ;
	endcase
always @ ( RG_rl_167_t1 or U_318 or TR_189 or U_317 or RG_rl_76 or U_06 or RG_quantized_block_rl_35 or 
	ST1_02d )
	RG_rl_167_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_35 )
		| ( { 9{ U_06 } } & RG_rl_76 )
		| ( { 9{ U_317 } } & TR_189 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_167_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_167_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_167_en )
		RG_rl_167 <= RG_rl_167_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a78_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h01 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h02 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h03 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h04 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h05 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h06 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h07 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h08 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h09 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h0a :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h0b :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h0c :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h0d :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h0e :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h0f :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h10 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h11 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h12 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h13 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h14 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h15 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h16 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h17 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h18 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h19 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h1a :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h1b :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h1c :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h1d :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h1e :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h1f :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h20 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h21 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h22 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h23 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h24 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h25 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h26 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h27 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h28 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h29 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h2a :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h2b :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h2c :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h2d :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h2e :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h2f :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h30 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h31 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h32 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h33 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h34 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h35 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h36 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h37 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h38 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h39 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h3a :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h3b :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h3c :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h3d :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h3e :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h3f :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h40 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h41 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h42 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h43 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h44 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h45 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h46 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h47 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h48 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h49 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h4a :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h4b :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h4c :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h4d :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h4e :
		RG_rl_168_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h4f :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h50 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h51 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h52 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h53 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h54 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h55 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h56 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h57 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h58 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h59 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h5a :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h5b :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h5c :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h5d :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h5e :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h5f :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h60 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h61 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h62 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h63 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h64 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h65 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h66 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h67 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h68 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h69 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h6a :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h6b :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h6c :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h6d :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h6e :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h6f :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h70 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h71 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h72 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h73 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h74 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h75 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h76 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h77 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h78 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h79 :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h7a :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h7b :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h7c :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h7d :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h7e :
		RG_rl_168_t1 = rl_a78_t8 ;
	7'h7f :
		RG_rl_168_t1 = rl_a78_t8 ;
	default :
		RG_rl_168_t1 = 9'hx ;
	endcase
always @ ( RG_rl_168_t1 or U_318 or TR_187 or U_317 or RG_rl_78 or U_06 or RG_quantized_block_rl_36 or 
	ST1_02d )
	RG_rl_168_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_36 )
		| ( { 9{ U_06 } } & RG_rl_78 )
		| ( { 9{ U_317 } } & TR_187 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_168_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_168_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_168_en )
		RG_rl_168 <= RG_rl_168_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a80_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h01 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h02 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h03 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h04 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h05 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h06 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h07 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h08 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h09 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h0a :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h0b :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h0c :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h0d :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h0e :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h0f :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h10 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h11 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h12 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h13 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h14 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h15 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h16 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h17 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h18 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h19 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h1a :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h1b :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h1c :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h1d :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h1e :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h1f :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h20 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h21 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h22 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h23 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h24 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h25 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h26 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h27 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h28 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h29 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h2a :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h2b :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h2c :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h2d :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h2e :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h2f :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h30 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h31 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h32 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h33 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h34 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h35 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h36 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h37 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h38 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h39 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h3a :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h3b :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h3c :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h3d :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h3e :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h3f :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h40 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h41 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h42 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h43 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h44 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h45 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h46 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h47 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h48 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h49 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h4a :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h4b :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h4c :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h4d :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h4e :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h4f :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h50 :
		RG_rl_169_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h51 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h52 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h53 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h54 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h55 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h56 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h57 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h58 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h59 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h5a :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h5b :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h5c :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h5d :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h5e :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h5f :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h60 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h61 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h62 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h63 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h64 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h65 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h66 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h67 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h68 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h69 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h6a :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h6b :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h6c :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h6d :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h6e :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h6f :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h70 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h71 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h72 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h73 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h74 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h75 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h76 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h77 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h78 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h79 :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h7a :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h7b :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h7c :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h7d :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h7e :
		RG_rl_169_t1 = rl_a80_t8 ;
	7'h7f :
		RG_rl_169_t1 = rl_a80_t8 ;
	default :
		RG_rl_169_t1 = 9'hx ;
	endcase
always @ ( RG_rl_169_t1 or U_318 or TR_185 or U_317 or RG_rl_80 or U_06 or RG_quantized_block_rl_37 or 
	ST1_02d )
	RG_rl_169_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_37 )
		| ( { 9{ U_06 } } & RG_rl_80 )
		| ( { 9{ U_317 } } & TR_185 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_169_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_169_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_169_en )
		RG_rl_169 <= RG_rl_169_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a82_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h01 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h02 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h03 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h04 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h05 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h06 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h07 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h08 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h09 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h0a :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h0b :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h0c :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h0d :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h0e :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h0f :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h10 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h11 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h12 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h13 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h14 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h15 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h16 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h17 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h18 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h19 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h1a :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h1b :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h1c :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h1d :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h1e :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h1f :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h20 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h21 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h22 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h23 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h24 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h25 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h26 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h27 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h28 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h29 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h2a :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h2b :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h2c :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h2d :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h2e :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h2f :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h30 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h31 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h32 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h33 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h34 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h35 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h36 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h37 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h38 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h39 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h3a :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h3b :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h3c :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h3d :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h3e :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h3f :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h40 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h41 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h42 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h43 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h44 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h45 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h46 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h47 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h48 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h49 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h4a :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h4b :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h4c :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h4d :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h4e :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h4f :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h50 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h51 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h52 :
		RG_rl_170_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h53 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h54 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h55 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h56 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h57 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h58 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h59 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h5a :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h5b :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h5c :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h5d :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h5e :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h5f :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h60 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h61 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h62 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h63 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h64 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h65 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h66 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h67 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h68 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h69 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h6a :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h6b :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h6c :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h6d :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h6e :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h6f :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h70 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h71 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h72 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h73 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h74 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h75 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h76 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h77 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h78 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h79 :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h7a :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h7b :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h7c :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h7d :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h7e :
		RG_rl_170_t1 = rl_a82_t8 ;
	7'h7f :
		RG_rl_170_t1 = rl_a82_t8 ;
	default :
		RG_rl_170_t1 = 9'hx ;
	endcase
always @ ( RG_rl_170_t1 or U_318 or TR_183 or U_317 or RG_rl_82 or U_06 or RG_quantized_block_rl_38 or 
	ST1_02d )
	RG_rl_170_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_38 )
		| ( { 9{ U_06 } } & RG_rl_82 )
		| ( { 9{ U_317 } } & TR_183 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_170_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_170_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_170_en )
		RG_rl_170 <= RG_rl_170_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a84_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h01 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h02 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h03 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h04 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h05 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h06 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h07 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h08 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h09 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h0a :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h0b :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h0c :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h0d :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h0e :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h0f :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h10 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h11 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h12 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h13 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h14 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h15 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h16 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h17 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h18 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h19 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h1a :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h1b :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h1c :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h1d :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h1e :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h1f :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h20 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h21 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h22 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h23 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h24 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h25 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h26 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h27 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h28 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h29 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h2a :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h2b :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h2c :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h2d :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h2e :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h2f :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h30 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h31 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h32 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h33 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h34 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h35 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h36 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h37 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h38 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h39 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h3a :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h3b :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h3c :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h3d :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h3e :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h3f :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h40 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h41 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h42 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h43 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h44 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h45 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h46 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h47 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h48 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h49 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h4a :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h4b :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h4c :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h4d :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h4e :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h4f :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h50 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h51 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h52 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h53 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h54 :
		RG_rl_171_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h55 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h56 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h57 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h58 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h59 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h5a :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h5b :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h5c :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h5d :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h5e :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h5f :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h60 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h61 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h62 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h63 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h64 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h65 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h66 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h67 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h68 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h69 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h6a :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h6b :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h6c :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h6d :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h6e :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h6f :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h70 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h71 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h72 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h73 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h74 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h75 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h76 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h77 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h78 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h79 :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h7a :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h7b :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h7c :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h7d :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h7e :
		RG_rl_171_t1 = rl_a84_t8 ;
	7'h7f :
		RG_rl_171_t1 = rl_a84_t8 ;
	default :
		RG_rl_171_t1 = 9'hx ;
	endcase
always @ ( RG_rl_171_t1 or U_318 or TR_181 or U_317 or RG_rl_84 or U_06 or RG_quantized_block_rl_39 or 
	ST1_02d )
	RG_rl_171_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_39 )
		| ( { 9{ U_06 } } & RG_rl_84 )
		| ( { 9{ U_317 } } & TR_181 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_171_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_171_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_171_en )
		RG_rl_171 <= RG_rl_171_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a86_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h01 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h02 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h03 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h04 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h05 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h06 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h07 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h08 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h09 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h0a :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h0b :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h0c :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h0d :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h0e :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h0f :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h10 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h11 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h12 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h13 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h14 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h15 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h16 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h17 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h18 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h19 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h1a :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h1b :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h1c :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h1d :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h1e :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h1f :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h20 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h21 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h22 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h23 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h24 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h25 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h26 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h27 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h28 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h29 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h2a :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h2b :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h2c :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h2d :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h2e :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h2f :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h30 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h31 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h32 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h33 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h34 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h35 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h36 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h37 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h38 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h39 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h3a :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h3b :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h3c :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h3d :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h3e :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h3f :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h40 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h41 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h42 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h43 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h44 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h45 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h46 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h47 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h48 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h49 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h4a :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h4b :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h4c :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h4d :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h4e :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h4f :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h50 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h51 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h52 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h53 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h54 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h55 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h56 :
		RG_rl_172_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h57 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h58 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h59 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h5a :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h5b :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h5c :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h5d :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h5e :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h5f :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h60 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h61 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h62 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h63 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h64 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h65 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h66 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h67 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h68 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h69 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h6a :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h6b :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h6c :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h6d :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h6e :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h6f :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h70 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h71 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h72 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h73 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h74 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h75 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h76 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h77 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h78 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h79 :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h7a :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h7b :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h7c :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h7d :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h7e :
		RG_rl_172_t1 = rl_a86_t8 ;
	7'h7f :
		RG_rl_172_t1 = rl_a86_t8 ;
	default :
		RG_rl_172_t1 = 9'hx ;
	endcase
always @ ( RG_rl_172_t1 or U_318 or TR_179 or U_317 or RG_rl_86 or U_06 or RG_quantized_block_rl_40 or 
	ST1_02d )
	RG_rl_172_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_40 )
		| ( { 9{ U_06 } } & RG_rl_86 )
		| ( { 9{ U_317 } } & TR_179 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_172_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_172_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_172_en )
		RG_rl_172 <= RG_rl_172_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a88_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h01 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h02 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h03 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h04 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h05 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h06 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h07 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h08 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h09 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h0a :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h0b :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h0c :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h0d :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h0e :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h0f :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h10 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h11 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h12 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h13 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h14 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h15 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h16 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h17 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h18 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h19 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h1a :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h1b :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h1c :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h1d :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h1e :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h1f :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h20 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h21 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h22 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h23 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h24 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h25 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h26 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h27 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h28 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h29 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h2a :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h2b :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h2c :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h2d :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h2e :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h2f :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h30 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h31 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h32 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h33 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h34 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h35 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h36 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h37 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h38 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h39 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h3a :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h3b :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h3c :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h3d :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h3e :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h3f :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h40 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h41 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h42 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h43 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h44 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h45 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h46 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h47 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h48 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h49 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h4a :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h4b :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h4c :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h4d :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h4e :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h4f :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h50 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h51 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h52 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h53 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h54 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h55 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h56 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h57 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h58 :
		RG_rl_173_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h59 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h5a :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h5b :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h5c :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h5d :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h5e :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h5f :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h60 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h61 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h62 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h63 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h64 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h65 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h66 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h67 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h68 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h69 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h6a :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h6b :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h6c :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h6d :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h6e :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h6f :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h70 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h71 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h72 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h73 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h74 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h75 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h76 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h77 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h78 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h79 :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h7a :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h7b :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h7c :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h7d :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h7e :
		RG_rl_173_t1 = rl_a88_t8 ;
	7'h7f :
		RG_rl_173_t1 = rl_a88_t8 ;
	default :
		RG_rl_173_t1 = 9'hx ;
	endcase
always @ ( RG_rl_173_t1 or U_318 or TR_177 or U_317 or RG_rl_88 or U_06 or RG_quantized_block_rl_41 or 
	ST1_02d )
	RG_rl_173_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_41 )
		| ( { 9{ U_06 } } & RG_rl_88 )
		| ( { 9{ U_317 } } & TR_177 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_173_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_173_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_173_en )
		RG_rl_173 <= RG_rl_173_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a90_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h01 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h02 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h03 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h04 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h05 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h06 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h07 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h08 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h09 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h0a :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h0b :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h0c :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h0d :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h0e :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h0f :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h10 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h11 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h12 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h13 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h14 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h15 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h16 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h17 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h18 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h19 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h1a :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h1b :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h1c :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h1d :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h1e :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h1f :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h20 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h21 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h22 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h23 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h24 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h25 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h26 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h27 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h28 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h29 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h2a :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h2b :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h2c :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h2d :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h2e :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h2f :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h30 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h31 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h32 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h33 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h34 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h35 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h36 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h37 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h38 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h39 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h3a :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h3b :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h3c :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h3d :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h3e :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h3f :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h40 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h41 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h42 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h43 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h44 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h45 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h46 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h47 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h48 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h49 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h4a :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h4b :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h4c :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h4d :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h4e :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h4f :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h50 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h51 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h52 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h53 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h54 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h55 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h56 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h57 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h58 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h59 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h5a :
		RG_rl_174_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h5b :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h5c :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h5d :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h5e :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h5f :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h60 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h61 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h62 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h63 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h64 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h65 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h66 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h67 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h68 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h69 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h6a :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h6b :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h6c :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h6d :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h6e :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h6f :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h70 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h71 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h72 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h73 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h74 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h75 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h76 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h77 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h78 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h79 :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h7a :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h7b :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h7c :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h7d :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h7e :
		RG_rl_174_t1 = rl_a90_t8 ;
	7'h7f :
		RG_rl_174_t1 = rl_a90_t8 ;
	default :
		RG_rl_174_t1 = 9'hx ;
	endcase
always @ ( RG_rl_174_t1 or U_318 or TR_175 or U_317 or RG_rl_90 or U_06 or RG_quantized_block_rl_42 or 
	ST1_02d )
	RG_rl_174_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_42 )
		| ( { 9{ U_06 } } & RG_rl_90 )
		| ( { 9{ U_317 } } & TR_175 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_174_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_174_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_174_en )
		RG_rl_174 <= RG_rl_174_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a92_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h01 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h02 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h03 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h04 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h05 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h06 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h07 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h08 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h09 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h0a :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h0b :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h0c :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h0d :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h0e :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h0f :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h10 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h11 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h12 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h13 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h14 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h15 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h16 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h17 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h18 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h19 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h1a :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h1b :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h1c :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h1d :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h1e :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h1f :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h20 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h21 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h22 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h23 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h24 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h25 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h26 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h27 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h28 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h29 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h2a :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h2b :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h2c :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h2d :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h2e :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h2f :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h30 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h31 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h32 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h33 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h34 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h35 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h36 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h37 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h38 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h39 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h3a :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h3b :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h3c :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h3d :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h3e :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h3f :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h40 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h41 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h42 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h43 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h44 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h45 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h46 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h47 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h48 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h49 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h4a :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h4b :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h4c :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h4d :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h4e :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h4f :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h50 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h51 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h52 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h53 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h54 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h55 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h56 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h57 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h58 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h59 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h5a :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h5b :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h5c :
		RG_rl_175_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h5d :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h5e :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h5f :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h60 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h61 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h62 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h63 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h64 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h65 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h66 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h67 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h68 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h69 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h6a :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h6b :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h6c :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h6d :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h6e :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h6f :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h70 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h71 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h72 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h73 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h74 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h75 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h76 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h77 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h78 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h79 :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h7a :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h7b :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h7c :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h7d :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h7e :
		RG_rl_175_t1 = rl_a92_t8 ;
	7'h7f :
		RG_rl_175_t1 = rl_a92_t8 ;
	default :
		RG_rl_175_t1 = 9'hx ;
	endcase
always @ ( RG_rl_175_t1 or U_318 or TR_173 or U_317 or RG_rl_92 or U_06 or RG_quantized_block_rl_43 or 
	ST1_02d )
	RG_rl_175_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_43 )
		| ( { 9{ U_06 } } & RG_rl_92 )
		| ( { 9{ U_317 } } & TR_173 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_175_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_175_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_175_en )
		RG_rl_175 <= RG_rl_175_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a94_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h01 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h02 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h03 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h04 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h05 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h06 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h07 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h08 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h09 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h0a :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h0b :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h0c :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h0d :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h0e :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h0f :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h10 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h11 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h12 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h13 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h14 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h15 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h16 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h17 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h18 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h19 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h1a :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h1b :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h1c :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h1d :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h1e :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h1f :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h20 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h21 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h22 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h23 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h24 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h25 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h26 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h27 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h28 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h29 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h2a :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h2b :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h2c :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h2d :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h2e :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h2f :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h30 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h31 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h32 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h33 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h34 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h35 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h36 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h37 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h38 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h39 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h3a :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h3b :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h3c :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h3d :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h3e :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h3f :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h40 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h41 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h42 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h43 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h44 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h45 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h46 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h47 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h48 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h49 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h4a :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h4b :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h4c :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h4d :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h4e :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h4f :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h50 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h51 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h52 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h53 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h54 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h55 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h56 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h57 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h58 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h59 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h5a :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h5b :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h5c :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h5d :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h5e :
		RG_rl_176_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h5f :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h60 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h61 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h62 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h63 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h64 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h65 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h66 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h67 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h68 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h69 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h6a :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h6b :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h6c :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h6d :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h6e :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h6f :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h70 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h71 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h72 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h73 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h74 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h75 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h76 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h77 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h78 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h79 :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h7a :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h7b :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h7c :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h7d :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h7e :
		RG_rl_176_t1 = rl_a94_t8 ;
	7'h7f :
		RG_rl_176_t1 = rl_a94_t8 ;
	default :
		RG_rl_176_t1 = 9'hx ;
	endcase
always @ ( RG_rl_176_t1 or U_318 or TR_171 or U_317 or RG_rl_94 or U_06 or RG_quantized_block_rl_44 or 
	ST1_02d )
	RG_rl_176_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_44 )
		| ( { 9{ U_06 } } & RG_rl_94 )
		| ( { 9{ U_317 } } & TR_171 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_176_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_176_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_176_en )
		RG_rl_176 <= RG_rl_176_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a96_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h01 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h02 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h03 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h04 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h05 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h06 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h07 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h08 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h09 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h0a :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h0b :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h0c :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h0d :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h0e :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h0f :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h10 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h11 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h12 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h13 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h14 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h15 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h16 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h17 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h18 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h19 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h1a :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h1b :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h1c :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h1d :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h1e :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h1f :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h20 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h21 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h22 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h23 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h24 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h25 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h26 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h27 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h28 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h29 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h2a :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h2b :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h2c :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h2d :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h2e :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h2f :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h30 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h31 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h32 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h33 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h34 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h35 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h36 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h37 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h38 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h39 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h3a :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h3b :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h3c :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h3d :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h3e :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h3f :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h40 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h41 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h42 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h43 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h44 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h45 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h46 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h47 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h48 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h49 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h4a :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h4b :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h4c :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h4d :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h4e :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h4f :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h50 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h51 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h52 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h53 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h54 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h55 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h56 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h57 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h58 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h59 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h5a :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h5b :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h5c :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h5d :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h5e :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h5f :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h60 :
		RG_rl_177_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h61 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h62 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h63 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h64 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h65 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h66 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h67 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h68 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h69 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h6a :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h6b :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h6c :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h6d :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h6e :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h6f :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h70 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h71 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h72 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h73 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h74 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h75 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h76 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h77 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h78 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h79 :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h7a :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h7b :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h7c :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h7d :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h7e :
		RG_rl_177_t1 = rl_a96_t8 ;
	7'h7f :
		RG_rl_177_t1 = rl_a96_t8 ;
	default :
		RG_rl_177_t1 = 9'hx ;
	endcase
always @ ( RG_rl_177_t1 or U_318 or TR_169 or U_317 or RG_rl_96 or U_06 or RG_quantized_block_rl_45 or 
	ST1_02d )
	RG_rl_177_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_45 )
		| ( { 9{ U_06 } } & RG_rl_96 )
		| ( { 9{ U_317 } } & TR_169 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_177_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_177_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_177_en )
		RG_rl_177 <= RG_rl_177_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a98_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h01 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h02 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h03 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h04 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h05 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h06 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h07 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h08 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h09 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h0a :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h0b :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h0c :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h0d :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h0e :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h0f :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h10 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h11 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h12 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h13 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h14 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h15 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h16 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h17 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h18 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h19 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h1a :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h1b :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h1c :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h1d :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h1e :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h1f :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h20 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h21 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h22 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h23 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h24 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h25 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h26 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h27 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h28 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h29 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h2a :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h2b :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h2c :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h2d :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h2e :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h2f :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h30 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h31 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h32 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h33 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h34 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h35 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h36 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h37 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h38 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h39 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h3a :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h3b :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h3c :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h3d :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h3e :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h3f :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h40 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h41 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h42 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h43 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h44 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h45 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h46 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h47 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h48 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h49 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h4a :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h4b :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h4c :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h4d :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h4e :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h4f :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h50 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h51 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h52 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h53 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h54 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h55 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h56 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h57 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h58 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h59 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h5a :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h5b :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h5c :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h5d :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h5e :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h5f :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h60 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h61 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h62 :
		RG_rl_178_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h63 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h64 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h65 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h66 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h67 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h68 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h69 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h6a :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h6b :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h6c :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h6d :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h6e :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h6f :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h70 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h71 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h72 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h73 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h74 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h75 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h76 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h77 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h78 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h79 :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h7a :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h7b :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h7c :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h7d :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h7e :
		RG_rl_178_t1 = rl_a98_t8 ;
	7'h7f :
		RG_rl_178_t1 = rl_a98_t8 ;
	default :
		RG_rl_178_t1 = 9'hx ;
	endcase
always @ ( RG_rl_178_t1 or U_318 or TR_167 or U_317 or RG_rl_98 or U_06 or RG_quantized_block_rl_46 or 
	ST1_02d )
	RG_rl_178_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_46 )
		| ( { 9{ U_06 } } & RG_rl_98 )
		| ( { 9{ U_317 } } & TR_167 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_178_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_178_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_178_en )
		RG_rl_178 <= RG_rl_178_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a100_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h01 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h02 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h03 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h04 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h05 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h06 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h07 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h08 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h09 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h0a :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h0b :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h0c :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h0d :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h0e :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h0f :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h10 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h11 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h12 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h13 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h14 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h15 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h16 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h17 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h18 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h19 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h1a :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h1b :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h1c :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h1d :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h1e :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h1f :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h20 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h21 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h22 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h23 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h24 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h25 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h26 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h27 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h28 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h29 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h2a :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h2b :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h2c :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h2d :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h2e :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h2f :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h30 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h31 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h32 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h33 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h34 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h35 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h36 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h37 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h38 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h39 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h3a :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h3b :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h3c :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h3d :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h3e :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h3f :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h40 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h41 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h42 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h43 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h44 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h45 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h46 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h47 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h48 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h49 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h4a :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h4b :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h4c :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h4d :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h4e :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h4f :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h50 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h51 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h52 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h53 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h54 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h55 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h56 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h57 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h58 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h59 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h5a :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h5b :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h5c :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h5d :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h5e :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h5f :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h60 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h61 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h62 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h63 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h64 :
		RG_rl_179_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h65 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h66 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h67 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h68 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h69 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h6a :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h6b :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h6c :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h6d :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h6e :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h6f :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h70 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h71 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h72 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h73 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h74 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h75 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h76 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h77 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h78 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h79 :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h7a :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h7b :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h7c :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h7d :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h7e :
		RG_rl_179_t1 = rl_a100_t8 ;
	7'h7f :
		RG_rl_179_t1 = rl_a100_t8 ;
	default :
		RG_rl_179_t1 = 9'hx ;
	endcase
always @ ( RG_rl_179_t1 or U_318 or TR_165 or U_317 or RG_rl_100 or U_06 or RG_quantized_block_rl_47 or 
	ST1_02d )
	RG_rl_179_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_47 )
		| ( { 9{ U_06 } } & RG_rl_100 )
		| ( { 9{ U_317 } } & TR_165 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_179_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_179_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_179_en )
		RG_rl_179 <= RG_rl_179_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a102_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h01 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h02 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h03 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h04 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h05 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h06 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h07 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h08 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h09 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h0a :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h0b :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h0c :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h0d :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h0e :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h0f :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h10 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h11 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h12 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h13 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h14 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h15 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h16 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h17 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h18 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h19 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h1a :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h1b :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h1c :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h1d :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h1e :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h1f :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h20 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h21 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h22 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h23 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h24 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h25 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h26 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h27 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h28 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h29 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h2a :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h2b :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h2c :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h2d :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h2e :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h2f :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h30 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h31 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h32 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h33 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h34 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h35 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h36 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h37 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h38 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h39 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h3a :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h3b :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h3c :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h3d :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h3e :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h3f :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h40 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h41 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h42 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h43 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h44 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h45 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h46 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h47 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h48 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h49 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h4a :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h4b :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h4c :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h4d :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h4e :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h4f :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h50 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h51 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h52 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h53 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h54 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h55 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h56 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h57 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h58 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h59 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h5a :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h5b :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h5c :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h5d :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h5e :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h5f :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h60 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h61 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h62 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h63 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h64 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h65 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h66 :
		RG_rl_180_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h67 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h68 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h69 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h6a :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h6b :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h6c :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h6d :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h6e :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h6f :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h70 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h71 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h72 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h73 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h74 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h75 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h76 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h77 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h78 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h79 :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h7a :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h7b :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h7c :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h7d :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h7e :
		RG_rl_180_t1 = rl_a102_t8 ;
	7'h7f :
		RG_rl_180_t1 = rl_a102_t8 ;
	default :
		RG_rl_180_t1 = 9'hx ;
	endcase
always @ ( RG_rl_180_t1 or U_318 or TR_163 or U_317 or RG_rl_102 or U_06 or RG_quantized_block_rl_48 or 
	ST1_02d )
	RG_rl_180_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_48 )
		| ( { 9{ U_06 } } & RG_rl_102 )
		| ( { 9{ U_317 } } & TR_163 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_180_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_180_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_180_en )
		RG_rl_180 <= RG_rl_180_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a104_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h01 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h02 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h03 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h04 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h05 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h06 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h07 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h08 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h09 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h0a :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h0b :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h0c :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h0d :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h0e :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h0f :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h10 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h11 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h12 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h13 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h14 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h15 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h16 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h17 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h18 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h19 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h1a :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h1b :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h1c :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h1d :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h1e :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h1f :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h20 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h21 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h22 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h23 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h24 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h25 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h26 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h27 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h28 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h29 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h2a :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h2b :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h2c :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h2d :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h2e :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h2f :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h30 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h31 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h32 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h33 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h34 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h35 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h36 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h37 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h38 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h39 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h3a :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h3b :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h3c :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h3d :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h3e :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h3f :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h40 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h41 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h42 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h43 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h44 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h45 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h46 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h47 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h48 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h49 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h4a :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h4b :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h4c :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h4d :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h4e :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h4f :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h50 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h51 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h52 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h53 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h54 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h55 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h56 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h57 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h58 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h59 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h5a :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h5b :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h5c :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h5d :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h5e :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h5f :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h60 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h61 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h62 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h63 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h64 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h65 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h66 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h67 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h68 :
		RG_rl_181_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h69 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h6a :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h6b :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h6c :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h6d :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h6e :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h6f :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h70 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h71 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h72 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h73 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h74 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h75 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h76 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h77 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h78 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h79 :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h7a :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h7b :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h7c :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h7d :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h7e :
		RG_rl_181_t1 = rl_a104_t8 ;
	7'h7f :
		RG_rl_181_t1 = rl_a104_t8 ;
	default :
		RG_rl_181_t1 = 9'hx ;
	endcase
always @ ( RG_rl_181_t1 or U_318 or TR_161 or U_317 or RG_rl_104 or U_06 or RG_quantized_block_rl_49 or 
	ST1_02d )
	RG_rl_181_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_49 )
		| ( { 9{ U_06 } } & RG_rl_104 )
		| ( { 9{ U_317 } } & TR_161 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_181_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_181_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_181_en )
		RG_rl_181 <= RG_rl_181_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a106_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h01 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h02 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h03 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h04 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h05 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h06 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h07 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h08 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h09 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h0a :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h0b :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h0c :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h0d :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h0e :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h0f :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h10 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h11 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h12 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h13 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h14 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h15 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h16 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h17 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h18 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h19 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h1a :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h1b :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h1c :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h1d :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h1e :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h1f :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h20 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h21 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h22 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h23 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h24 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h25 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h26 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h27 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h28 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h29 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h2a :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h2b :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h2c :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h2d :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h2e :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h2f :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h30 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h31 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h32 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h33 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h34 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h35 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h36 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h37 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h38 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h39 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h3a :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h3b :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h3c :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h3d :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h3e :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h3f :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h40 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h41 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h42 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h43 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h44 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h45 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h46 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h47 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h48 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h49 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h4a :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h4b :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h4c :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h4d :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h4e :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h4f :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h50 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h51 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h52 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h53 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h54 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h55 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h56 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h57 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h58 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h59 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h5a :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h5b :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h5c :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h5d :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h5e :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h5f :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h60 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h61 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h62 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h63 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h64 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h65 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h66 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h67 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h68 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h69 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h6a :
		RG_rl_182_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h6b :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h6c :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h6d :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h6e :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h6f :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h70 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h71 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h72 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h73 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h74 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h75 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h76 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h77 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h78 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h79 :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h7a :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h7b :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h7c :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h7d :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h7e :
		RG_rl_182_t1 = rl_a106_t8 ;
	7'h7f :
		RG_rl_182_t1 = rl_a106_t8 ;
	default :
		RG_rl_182_t1 = 9'hx ;
	endcase
always @ ( RG_rl_182_t1 or U_318 or TR_159 or U_317 or RG_rl_106 or U_06 or RG_quantized_block_rl_50 or 
	ST1_02d )
	RG_rl_182_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_50 )
		| ( { 9{ U_06 } } & RG_rl_106 )
		| ( { 9{ U_317 } } & TR_159 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_182_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_182_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_182_en )
		RG_rl_182 <= RG_rl_182_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a108_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h01 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h02 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h03 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h04 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h05 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h06 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h07 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h08 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h09 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h0a :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h0b :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h0c :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h0d :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h0e :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h0f :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h10 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h11 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h12 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h13 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h14 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h15 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h16 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h17 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h18 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h19 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h1a :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h1b :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h1c :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h1d :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h1e :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h1f :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h20 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h21 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h22 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h23 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h24 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h25 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h26 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h27 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h28 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h29 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h2a :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h2b :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h2c :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h2d :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h2e :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h2f :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h30 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h31 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h32 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h33 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h34 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h35 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h36 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h37 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h38 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h39 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h3a :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h3b :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h3c :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h3d :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h3e :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h3f :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h40 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h41 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h42 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h43 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h44 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h45 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h46 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h47 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h48 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h49 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h4a :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h4b :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h4c :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h4d :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h4e :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h4f :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h50 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h51 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h52 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h53 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h54 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h55 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h56 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h57 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h58 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h59 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h5a :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h5b :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h5c :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h5d :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h5e :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h5f :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h60 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h61 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h62 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h63 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h64 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h65 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h66 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h67 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h68 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h69 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h6a :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h6b :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h6c :
		RG_rl_183_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h6d :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h6e :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h6f :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h70 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h71 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h72 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h73 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h74 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h75 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h76 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h77 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h78 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h79 :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h7a :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h7b :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h7c :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h7d :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h7e :
		RG_rl_183_t1 = rl_a108_t8 ;
	7'h7f :
		RG_rl_183_t1 = rl_a108_t8 ;
	default :
		RG_rl_183_t1 = 9'hx ;
	endcase
always @ ( RG_rl_183_t1 or U_318 or TR_157 or U_317 or RG_rl_108 or U_06 or RG_quantized_block_rl_51 or 
	ST1_02d )
	RG_rl_183_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_51 )
		| ( { 9{ U_06 } } & RG_rl_108 )
		| ( { 9{ U_317 } } & TR_157 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_183_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_183_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_183_en )
		RG_rl_183 <= RG_rl_183_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a110_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h01 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h02 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h03 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h04 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h05 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h06 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h07 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h08 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h09 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h0a :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h0b :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h0c :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h0d :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h0e :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h0f :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h10 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h11 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h12 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h13 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h14 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h15 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h16 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h17 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h18 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h19 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h1a :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h1b :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h1c :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h1d :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h1e :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h1f :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h20 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h21 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h22 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h23 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h24 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h25 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h26 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h27 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h28 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h29 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h2a :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h2b :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h2c :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h2d :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h2e :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h2f :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h30 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h31 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h32 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h33 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h34 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h35 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h36 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h37 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h38 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h39 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h3a :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h3b :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h3c :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h3d :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h3e :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h3f :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h40 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h41 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h42 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h43 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h44 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h45 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h46 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h47 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h48 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h49 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h4a :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h4b :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h4c :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h4d :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h4e :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h4f :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h50 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h51 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h52 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h53 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h54 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h55 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h56 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h57 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h58 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h59 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h5a :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h5b :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h5c :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h5d :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h5e :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h5f :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h60 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h61 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h62 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h63 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h64 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h65 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h66 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h67 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h68 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h69 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h6a :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h6b :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h6c :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h6d :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h6e :
		RG_rl_184_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h6f :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h70 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h71 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h72 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h73 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h74 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h75 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h76 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h77 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h78 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h79 :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h7a :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h7b :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h7c :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h7d :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h7e :
		RG_rl_184_t1 = rl_a110_t8 ;
	7'h7f :
		RG_rl_184_t1 = rl_a110_t8 ;
	default :
		RG_rl_184_t1 = 9'hx ;
	endcase
always @ ( RG_rl_184_t1 or U_318 or TR_155 or U_317 or RG_rl_110 or U_06 or RG_quantized_block_rl_52 or 
	ST1_02d )
	RG_rl_184_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_52 )
		| ( { 9{ U_06 } } & RG_rl_110 )
		| ( { 9{ U_317 } } & TR_155 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_184_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_184_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_184_en )
		RG_rl_184 <= RG_rl_184_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a112_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h01 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h02 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h03 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h04 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h05 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h06 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h07 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h08 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h09 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h0a :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h0b :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h0c :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h0d :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h0e :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h0f :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h10 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h11 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h12 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h13 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h14 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h15 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h16 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h17 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h18 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h19 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h1a :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h1b :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h1c :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h1d :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h1e :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h1f :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h20 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h21 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h22 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h23 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h24 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h25 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h26 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h27 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h28 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h29 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h2a :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h2b :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h2c :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h2d :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h2e :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h2f :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h30 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h31 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h32 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h33 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h34 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h35 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h36 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h37 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h38 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h39 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h3a :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h3b :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h3c :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h3d :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h3e :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h3f :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h40 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h41 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h42 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h43 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h44 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h45 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h46 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h47 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h48 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h49 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h4a :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h4b :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h4c :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h4d :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h4e :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h4f :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h50 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h51 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h52 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h53 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h54 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h55 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h56 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h57 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h58 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h59 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h5a :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h5b :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h5c :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h5d :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h5e :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h5f :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h60 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h61 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h62 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h63 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h64 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h65 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h66 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h67 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h68 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h69 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h6a :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h6b :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h6c :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h6d :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h6e :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h6f :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h70 :
		RG_rl_185_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h71 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h72 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h73 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h74 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h75 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h76 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h77 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h78 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h79 :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h7a :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h7b :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h7c :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h7d :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h7e :
		RG_rl_185_t1 = rl_a112_t8 ;
	7'h7f :
		RG_rl_185_t1 = rl_a112_t8 ;
	default :
		RG_rl_185_t1 = 9'hx ;
	endcase
always @ ( RG_rl_185_t1 or U_318 or TR_153 or U_317 or RG_rl_112 or U_06 or RG_quantized_block_rl_53 or 
	ST1_02d )
	RG_rl_185_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_53 )
		| ( { 9{ U_06 } } & RG_rl_112 )
		| ( { 9{ U_317 } } & TR_153 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_185_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_185_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_185_en )
		RG_rl_185 <= RG_rl_185_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a114_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h01 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h02 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h03 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h04 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h05 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h06 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h07 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h08 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h09 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h0a :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h0b :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h0c :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h0d :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h0e :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h0f :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h10 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h11 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h12 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h13 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h14 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h15 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h16 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h17 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h18 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h19 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h1a :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h1b :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h1c :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h1d :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h1e :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h1f :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h20 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h21 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h22 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h23 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h24 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h25 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h26 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h27 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h28 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h29 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h2a :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h2b :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h2c :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h2d :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h2e :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h2f :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h30 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h31 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h32 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h33 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h34 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h35 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h36 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h37 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h38 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h39 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h3a :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h3b :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h3c :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h3d :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h3e :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h3f :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h40 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h41 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h42 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h43 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h44 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h45 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h46 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h47 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h48 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h49 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h4a :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h4b :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h4c :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h4d :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h4e :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h4f :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h50 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h51 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h52 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h53 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h54 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h55 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h56 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h57 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h58 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h59 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h5a :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h5b :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h5c :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h5d :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h5e :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h5f :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h60 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h61 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h62 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h63 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h64 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h65 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h66 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h67 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h68 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h69 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h6a :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h6b :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h6c :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h6d :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h6e :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h6f :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h70 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h71 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h72 :
		RG_rl_186_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h73 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h74 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h75 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h76 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h77 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h78 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h79 :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h7a :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h7b :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h7c :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h7d :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h7e :
		RG_rl_186_t1 = rl_a114_t8 ;
	7'h7f :
		RG_rl_186_t1 = rl_a114_t8 ;
	default :
		RG_rl_186_t1 = 9'hx ;
	endcase
always @ ( RG_rl_186_t1 or U_318 or TR_151 or U_317 or RG_rl_114 or U_06 or RG_quantized_block_rl_54 or 
	ST1_02d )
	RG_rl_186_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_54 )
		| ( { 9{ U_06 } } & RG_rl_114 )
		| ( { 9{ U_317 } } & TR_151 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_186_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_186_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_186_en )
		RG_rl_186 <= RG_rl_186_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a116_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h01 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h02 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h03 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h04 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h05 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h06 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h07 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h08 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h09 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h0a :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h0b :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h0c :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h0d :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h0e :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h0f :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h10 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h11 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h12 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h13 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h14 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h15 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h16 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h17 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h18 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h19 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h1a :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h1b :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h1c :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h1d :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h1e :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h1f :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h20 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h21 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h22 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h23 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h24 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h25 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h26 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h27 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h28 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h29 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h2a :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h2b :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h2c :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h2d :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h2e :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h2f :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h30 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h31 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h32 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h33 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h34 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h35 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h36 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h37 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h38 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h39 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h3a :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h3b :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h3c :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h3d :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h3e :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h3f :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h40 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h41 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h42 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h43 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h44 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h45 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h46 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h47 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h48 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h49 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h4a :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h4b :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h4c :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h4d :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h4e :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h4f :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h50 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h51 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h52 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h53 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h54 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h55 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h56 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h57 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h58 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h59 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h5a :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h5b :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h5c :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h5d :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h5e :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h5f :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h60 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h61 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h62 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h63 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h64 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h65 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h66 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h67 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h68 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h69 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h6a :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h6b :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h6c :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h6d :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h6e :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h6f :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h70 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h71 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h72 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h73 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h74 :
		RG_rl_187_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h75 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h76 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h77 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h78 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h79 :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h7a :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h7b :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h7c :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h7d :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h7e :
		RG_rl_187_t1 = rl_a116_t8 ;
	7'h7f :
		RG_rl_187_t1 = rl_a116_t8 ;
	default :
		RG_rl_187_t1 = 9'hx ;
	endcase
always @ ( RG_rl_187_t1 or U_318 or TR_149 or U_317 or RG_rl_116 or U_06 or RG_quantized_block_rl_55 or 
	ST1_02d )
	RG_rl_187_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_55 )
		| ( { 9{ U_06 } } & RG_rl_116 )
		| ( { 9{ U_317 } } & TR_149 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_187_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_187_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_187_en )
		RG_rl_187 <= RG_rl_187_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a118_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h01 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h02 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h03 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h04 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h05 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h06 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h07 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h08 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h09 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h0a :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h0b :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h0c :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h0d :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h0e :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h0f :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h10 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h11 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h12 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h13 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h14 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h15 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h16 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h17 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h18 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h19 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h1a :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h1b :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h1c :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h1d :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h1e :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h1f :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h20 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h21 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h22 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h23 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h24 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h25 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h26 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h27 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h28 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h29 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h2a :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h2b :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h2c :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h2d :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h2e :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h2f :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h30 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h31 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h32 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h33 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h34 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h35 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h36 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h37 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h38 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h39 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h3a :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h3b :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h3c :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h3d :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h3e :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h3f :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h40 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h41 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h42 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h43 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h44 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h45 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h46 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h47 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h48 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h49 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h4a :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h4b :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h4c :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h4d :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h4e :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h4f :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h50 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h51 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h52 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h53 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h54 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h55 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h56 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h57 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h58 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h59 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h5a :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h5b :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h5c :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h5d :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h5e :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h5f :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h60 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h61 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h62 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h63 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h64 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h65 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h66 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h67 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h68 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h69 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h6a :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h6b :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h6c :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h6d :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h6e :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h6f :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h70 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h71 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h72 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h73 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h74 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h75 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h76 :
		RG_rl_188_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h77 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h78 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h79 :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h7a :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h7b :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h7c :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h7d :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h7e :
		RG_rl_188_t1 = rl_a118_t8 ;
	7'h7f :
		RG_rl_188_t1 = rl_a118_t8 ;
	default :
		RG_rl_188_t1 = 9'hx ;
	endcase
always @ ( RG_rl_188_t1 or U_318 or TR_147 or U_317 or RG_rl_118 or U_06 or RG_quantized_block_rl_56 or 
	ST1_02d )
	RG_rl_188_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_56 )
		| ( { 9{ U_06 } } & RG_rl_118 )
		| ( { 9{ U_317 } } & TR_147 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_188_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_188_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_188_en )
		RG_rl_188 <= RG_rl_188_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a120_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h01 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h02 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h03 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h04 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h05 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h06 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h07 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h08 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h09 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h0a :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h0b :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h0c :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h0d :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h0e :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h0f :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h10 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h11 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h12 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h13 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h14 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h15 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h16 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h17 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h18 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h19 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h1a :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h1b :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h1c :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h1d :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h1e :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h1f :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h20 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h21 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h22 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h23 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h24 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h25 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h26 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h27 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h28 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h29 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h2a :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h2b :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h2c :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h2d :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h2e :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h2f :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h30 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h31 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h32 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h33 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h34 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h35 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h36 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h37 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h38 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h39 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h3a :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h3b :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h3c :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h3d :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h3e :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h3f :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h40 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h41 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h42 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h43 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h44 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h45 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h46 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h47 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h48 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h49 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h4a :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h4b :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h4c :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h4d :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h4e :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h4f :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h50 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h51 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h52 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h53 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h54 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h55 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h56 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h57 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h58 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h59 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h5a :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h5b :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h5c :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h5d :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h5e :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h5f :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h60 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h61 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h62 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h63 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h64 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h65 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h66 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h67 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h68 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h69 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h6a :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h6b :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h6c :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h6d :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h6e :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h6f :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h70 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h71 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h72 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h73 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h74 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h75 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h76 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h77 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h78 :
		RG_rl_189_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h79 :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h7a :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h7b :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h7c :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h7d :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h7e :
		RG_rl_189_t1 = rl_a120_t8 ;
	7'h7f :
		RG_rl_189_t1 = rl_a120_t8 ;
	default :
		RG_rl_189_t1 = 9'hx ;
	endcase
always @ ( RG_rl_189_t1 or U_318 or TR_145 or U_317 or RG_rl_120 or U_06 or RG_quantized_block_rl_57 or 
	ST1_02d )
	RG_rl_189_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_57 )
		| ( { 9{ U_06 } } & RG_rl_120 )
		| ( { 9{ U_317 } } & TR_145 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_189_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_189_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_189_en )
		RG_rl_189 <= RG_rl_189_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a122_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h01 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h02 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h03 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h04 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h05 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h06 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h07 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h08 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h09 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h0a :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h0b :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h0c :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h0d :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h0e :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h0f :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h10 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h11 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h12 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h13 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h14 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h15 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h16 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h17 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h18 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h19 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h1a :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h1b :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h1c :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h1d :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h1e :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h1f :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h20 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h21 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h22 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h23 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h24 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h25 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h26 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h27 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h28 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h29 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h2a :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h2b :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h2c :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h2d :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h2e :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h2f :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h30 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h31 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h32 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h33 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h34 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h35 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h36 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h37 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h38 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h39 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h3a :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h3b :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h3c :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h3d :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h3e :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h3f :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h40 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h41 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h42 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h43 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h44 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h45 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h46 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h47 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h48 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h49 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h4a :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h4b :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h4c :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h4d :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h4e :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h4f :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h50 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h51 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h52 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h53 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h54 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h55 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h56 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h57 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h58 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h59 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h5a :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h5b :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h5c :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h5d :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h5e :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h5f :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h60 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h61 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h62 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h63 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h64 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h65 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h66 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h67 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h68 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h69 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h6a :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h6b :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h6c :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h6d :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h6e :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h6f :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h70 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h71 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h72 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h73 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h74 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h75 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h76 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h77 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h78 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h79 :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h7a :
		RG_rl_190_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h7b :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h7c :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h7d :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h7e :
		RG_rl_190_t1 = rl_a122_t8 ;
	7'h7f :
		RG_rl_190_t1 = rl_a122_t8 ;
	default :
		RG_rl_190_t1 = 9'hx ;
	endcase
always @ ( RG_rl_190_t1 or U_318 or TR_143 or U_317 or RG_rl_122 or U_06 or RG_quantized_block_rl_58 or 
	ST1_02d )
	RG_rl_190_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_58 )
		| ( { 9{ U_06 } } & RG_rl_122 )
		| ( { 9{ U_317 } } & TR_143 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_190_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_190_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_190_en )
		RG_rl_190 <= RG_rl_190_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( M_16_t or rl_a124_t8 or incr8u2ot )	// line#=../rle.cpp:73,74
	case ( incr8u2ot [6:0] )
	7'h00 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h01 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h02 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h03 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h04 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h05 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h06 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h07 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h08 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h09 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h0a :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h0b :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h0c :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h0d :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h0e :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h0f :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h10 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h11 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h12 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h13 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h14 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h15 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h16 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h17 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h18 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h19 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h1a :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h1b :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h1c :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h1d :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h1e :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h1f :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h20 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h21 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h22 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h23 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h24 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h25 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h26 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h27 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h28 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h29 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h2a :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h2b :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h2c :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h2d :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h2e :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h2f :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h30 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h31 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h32 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h33 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h34 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h35 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h36 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h37 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h38 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h39 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h3a :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h3b :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h3c :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h3d :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h3e :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h3f :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h40 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h41 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h42 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h43 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h44 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h45 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h46 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h47 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h48 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h49 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h4a :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h4b :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h4c :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h4d :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h4e :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h4f :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h50 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h51 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h52 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h53 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h54 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h55 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h56 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h57 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h58 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h59 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h5a :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h5b :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h5c :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h5d :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h5e :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h5f :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h60 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h61 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h62 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h63 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h64 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h65 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h66 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h67 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h68 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h69 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h6a :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h6b :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h6c :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h6d :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h6e :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h6f :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h70 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h71 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h72 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h73 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h74 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h75 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h76 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h77 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h78 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h79 :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h7a :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h7b :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h7c :
		RG_rl_191_t1 = M_16_t ;	// line#=../rle.cpp:74
	7'h7d :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h7e :
		RG_rl_191_t1 = rl_a124_t8 ;
	7'h7f :
		RG_rl_191_t1 = rl_a124_t8 ;
	default :
		RG_rl_191_t1 = 9'hx ;
	endcase
always @ ( RG_rl_191_t1 or U_318 or TR_141 or U_317 or RG_rl_124 or U_06 or RG_quantized_block_rl_zz or 
	ST1_02d )
	RG_rl_191_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl_zz )
		| ( { 9{ U_06 } } & RG_rl_124 )
		| ( { 9{ U_317 } } & TR_141 )		// line#=../rle.cpp:68,69
		| ( { 9{ U_318 } } & RG_rl_191_t1 )	// line#=../rle.cpp:73,74
		) ;
assign	RG_rl_191_en = ( ST1_02d | U_06 | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_rl_191_en )
		RG_rl_191 <= RG_rl_191_t ;	// line#=../rle.cpp:68,69,73,74
always @ ( incr8u3ot or U_318 or incr8u4ot or U_317 or FF_i or ST1_04d )
	RG_len_t = ( ( { 8{ ST1_04d } } & { 7'h00 , FF_i } )
		| ( { 8{ U_317 } } & incr8u4ot )	// line#=../rle.cpp:69
		| ( { 8{ U_318 } } & incr8u3ot )	// line#=../rle.cpp:74
		) ;
assign	RG_len_en = ( ST1_04d | U_317 | U_318 ) ;
always @ ( posedge clk )
	if ( RG_len_en )
		RG_len <= RG_len_t ;	// line#=../rle.cpp:69,74
always @ ( sub8u1ot or ST1_07d or RG_len or U_174 or incr8u4ot or U_173 )
	RG_len_1_t = ( ( { 8{ U_173 } } & incr8u4ot )	// line#=../rle.cpp:80
		| ( { 8{ U_174 } } & RG_len )
		| ( { 8{ ST1_07d } } & sub8u1ot )	// line#=../rle.cpp:86
		) ;
always @ ( posedge clk )
	RG_len_1 <= RG_len_1_t ;	// line#=../rle.cpp:80,86
always @ ( incr8u3ot or ST1_04d or RG_k or ST1_03d )
	RG_k_1_t = ( ( { 7{ ST1_03d } } & { 1'h0 , RG_k } )
		| ( { 7{ ST1_04d } } & incr8u3ot [6:0] )	// line#=../rle.cpp:142
		) ;
always @ ( posedge clk )
	RG_k_1 <= RG_k_1_t ;	// line#=../rle.cpp:142
assign	JF_01 = ~C_01 ;	// line#=../rle.cpp:35
always @ ( RG_quantized_block_rl_7 or RG_quantized_block_rl_6 or RG_quantized_block_rl_5 or 
	RG_quantized_block_rl_4 or RG_quantized_block_rl_3 or RG_quantized_block_rl_2 or 
	RG_quantized_block_rl_1 or RG_quantized_block_rl or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_04 = RG_quantized_block_rl ;	// line#=../rle.cpp:111
	3'h1 :
		TR_04 = RG_quantized_block_rl_1 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_04 = RG_quantized_block_rl_2 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_04 = RG_quantized_block_rl_3 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_04 = RG_quantized_block_rl_4 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_04 = RG_quantized_block_rl_5 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_04 = RG_quantized_block_rl_6 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_04 = RG_quantized_block_rl_7 ;	// line#=../rle.cpp:111
	default :
		TR_04 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_15 or RG_quantized_block_rl_14 or RG_quantized_block_rl_13 or 
	RG_quantized_block_rl_12 or RG_quantized_block_rl_11 or RG_quantized_block_rl_10 or 
	RG_quantized_block_rl_9 or RG_quantized_block_rl_8 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_05 = RG_quantized_block_rl_8 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_05 = RG_quantized_block_rl_9 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_05 = RG_quantized_block_rl_10 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_05 = RG_quantized_block_rl_11 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_05 = RG_quantized_block_rl_12 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_05 = RG_quantized_block_rl_13 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_05 = RG_quantized_block_rl_14 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_05 = RG_quantized_block_rl_15 ;	// line#=../rle.cpp:111
	default :
		TR_05 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_23 or RG_quantized_block_rl_22 or RG_quantized_block_rl_21 or 
	RG_quantized_block_rl_20 or RG_quantized_block_rl_19 or RG_quantized_block_rl_18 or 
	RG_quantized_block_rl_17 or RG_quantized_block_rl_16 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_06 = RG_quantized_block_rl_16 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_06 = RG_quantized_block_rl_17 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_06 = RG_quantized_block_rl_18 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_06 = RG_quantized_block_rl_19 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_06 = RG_quantized_block_rl_20 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_06 = RG_quantized_block_rl_21 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_06 = RG_quantized_block_rl_22 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_06 = RG_quantized_block_rl_23 ;	// line#=../rle.cpp:111
	default :
		TR_06 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_31 or RG_quantized_block_rl_30 or RG_quantized_block_rl_29 or 
	RG_quantized_block_rl_28 or RG_quantized_block_rl_27 or RG_quantized_block_rl_26 or 
	RG_quantized_block_rl_25 or RG_quantized_block_rl_24 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_07 = RG_quantized_block_rl_24 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_07 = RG_quantized_block_rl_25 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_07 = RG_quantized_block_rl_26 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_07 = RG_quantized_block_rl_27 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_07 = RG_quantized_block_rl_28 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_07 = RG_quantized_block_rl_29 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_07 = RG_quantized_block_rl_30 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_07 = RG_quantized_block_rl_31 ;	// line#=../rle.cpp:111
	default :
		TR_07 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_39 or RG_quantized_block_rl_38 or RG_quantized_block_rl_37 or 
	RG_quantized_block_rl_36 or RG_quantized_block_rl_35 or RG_quantized_block_rl_34 or 
	RG_quantized_block_rl_33 or RG_quantized_block_rl_32 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_08 = RG_quantized_block_rl_32 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_08 = RG_quantized_block_rl_33 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_08 = RG_quantized_block_rl_34 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_08 = RG_quantized_block_rl_35 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_08 = RG_quantized_block_rl_36 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_08 = RG_quantized_block_rl_37 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_08 = RG_quantized_block_rl_38 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_08 = RG_quantized_block_rl_39 ;	// line#=../rle.cpp:111
	default :
		TR_08 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_47 or RG_quantized_block_rl_46 or RG_quantized_block_rl_45 or 
	RG_quantized_block_rl_44 or RG_quantized_block_rl_43 or RG_quantized_block_rl_42 or 
	RG_quantized_block_rl_41 or RG_quantized_block_rl_40 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_09 = RG_quantized_block_rl_40 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_09 = RG_quantized_block_rl_41 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_09 = RG_quantized_block_rl_42 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_09 = RG_quantized_block_rl_43 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_09 = RG_quantized_block_rl_44 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_09 = RG_quantized_block_rl_45 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_09 = RG_quantized_block_rl_46 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_09 = RG_quantized_block_rl_47 ;	// line#=../rle.cpp:111
	default :
		TR_09 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_55 or RG_quantized_block_rl_54 or RG_quantized_block_rl_53 or 
	RG_quantized_block_rl_52 or RG_quantized_block_rl_51 or RG_quantized_block_rl_50 or 
	RG_quantized_block_rl_49 or RG_quantized_block_rl_48 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_10 = RG_quantized_block_rl_48 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_10 = RG_quantized_block_rl_49 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_10 = RG_quantized_block_rl_50 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_10 = RG_quantized_block_rl_51 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_10 = RG_quantized_block_rl_52 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_10 = RG_quantized_block_rl_53 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_10 = RG_quantized_block_rl_54 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_10 = RG_quantized_block_rl_55 ;	// line#=../rle.cpp:111
	default :
		TR_10 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_zz or RG_k_quantized_block_rl_01 or RG_quantized_block_rl_61 or 
	RG_quantized_block_rl_60 or RG_quantized_block_rl_59 or RG_quantized_block_rl_58 or 
	RG_quantized_block_rl_57 or RG_quantized_block_rl_56 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_11 = RG_quantized_block_rl_56 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_11 = RG_quantized_block_rl_57 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_11 = RG_quantized_block_rl_58 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_11 = RG_quantized_block_rl_59 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_11 = RG_quantized_block_rl_60 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_11 = RG_quantized_block_rl_61 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_11 = RG_k_quantized_block_rl_01 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_11 = RG_quantized_block_rl_zz ;	// line#=../rle.cpp:111
	default :
		TR_11 = 9'hx ;
	endcase
always @ ( TR_11 or TR_10 or TR_09 or TR_08 or TR_07 or TR_06 or TR_05 or TR_04 or 
	RG_i_k_01 )	// line#=../rle.cpp:111,142
	begin
	M_184_c1 = ~|RG_i_k_01 [2:0] ;	// line#=../rle.cpp:111,142
	M_184_c2 = ~|( RG_i_k_01 [2:0] ^ 3'h1 ) ;	// line#=../rle.cpp:111,142
	M_184_c3 = ~|( RG_i_k_01 [2:0] ^ 3'h2 ) ;	// line#=../rle.cpp:111,142
	M_184_c4 = ~|( RG_i_k_01 [2:0] ^ 3'h3 ) ;	// line#=../rle.cpp:111,142
	M_184_c5 = ~|( RG_i_k_01 [2:0] ^ 3'h4 ) ;	// line#=../rle.cpp:111,142
	M_184_c6 = ~|( RG_i_k_01 [2:0] ^ 3'h5 ) ;	// line#=../rle.cpp:111,142
	M_184_c7 = ~|( RG_i_k_01 [2:0] ^ 3'h6 ) ;	// line#=../rle.cpp:111,142
	M_184_c8 = ~|( RG_i_k_01 [2:0] ^ 3'h7 ) ;	// line#=../rle.cpp:111,142
	M_184 = ( ( { 9{ M_184_c1 } } & TR_04 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_184_c2 } } & TR_05 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_184_c3 } } & TR_06 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_184_c4 } } & TR_07 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_184_c5 } } & TR_08 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_184_c6 } } & TR_09 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_184_c7 } } & TR_10 )	// line#=../rle.cpp:111,142
		| ( { 9{ M_184_c8 } } & TR_11 )	// line#=../rle.cpp:111,142
		) ;
	end
assign	JF_03 = ~RG_k_1 [6] ;
always @ ( M_113 or M_112 or M_110 or M_179 or M_109 or M_178 or M_108 or M_177 or 
	M_107 or M_176 or M_106 or M_175 or M_105 or M_174 or M_104 or M_173 or 
	M_103 or M_172 or M_102 or M_171 or M_100 or M_170 or M_99 or M_169 or M_98 or 
	M_168 or M_97 or M_167 or M_96 or M_166 or M_95 or M_165 or M_94 or M_164 or 
	M_93 or M_163 or M_92 or M_162 or M_91 or M_161 or M_90 or M_160 or M_89 or 
	M_159 or M_88 or M_158 or M_87 or M_157 or M_86 or M_156 or M_85 or M_155 or 
	M_84 or M_154 or M_83 or M_153 or M_82 or M_152 or M_81 or M_151 or M_80 or 
	M_150 or M_79 or M_149 or M_78 or M_148 or M_77 or M_147 or M_76 or M_146 or 
	M_75 or M_145 or M_74 or M_144 or M_73 or M_143 or M_72 or M_142 or M_71 or 
	M_141 or M_70 or M_140 or M_69 or M_139 or M_68 or M_138 or M_67 or M_137 or 
	M_66 or M_136 or M_65 or M_135 or M_64 or M_134 or M_63 or M_133 or M_62 or 
	M_132 or M_61 or M_131 or M_60 or M_130 or M_59 or M_129 or M_58 or M_128 or 
	M_57 or M_127 or M_56 or M_126 or M_55 or M_125 or M_54 or M_124 or M_53 or 
	M_123 or M_52 or M_122 or M_51 or M_120 or M_50 or M_119 or M_49 or M_118 or 
	M_117 or M_116 or M_115 or M_114 or sub8u_7_11ot )	// line#=../rle.cpp:77,78
	case ( sub8u_7_11ot )
	7'h00 :
		M_02_t128_t1 = M_114 ;	// line#=../rle.cpp:77,78
	7'h01 :
		M_02_t128_t1 = M_115 ;	// line#=../rle.cpp:77,78
	7'h02 :
		M_02_t128_t1 = M_116 ;	// line#=../rle.cpp:77,78
	7'h03 :
		M_02_t128_t1 = M_117 ;	// line#=../rle.cpp:77,78
	7'h04 :
		M_02_t128_t1 = M_118 ;	// line#=../rle.cpp:77,78
	7'h05 :
		M_02_t128_t1 = M_49 ;	// line#=../rle.cpp:77,78
	7'h06 :
		M_02_t128_t1 = M_119 ;	// line#=../rle.cpp:77,78
	7'h07 :
		M_02_t128_t1 = M_50 ;	// line#=../rle.cpp:77,78
	7'h08 :
		M_02_t128_t1 = M_120 ;	// line#=../rle.cpp:77,78
	7'h09 :
		M_02_t128_t1 = M_51 ;	// line#=../rle.cpp:77,78
	7'h0a :
		M_02_t128_t1 = M_122 ;	// line#=../rle.cpp:77,78
	7'h0b :
		M_02_t128_t1 = M_52 ;	// line#=../rle.cpp:77,78
	7'h0c :
		M_02_t128_t1 = M_123 ;	// line#=../rle.cpp:77,78
	7'h0d :
		M_02_t128_t1 = M_53 ;	// line#=../rle.cpp:77,78
	7'h0e :
		M_02_t128_t1 = M_124 ;	// line#=../rle.cpp:77,78
	7'h0f :
		M_02_t128_t1 = M_54 ;	// line#=../rle.cpp:77,78
	7'h10 :
		M_02_t128_t1 = M_125 ;	// line#=../rle.cpp:77,78
	7'h11 :
		M_02_t128_t1 = M_55 ;	// line#=../rle.cpp:77,78
	7'h12 :
		M_02_t128_t1 = M_126 ;	// line#=../rle.cpp:77,78
	7'h13 :
		M_02_t128_t1 = M_56 ;	// line#=../rle.cpp:77,78
	7'h14 :
		M_02_t128_t1 = M_127 ;	// line#=../rle.cpp:77,78
	7'h15 :
		M_02_t128_t1 = M_57 ;	// line#=../rle.cpp:77,78
	7'h16 :
		M_02_t128_t1 = M_128 ;	// line#=../rle.cpp:77,78
	7'h17 :
		M_02_t128_t1 = M_58 ;	// line#=../rle.cpp:77,78
	7'h18 :
		M_02_t128_t1 = M_129 ;	// line#=../rle.cpp:77,78
	7'h19 :
		M_02_t128_t1 = M_59 ;	// line#=../rle.cpp:77,78
	7'h1a :
		M_02_t128_t1 = M_130 ;	// line#=../rle.cpp:77,78
	7'h1b :
		M_02_t128_t1 = M_60 ;	// line#=../rle.cpp:77,78
	7'h1c :
		M_02_t128_t1 = M_131 ;	// line#=../rle.cpp:77,78
	7'h1d :
		M_02_t128_t1 = M_61 ;	// line#=../rle.cpp:77,78
	7'h1e :
		M_02_t128_t1 = M_132 ;	// line#=../rle.cpp:77,78
	7'h1f :
		M_02_t128_t1 = M_62 ;	// line#=../rle.cpp:77,78
	7'h20 :
		M_02_t128_t1 = M_133 ;	// line#=../rle.cpp:77,78
	7'h21 :
		M_02_t128_t1 = M_63 ;	// line#=../rle.cpp:77,78
	7'h22 :
		M_02_t128_t1 = M_134 ;	// line#=../rle.cpp:77,78
	7'h23 :
		M_02_t128_t1 = M_64 ;	// line#=../rle.cpp:77,78
	7'h24 :
		M_02_t128_t1 = M_135 ;	// line#=../rle.cpp:77,78
	7'h25 :
		M_02_t128_t1 = M_65 ;	// line#=../rle.cpp:77,78
	7'h26 :
		M_02_t128_t1 = M_136 ;	// line#=../rle.cpp:77,78
	7'h27 :
		M_02_t128_t1 = M_66 ;	// line#=../rle.cpp:77,78
	7'h28 :
		M_02_t128_t1 = M_137 ;	// line#=../rle.cpp:77,78
	7'h29 :
		M_02_t128_t1 = M_67 ;	// line#=../rle.cpp:77,78
	7'h2a :
		M_02_t128_t1 = M_138 ;	// line#=../rle.cpp:77,78
	7'h2b :
		M_02_t128_t1 = M_68 ;	// line#=../rle.cpp:77,78
	7'h2c :
		M_02_t128_t1 = M_139 ;	// line#=../rle.cpp:77,78
	7'h2d :
		M_02_t128_t1 = M_69 ;	// line#=../rle.cpp:77,78
	7'h2e :
		M_02_t128_t1 = M_140 ;	// line#=../rle.cpp:77,78
	7'h2f :
		M_02_t128_t1 = M_70 ;	// line#=../rle.cpp:77,78
	7'h30 :
		M_02_t128_t1 = M_141 ;	// line#=../rle.cpp:77,78
	7'h31 :
		M_02_t128_t1 = M_71 ;	// line#=../rle.cpp:77,78
	7'h32 :
		M_02_t128_t1 = M_142 ;	// line#=../rle.cpp:77,78
	7'h33 :
		M_02_t128_t1 = M_72 ;	// line#=../rle.cpp:77,78
	7'h34 :
		M_02_t128_t1 = M_143 ;	// line#=../rle.cpp:77,78
	7'h35 :
		M_02_t128_t1 = M_73 ;	// line#=../rle.cpp:77,78
	7'h36 :
		M_02_t128_t1 = M_144 ;	// line#=../rle.cpp:77,78
	7'h37 :
		M_02_t128_t1 = M_74 ;	// line#=../rle.cpp:77,78
	7'h38 :
		M_02_t128_t1 = M_145 ;	// line#=../rle.cpp:77,78
	7'h39 :
		M_02_t128_t1 = M_75 ;	// line#=../rle.cpp:77,78
	7'h3a :
		M_02_t128_t1 = M_146 ;	// line#=../rle.cpp:77,78
	7'h3b :
		M_02_t128_t1 = M_76 ;	// line#=../rle.cpp:77,78
	7'h3c :
		M_02_t128_t1 = M_147 ;	// line#=../rle.cpp:77,78
	7'h3d :
		M_02_t128_t1 = M_77 ;	// line#=../rle.cpp:77,78
	7'h3e :
		M_02_t128_t1 = M_148 ;	// line#=../rle.cpp:77,78
	7'h3f :
		M_02_t128_t1 = M_78 ;	// line#=../rle.cpp:77,78
	7'h40 :
		M_02_t128_t1 = M_149 ;	// line#=../rle.cpp:77,78
	7'h41 :
		M_02_t128_t1 = M_79 ;	// line#=../rle.cpp:77,78
	7'h42 :
		M_02_t128_t1 = M_150 ;	// line#=../rle.cpp:77,78
	7'h43 :
		M_02_t128_t1 = M_80 ;	// line#=../rle.cpp:77,78
	7'h44 :
		M_02_t128_t1 = M_151 ;	// line#=../rle.cpp:77,78
	7'h45 :
		M_02_t128_t1 = M_81 ;	// line#=../rle.cpp:77,78
	7'h46 :
		M_02_t128_t1 = M_152 ;	// line#=../rle.cpp:77,78
	7'h47 :
		M_02_t128_t1 = M_82 ;	// line#=../rle.cpp:77,78
	7'h48 :
		M_02_t128_t1 = M_153 ;	// line#=../rle.cpp:77,78
	7'h49 :
		M_02_t128_t1 = M_83 ;	// line#=../rle.cpp:77,78
	7'h4a :
		M_02_t128_t1 = M_154 ;	// line#=../rle.cpp:77,78
	7'h4b :
		M_02_t128_t1 = M_84 ;	// line#=../rle.cpp:77,78
	7'h4c :
		M_02_t128_t1 = M_155 ;	// line#=../rle.cpp:77,78
	7'h4d :
		M_02_t128_t1 = M_85 ;	// line#=../rle.cpp:77,78
	7'h4e :
		M_02_t128_t1 = M_156 ;	// line#=../rle.cpp:77,78
	7'h4f :
		M_02_t128_t1 = M_86 ;	// line#=../rle.cpp:77,78
	7'h50 :
		M_02_t128_t1 = M_157 ;	// line#=../rle.cpp:77,78
	7'h51 :
		M_02_t128_t1 = M_87 ;	// line#=../rle.cpp:77,78
	7'h52 :
		M_02_t128_t1 = M_158 ;	// line#=../rle.cpp:77,78
	7'h53 :
		M_02_t128_t1 = M_88 ;	// line#=../rle.cpp:77,78
	7'h54 :
		M_02_t128_t1 = M_159 ;	// line#=../rle.cpp:77,78
	7'h55 :
		M_02_t128_t1 = M_89 ;	// line#=../rle.cpp:77,78
	7'h56 :
		M_02_t128_t1 = M_160 ;	// line#=../rle.cpp:77,78
	7'h57 :
		M_02_t128_t1 = M_90 ;	// line#=../rle.cpp:77,78
	7'h58 :
		M_02_t128_t1 = M_161 ;	// line#=../rle.cpp:77,78
	7'h59 :
		M_02_t128_t1 = M_91 ;	// line#=../rle.cpp:77,78
	7'h5a :
		M_02_t128_t1 = M_162 ;	// line#=../rle.cpp:77,78
	7'h5b :
		M_02_t128_t1 = M_92 ;	// line#=../rle.cpp:77,78
	7'h5c :
		M_02_t128_t1 = M_163 ;	// line#=../rle.cpp:77,78
	7'h5d :
		M_02_t128_t1 = M_93 ;	// line#=../rle.cpp:77,78
	7'h5e :
		M_02_t128_t1 = M_164 ;	// line#=../rle.cpp:77,78
	7'h5f :
		M_02_t128_t1 = M_94 ;	// line#=../rle.cpp:77,78
	7'h60 :
		M_02_t128_t1 = M_165 ;	// line#=../rle.cpp:77,78
	7'h61 :
		M_02_t128_t1 = M_95 ;	// line#=../rle.cpp:77,78
	7'h62 :
		M_02_t128_t1 = M_166 ;	// line#=../rle.cpp:77,78
	7'h63 :
		M_02_t128_t1 = M_96 ;	// line#=../rle.cpp:77,78
	7'h64 :
		M_02_t128_t1 = M_167 ;	// line#=../rle.cpp:77,78
	7'h65 :
		M_02_t128_t1 = M_97 ;	// line#=../rle.cpp:77,78
	7'h66 :
		M_02_t128_t1 = M_168 ;	// line#=../rle.cpp:77,78
	7'h67 :
		M_02_t128_t1 = M_98 ;	// line#=../rle.cpp:77,78
	7'h68 :
		M_02_t128_t1 = M_169 ;	// line#=../rle.cpp:77,78
	7'h69 :
		M_02_t128_t1 = M_99 ;	// line#=../rle.cpp:77,78
	7'h6a :
		M_02_t128_t1 = M_170 ;	// line#=../rle.cpp:77,78
	7'h6b :
		M_02_t128_t1 = M_100 ;	// line#=../rle.cpp:77,78
	7'h6c :
		M_02_t128_t1 = M_171 ;	// line#=../rle.cpp:77,78
	7'h6d :
		M_02_t128_t1 = M_102 ;	// line#=../rle.cpp:77,78
	7'h6e :
		M_02_t128_t1 = M_172 ;	// line#=../rle.cpp:77,78
	7'h6f :
		M_02_t128_t1 = M_103 ;	// line#=../rle.cpp:77,78
	7'h70 :
		M_02_t128_t1 = M_173 ;	// line#=../rle.cpp:77,78
	7'h71 :
		M_02_t128_t1 = M_104 ;	// line#=../rle.cpp:77,78
	7'h72 :
		M_02_t128_t1 = M_174 ;	// line#=../rle.cpp:77,78
	7'h73 :
		M_02_t128_t1 = M_105 ;	// line#=../rle.cpp:77,78
	7'h74 :
		M_02_t128_t1 = M_175 ;	// line#=../rle.cpp:77,78
	7'h75 :
		M_02_t128_t1 = M_106 ;	// line#=../rle.cpp:77,78
	7'h76 :
		M_02_t128_t1 = M_176 ;	// line#=../rle.cpp:77,78
	7'h77 :
		M_02_t128_t1 = M_107 ;	// line#=../rle.cpp:77,78
	7'h78 :
		M_02_t128_t1 = M_177 ;	// line#=../rle.cpp:77,78
	7'h79 :
		M_02_t128_t1 = M_108 ;	// line#=../rle.cpp:77,78
	7'h7a :
		M_02_t128_t1 = M_178 ;	// line#=../rle.cpp:77,78
	7'h7b :
		M_02_t128_t1 = M_109 ;	// line#=../rle.cpp:77,78
	7'h7c :
		M_02_t128_t1 = M_179 ;	// line#=../rle.cpp:77,78
	7'h7d :
		M_02_t128_t1 = M_110 ;	// line#=../rle.cpp:77,78
	7'h7e :
		M_02_t128_t1 = M_112 ;	// line#=../rle.cpp:77,78
	7'h7f :
		M_02_t128_t1 = M_113 ;	// line#=../rle.cpp:77,78
	default :
		M_02_t128_t1 = 1'hx ;
	endcase
always @ ( M_02_t128_t1 or M_14_t128 )	// line#=../rle.cpp:77,78
	M_02_t128 = ( { 1{ M_14_t128 } } & M_02_t128_t1 )	// line#=../rle.cpp:77,78
		 ;	// line#=../rle.cpp:77,78
always @ ( RG_zz_62 or RG_zz_61 or RG_zz_60 or RG_zz_59 or RG_zz_58 or RG_zz_57 or 
	RG_zz_56 or RG_zz_55 or RG_zz_54 or RG_zz_53 or RG_zz_52 or RG_zz_51 or 
	RG_zz_50 or RG_zz_49 or RG_zz_48 or RG_zz_47 or RG_zz_46 or RG_zz_45 or 
	RG_zz_44 or RG_zz_43 or RG_zz_42 or RG_zz_41 or RG_zz_40 or RG_zz_39 or 
	RG_zz_38 or RG_zz_37 or RG_zz_36 or RG_zz_35 or RG_zz_34 or RG_zz_33 or 
	RG_zz_32 or RG_zz_31 or RG_zz_30 or RG_zz_29 or RG_zz_28 or RG_zz_27 or 
	RG_zz_26 or RG_zz_25 or RG_zz_24 or RG_zz_23 or RG_zz_22 or RG_zz_21 or 
	RG_zz_20 or RG_zz_19 or RG_zz_18 or RG_zz_17 or RG_zz_16 or RG_zz_15 or 
	RG_zz_14 or RG_zz_13 or RG_zz_12 or RG_zz_11 or RG_zz_10 or RG_zz_9 or RG_zz_8 or 
	RG_zz_7 or RG_zz_6 or RG_zz_5 or RG_zz_4 or RG_zz_3 or RG_zz_2 or RG_zz_1 or 
	RG_zz or RG_quantized_block_rl_zz or RG_i_j_01 )	// line#=../rle.cpp:61,62
	case ( RG_i_j_01 [5:0] )
	6'h00 :
		M_01_t64_t1 = ~|RG_quantized_block_rl_zz ;	// line#=../rle.cpp:61,62
	6'h01 :
		M_01_t64_t1 = ~|RG_zz ;	// line#=../rle.cpp:61,62
	6'h02 :
		M_01_t64_t1 = ~|RG_zz_1 ;	// line#=../rle.cpp:61,62
	6'h03 :
		M_01_t64_t1 = ~|RG_zz_2 ;	// line#=../rle.cpp:61,62
	6'h04 :
		M_01_t64_t1 = ~|RG_zz_3 ;	// line#=../rle.cpp:61,62
	6'h05 :
		M_01_t64_t1 = ~|RG_zz_4 ;	// line#=../rle.cpp:61,62
	6'h06 :
		M_01_t64_t1 = ~|RG_zz_5 ;	// line#=../rle.cpp:61,62
	6'h07 :
		M_01_t64_t1 = ~|RG_zz_6 ;	// line#=../rle.cpp:61,62
	6'h08 :
		M_01_t64_t1 = ~|RG_zz_7 ;	// line#=../rle.cpp:61,62
	6'h09 :
		M_01_t64_t1 = ~|RG_zz_8 ;	// line#=../rle.cpp:61,62
	6'h0a :
		M_01_t64_t1 = ~|RG_zz_9 ;	// line#=../rle.cpp:61,62
	6'h0b :
		M_01_t64_t1 = ~|RG_zz_10 ;	// line#=../rle.cpp:61,62
	6'h0c :
		M_01_t64_t1 = ~|RG_zz_11 ;	// line#=../rle.cpp:61,62
	6'h0d :
		M_01_t64_t1 = ~|RG_zz_12 ;	// line#=../rle.cpp:61,62
	6'h0e :
		M_01_t64_t1 = ~|RG_zz_13 ;	// line#=../rle.cpp:61,62
	6'h0f :
		M_01_t64_t1 = ~|RG_zz_14 ;	// line#=../rle.cpp:61,62
	6'h10 :
		M_01_t64_t1 = ~|RG_zz_15 ;	// line#=../rle.cpp:61,62
	6'h11 :
		M_01_t64_t1 = ~|RG_zz_16 ;	// line#=../rle.cpp:61,62
	6'h12 :
		M_01_t64_t1 = ~|RG_zz_17 ;	// line#=../rle.cpp:61,62
	6'h13 :
		M_01_t64_t1 = ~|RG_zz_18 ;	// line#=../rle.cpp:61,62
	6'h14 :
		M_01_t64_t1 = ~|RG_zz_19 ;	// line#=../rle.cpp:61,62
	6'h15 :
		M_01_t64_t1 = ~|RG_zz_20 ;	// line#=../rle.cpp:61,62
	6'h16 :
		M_01_t64_t1 = ~|RG_zz_21 ;	// line#=../rle.cpp:61,62
	6'h17 :
		M_01_t64_t1 = ~|RG_zz_22 ;	// line#=../rle.cpp:61,62
	6'h18 :
		M_01_t64_t1 = ~|RG_zz_23 ;	// line#=../rle.cpp:61,62
	6'h19 :
		M_01_t64_t1 = ~|RG_zz_24 ;	// line#=../rle.cpp:61,62
	6'h1a :
		M_01_t64_t1 = ~|RG_zz_25 ;	// line#=../rle.cpp:61,62
	6'h1b :
		M_01_t64_t1 = ~|RG_zz_26 ;	// line#=../rle.cpp:61,62
	6'h1c :
		M_01_t64_t1 = ~|RG_zz_27 ;	// line#=../rle.cpp:61,62
	6'h1d :
		M_01_t64_t1 = ~|RG_zz_28 ;	// line#=../rle.cpp:61,62
	6'h1e :
		M_01_t64_t1 = ~|RG_zz_29 ;	// line#=../rle.cpp:61,62
	6'h1f :
		M_01_t64_t1 = ~|RG_zz_30 ;	// line#=../rle.cpp:61,62
	6'h20 :
		M_01_t64_t1 = ~|RG_zz_31 ;	// line#=../rle.cpp:61,62
	6'h21 :
		M_01_t64_t1 = ~|RG_zz_32 ;	// line#=../rle.cpp:61,62
	6'h22 :
		M_01_t64_t1 = ~|RG_zz_33 ;	// line#=../rle.cpp:61,62
	6'h23 :
		M_01_t64_t1 = ~|RG_zz_34 ;	// line#=../rle.cpp:61,62
	6'h24 :
		M_01_t64_t1 = ~|RG_zz_35 ;	// line#=../rle.cpp:61,62
	6'h25 :
		M_01_t64_t1 = ~|RG_zz_36 ;	// line#=../rle.cpp:61,62
	6'h26 :
		M_01_t64_t1 = ~|RG_zz_37 ;	// line#=../rle.cpp:61,62
	6'h27 :
		M_01_t64_t1 = ~|RG_zz_38 ;	// line#=../rle.cpp:61,62
	6'h28 :
		M_01_t64_t1 = ~|RG_zz_39 ;	// line#=../rle.cpp:61,62
	6'h29 :
		M_01_t64_t1 = ~|RG_zz_40 ;	// line#=../rle.cpp:61,62
	6'h2a :
		M_01_t64_t1 = ~|RG_zz_41 ;	// line#=../rle.cpp:61,62
	6'h2b :
		M_01_t64_t1 = ~|RG_zz_42 ;	// line#=../rle.cpp:61,62
	6'h2c :
		M_01_t64_t1 = ~|RG_zz_43 ;	// line#=../rle.cpp:61,62
	6'h2d :
		M_01_t64_t1 = ~|RG_zz_44 ;	// line#=../rle.cpp:61,62
	6'h2e :
		M_01_t64_t1 = ~|RG_zz_45 ;	// line#=../rle.cpp:61,62
	6'h2f :
		M_01_t64_t1 = ~|RG_zz_46 ;	// line#=../rle.cpp:61,62
	6'h30 :
		M_01_t64_t1 = ~|RG_zz_47 ;	// line#=../rle.cpp:61,62
	6'h31 :
		M_01_t64_t1 = ~|RG_zz_48 ;	// line#=../rle.cpp:61,62
	6'h32 :
		M_01_t64_t1 = ~|RG_zz_49 ;	// line#=../rle.cpp:61,62
	6'h33 :
		M_01_t64_t1 = ~|RG_zz_50 ;	// line#=../rle.cpp:61,62
	6'h34 :
		M_01_t64_t1 = ~|RG_zz_51 ;	// line#=../rle.cpp:61,62
	6'h35 :
		M_01_t64_t1 = ~|RG_zz_52 ;	// line#=../rle.cpp:61,62
	6'h36 :
		M_01_t64_t1 = ~|RG_zz_53 ;	// line#=../rle.cpp:61,62
	6'h37 :
		M_01_t64_t1 = ~|RG_zz_54 ;	// line#=../rle.cpp:61,62
	6'h38 :
		M_01_t64_t1 = ~|RG_zz_55 ;	// line#=../rle.cpp:61,62
	6'h39 :
		M_01_t64_t1 = ~|RG_zz_56 ;	// line#=../rle.cpp:61,62
	6'h3a :
		M_01_t64_t1 = ~|RG_zz_57 ;	// line#=../rle.cpp:61,62
	6'h3b :
		M_01_t64_t1 = ~|RG_zz_58 ;	// line#=../rle.cpp:61,62
	6'h3c :
		M_01_t64_t1 = ~|RG_zz_59 ;	// line#=../rle.cpp:61,62
	6'h3d :
		M_01_t64_t1 = ~|RG_zz_60 ;	// line#=../rle.cpp:61,62
	6'h3e :
		M_01_t64_t1 = ~|RG_zz_61 ;	// line#=../rle.cpp:61,62
	6'h3f :
		M_01_t64_t1 = ~|RG_zz_62 ;	// line#=../rle.cpp:61,62
	default :
		M_01_t64_t1 = 1'hx ;
	endcase
always @ ( M_01_t64_t1 or C_07 )	// line#=../rle.cpp:61,62
	M_01_t64 = ( { 1{ C_07 } } & M_01_t64_t1 )	// line#=../rle.cpp:61,62
		 ;	// line#=../rle.cpp:61,62
always @ ( RG_rl_127 or RG_rl_126 or RG_rl_125 or RG_rl_124 or RG_rl_123 or RG_rl_122 or 
	RG_rl_121 or RG_rl_120 or RG_rl_119 or RG_rl_118 or RG_rl_117 or RG_rl_116 or 
	RG_rl_115 or RG_rl_114 or RG_rl_113 or RG_rl_112 or RG_rl_111 or RG_rl_110 or 
	RG_rl_109 or RG_rl_108 or RG_rl_107 or RG_rl_106 or RG_rl_105 or RG_rl_104 or 
	RG_rl_103 or RG_rl_102 or RG_rl_101 or RG_rl_100 or RG_rl_99 or RG_rl_98 or 
	RG_rl_97 or RG_rl_96 or RG_rl_95 or RG_rl_94 or RG_rl_93 or RG_rl_92 or 
	RG_rl_91 or RG_rl_90 or RG_rl_89 or RG_rl_88 or RG_rl_87 or RG_rl_86 or 
	RG_rl_85 or RG_rl_84 or RG_rl_83 or RG_rl_82 or RG_rl_81 or RG_rl_80 or 
	RG_rl_79 or RG_rl_78 or RG_rl_77 or RG_rl_76 or RG_rl_75 or RG_rl_74 or 
	RG_rl_73 or RG_rl_72 or RG_rl_71 or RG_rl_70 or RG_rl_69 or RG_rl_68 or 
	RG_rl_67 or RG_rl_66 or RG_rl_65 or RG_rl_64 or RG_rl_63 or RG_rl_62 or 
	RG_rl_61 or RG_rl_60 or RG_rl_59 or RG_rl_58 or RG_rl_57 or RG_rl_56 or 
	RG_rl_55 or RG_rl_54 or RG_rl_53 or RG_rl_52 or RG_rl_51 or RG_rl_50 or 
	RG_rl_49 or RG_rl_48 or RG_rl_47 or RG_rl_46 or RG_rl_45 or RG_rl_44 or 
	RG_rl_43 or RG_rl_42 or RG_rl_41 or RG_rl_40 or RG_rl_39 or RG_rl_38 or 
	RG_rl_37 or RG_rl_36 or RG_rl_35 or RG_rl_34 or RG_rl_33 or RG_rl_32 or 
	RG_rl_31 or RG_rl_30 or RG_rl_29 or RG_rl_28 or RG_rl_27 or RG_rl_26 or 
	RG_rl_25 or RG_rl_24 or RG_rl_23 or RG_rl_22 or RG_rl_21 or RG_rl_20 or 
	RG_rl_19 or RG_rl_18 or RG_rl_17 or RG_rl_16 or RG_rl_15 or RG_rl_14 or 
	RG_rl_13 or RG_rl_12 or RG_rl_11 or RG_rl_10 or RG_rl_9 or RG_rl_8 or RG_rl_7 or 
	RG_rl_6 or RG_rl_5 or RG_rl_4 or RG_rl_3 or RG_rl_2 or RG_rl_1 or RG_rl or 
	sub8u_7_11ot )	// line#=../rle.cpp:83,84
	case ( sub8u_7_11ot )
	7'h00 :
		M_03_t128_t1 = ~|RG_rl ;	// line#=../rle.cpp:83,84
	7'h01 :
		M_03_t128_t1 = ~|RG_rl_1 ;	// line#=../rle.cpp:83,84
	7'h02 :
		M_03_t128_t1 = ~|RG_rl_2 ;	// line#=../rle.cpp:83,84
	7'h03 :
		M_03_t128_t1 = ~|RG_rl_3 ;	// line#=../rle.cpp:83,84
	7'h04 :
		M_03_t128_t1 = ~|RG_rl_4 ;	// line#=../rle.cpp:83,84
	7'h05 :
		M_03_t128_t1 = ~|RG_rl_5 ;	// line#=../rle.cpp:83,84
	7'h06 :
		M_03_t128_t1 = ~|RG_rl_6 ;	// line#=../rle.cpp:83,84
	7'h07 :
		M_03_t128_t1 = ~|RG_rl_7 ;	// line#=../rle.cpp:83,84
	7'h08 :
		M_03_t128_t1 = ~|RG_rl_8 ;	// line#=../rle.cpp:83,84
	7'h09 :
		M_03_t128_t1 = ~|RG_rl_9 ;	// line#=../rle.cpp:83,84
	7'h0a :
		M_03_t128_t1 = ~|RG_rl_10 ;	// line#=../rle.cpp:83,84
	7'h0b :
		M_03_t128_t1 = ~|RG_rl_11 ;	// line#=../rle.cpp:83,84
	7'h0c :
		M_03_t128_t1 = ~|RG_rl_12 ;	// line#=../rle.cpp:83,84
	7'h0d :
		M_03_t128_t1 = ~|RG_rl_13 ;	// line#=../rle.cpp:83,84
	7'h0e :
		M_03_t128_t1 = ~|RG_rl_14 ;	// line#=../rle.cpp:83,84
	7'h0f :
		M_03_t128_t1 = ~|RG_rl_15 ;	// line#=../rle.cpp:83,84
	7'h10 :
		M_03_t128_t1 = ~|RG_rl_16 ;	// line#=../rle.cpp:83,84
	7'h11 :
		M_03_t128_t1 = ~|RG_rl_17 ;	// line#=../rle.cpp:83,84
	7'h12 :
		M_03_t128_t1 = ~|RG_rl_18 ;	// line#=../rle.cpp:83,84
	7'h13 :
		M_03_t128_t1 = ~|RG_rl_19 ;	// line#=../rle.cpp:83,84
	7'h14 :
		M_03_t128_t1 = ~|RG_rl_20 ;	// line#=../rle.cpp:83,84
	7'h15 :
		M_03_t128_t1 = ~|RG_rl_21 ;	// line#=../rle.cpp:83,84
	7'h16 :
		M_03_t128_t1 = ~|RG_rl_22 ;	// line#=../rle.cpp:83,84
	7'h17 :
		M_03_t128_t1 = ~|RG_rl_23 ;	// line#=../rle.cpp:83,84
	7'h18 :
		M_03_t128_t1 = ~|RG_rl_24 ;	// line#=../rle.cpp:83,84
	7'h19 :
		M_03_t128_t1 = ~|RG_rl_25 ;	// line#=../rle.cpp:83,84
	7'h1a :
		M_03_t128_t1 = ~|RG_rl_26 ;	// line#=../rle.cpp:83,84
	7'h1b :
		M_03_t128_t1 = ~|RG_rl_27 ;	// line#=../rle.cpp:83,84
	7'h1c :
		M_03_t128_t1 = ~|RG_rl_28 ;	// line#=../rle.cpp:83,84
	7'h1d :
		M_03_t128_t1 = ~|RG_rl_29 ;	// line#=../rle.cpp:83,84
	7'h1e :
		M_03_t128_t1 = ~|RG_rl_30 ;	// line#=../rle.cpp:83,84
	7'h1f :
		M_03_t128_t1 = ~|RG_rl_31 ;	// line#=../rle.cpp:83,84
	7'h20 :
		M_03_t128_t1 = ~|RG_rl_32 ;	// line#=../rle.cpp:83,84
	7'h21 :
		M_03_t128_t1 = ~|RG_rl_33 ;	// line#=../rle.cpp:83,84
	7'h22 :
		M_03_t128_t1 = ~|RG_rl_34 ;	// line#=../rle.cpp:83,84
	7'h23 :
		M_03_t128_t1 = ~|RG_rl_35 ;	// line#=../rle.cpp:83,84
	7'h24 :
		M_03_t128_t1 = ~|RG_rl_36 ;	// line#=../rle.cpp:83,84
	7'h25 :
		M_03_t128_t1 = ~|RG_rl_37 ;	// line#=../rle.cpp:83,84
	7'h26 :
		M_03_t128_t1 = ~|RG_rl_38 ;	// line#=../rle.cpp:83,84
	7'h27 :
		M_03_t128_t1 = ~|RG_rl_39 ;	// line#=../rle.cpp:83,84
	7'h28 :
		M_03_t128_t1 = ~|RG_rl_40 ;	// line#=../rle.cpp:83,84
	7'h29 :
		M_03_t128_t1 = ~|RG_rl_41 ;	// line#=../rle.cpp:83,84
	7'h2a :
		M_03_t128_t1 = ~|RG_rl_42 ;	// line#=../rle.cpp:83,84
	7'h2b :
		M_03_t128_t1 = ~|RG_rl_43 ;	// line#=../rle.cpp:83,84
	7'h2c :
		M_03_t128_t1 = ~|RG_rl_44 ;	// line#=../rle.cpp:83,84
	7'h2d :
		M_03_t128_t1 = ~|RG_rl_45 ;	// line#=../rle.cpp:83,84
	7'h2e :
		M_03_t128_t1 = ~|RG_rl_46 ;	// line#=../rle.cpp:83,84
	7'h2f :
		M_03_t128_t1 = ~|RG_rl_47 ;	// line#=../rle.cpp:83,84
	7'h30 :
		M_03_t128_t1 = ~|RG_rl_48 ;	// line#=../rle.cpp:83,84
	7'h31 :
		M_03_t128_t1 = ~|RG_rl_49 ;	// line#=../rle.cpp:83,84
	7'h32 :
		M_03_t128_t1 = ~|RG_rl_50 ;	// line#=../rle.cpp:83,84
	7'h33 :
		M_03_t128_t1 = ~|RG_rl_51 ;	// line#=../rle.cpp:83,84
	7'h34 :
		M_03_t128_t1 = ~|RG_rl_52 ;	// line#=../rle.cpp:83,84
	7'h35 :
		M_03_t128_t1 = ~|RG_rl_53 ;	// line#=../rle.cpp:83,84
	7'h36 :
		M_03_t128_t1 = ~|RG_rl_54 ;	// line#=../rle.cpp:83,84
	7'h37 :
		M_03_t128_t1 = ~|RG_rl_55 ;	// line#=../rle.cpp:83,84
	7'h38 :
		M_03_t128_t1 = ~|RG_rl_56 ;	// line#=../rle.cpp:83,84
	7'h39 :
		M_03_t128_t1 = ~|RG_rl_57 ;	// line#=../rle.cpp:83,84
	7'h3a :
		M_03_t128_t1 = ~|RG_rl_58 ;	// line#=../rle.cpp:83,84
	7'h3b :
		M_03_t128_t1 = ~|RG_rl_59 ;	// line#=../rle.cpp:83,84
	7'h3c :
		M_03_t128_t1 = ~|RG_rl_60 ;	// line#=../rle.cpp:83,84
	7'h3d :
		M_03_t128_t1 = ~|RG_rl_61 ;	// line#=../rle.cpp:83,84
	7'h3e :
		M_03_t128_t1 = ~|RG_rl_62 ;	// line#=../rle.cpp:83,84
	7'h3f :
		M_03_t128_t1 = ~|RG_rl_63 ;	// line#=../rle.cpp:83,84
	7'h40 :
		M_03_t128_t1 = ~|RG_rl_64 ;	// line#=../rle.cpp:83,84
	7'h41 :
		M_03_t128_t1 = ~|RG_rl_65 ;	// line#=../rle.cpp:83,84
	7'h42 :
		M_03_t128_t1 = ~|RG_rl_66 ;	// line#=../rle.cpp:83,84
	7'h43 :
		M_03_t128_t1 = ~|RG_rl_67 ;	// line#=../rle.cpp:83,84
	7'h44 :
		M_03_t128_t1 = ~|RG_rl_68 ;	// line#=../rle.cpp:83,84
	7'h45 :
		M_03_t128_t1 = ~|RG_rl_69 ;	// line#=../rle.cpp:83,84
	7'h46 :
		M_03_t128_t1 = ~|RG_rl_70 ;	// line#=../rle.cpp:83,84
	7'h47 :
		M_03_t128_t1 = ~|RG_rl_71 ;	// line#=../rle.cpp:83,84
	7'h48 :
		M_03_t128_t1 = ~|RG_rl_72 ;	// line#=../rle.cpp:83,84
	7'h49 :
		M_03_t128_t1 = ~|RG_rl_73 ;	// line#=../rle.cpp:83,84
	7'h4a :
		M_03_t128_t1 = ~|RG_rl_74 ;	// line#=../rle.cpp:83,84
	7'h4b :
		M_03_t128_t1 = ~|RG_rl_75 ;	// line#=../rle.cpp:83,84
	7'h4c :
		M_03_t128_t1 = ~|RG_rl_76 ;	// line#=../rle.cpp:83,84
	7'h4d :
		M_03_t128_t1 = ~|RG_rl_77 ;	// line#=../rle.cpp:83,84
	7'h4e :
		M_03_t128_t1 = ~|RG_rl_78 ;	// line#=../rle.cpp:83,84
	7'h4f :
		M_03_t128_t1 = ~|RG_rl_79 ;	// line#=../rle.cpp:83,84
	7'h50 :
		M_03_t128_t1 = ~|RG_rl_80 ;	// line#=../rle.cpp:83,84
	7'h51 :
		M_03_t128_t1 = ~|RG_rl_81 ;	// line#=../rle.cpp:83,84
	7'h52 :
		M_03_t128_t1 = ~|RG_rl_82 ;	// line#=../rle.cpp:83,84
	7'h53 :
		M_03_t128_t1 = ~|RG_rl_83 ;	// line#=../rle.cpp:83,84
	7'h54 :
		M_03_t128_t1 = ~|RG_rl_84 ;	// line#=../rle.cpp:83,84
	7'h55 :
		M_03_t128_t1 = ~|RG_rl_85 ;	// line#=../rle.cpp:83,84
	7'h56 :
		M_03_t128_t1 = ~|RG_rl_86 ;	// line#=../rle.cpp:83,84
	7'h57 :
		M_03_t128_t1 = ~|RG_rl_87 ;	// line#=../rle.cpp:83,84
	7'h58 :
		M_03_t128_t1 = ~|RG_rl_88 ;	// line#=../rle.cpp:83,84
	7'h59 :
		M_03_t128_t1 = ~|RG_rl_89 ;	// line#=../rle.cpp:83,84
	7'h5a :
		M_03_t128_t1 = ~|RG_rl_90 ;	// line#=../rle.cpp:83,84
	7'h5b :
		M_03_t128_t1 = ~|RG_rl_91 ;	// line#=../rle.cpp:83,84
	7'h5c :
		M_03_t128_t1 = ~|RG_rl_92 ;	// line#=../rle.cpp:83,84
	7'h5d :
		M_03_t128_t1 = ~|RG_rl_93 ;	// line#=../rle.cpp:83,84
	7'h5e :
		M_03_t128_t1 = ~|RG_rl_94 ;	// line#=../rle.cpp:83,84
	7'h5f :
		M_03_t128_t1 = ~|RG_rl_95 ;	// line#=../rle.cpp:83,84
	7'h60 :
		M_03_t128_t1 = ~|RG_rl_96 ;	// line#=../rle.cpp:83,84
	7'h61 :
		M_03_t128_t1 = ~|RG_rl_97 ;	// line#=../rle.cpp:83,84
	7'h62 :
		M_03_t128_t1 = ~|RG_rl_98 ;	// line#=../rle.cpp:83,84
	7'h63 :
		M_03_t128_t1 = ~|RG_rl_99 ;	// line#=../rle.cpp:83,84
	7'h64 :
		M_03_t128_t1 = ~|RG_rl_100 ;	// line#=../rle.cpp:83,84
	7'h65 :
		M_03_t128_t1 = ~|RG_rl_101 ;	// line#=../rle.cpp:83,84
	7'h66 :
		M_03_t128_t1 = ~|RG_rl_102 ;	// line#=../rle.cpp:83,84
	7'h67 :
		M_03_t128_t1 = ~|RG_rl_103 ;	// line#=../rle.cpp:83,84
	7'h68 :
		M_03_t128_t1 = ~|RG_rl_104 ;	// line#=../rle.cpp:83,84
	7'h69 :
		M_03_t128_t1 = ~|RG_rl_105 ;	// line#=../rle.cpp:83,84
	7'h6a :
		M_03_t128_t1 = ~|RG_rl_106 ;	// line#=../rle.cpp:83,84
	7'h6b :
		M_03_t128_t1 = ~|RG_rl_107 ;	// line#=../rle.cpp:83,84
	7'h6c :
		M_03_t128_t1 = ~|RG_rl_108 ;	// line#=../rle.cpp:83,84
	7'h6d :
		M_03_t128_t1 = ~|RG_rl_109 ;	// line#=../rle.cpp:83,84
	7'h6e :
		M_03_t128_t1 = ~|RG_rl_110 ;	// line#=../rle.cpp:83,84
	7'h6f :
		M_03_t128_t1 = ~|RG_rl_111 ;	// line#=../rle.cpp:83,84
	7'h70 :
		M_03_t128_t1 = ~|RG_rl_112 ;	// line#=../rle.cpp:83,84
	7'h71 :
		M_03_t128_t1 = ~|RG_rl_113 ;	// line#=../rle.cpp:83,84
	7'h72 :
		M_03_t128_t1 = ~|RG_rl_114 ;	// line#=../rle.cpp:83,84
	7'h73 :
		M_03_t128_t1 = ~|RG_rl_115 ;	// line#=../rle.cpp:83,84
	7'h74 :
		M_03_t128_t1 = ~|RG_rl_116 ;	// line#=../rle.cpp:83,84
	7'h75 :
		M_03_t128_t1 = ~|RG_rl_117 ;	// line#=../rle.cpp:83,84
	7'h76 :
		M_03_t128_t1 = ~|RG_rl_118 ;	// line#=../rle.cpp:83,84
	7'h77 :
		M_03_t128_t1 = ~|RG_rl_119 ;	// line#=../rle.cpp:83,84
	7'h78 :
		M_03_t128_t1 = ~|RG_rl_120 ;	// line#=../rle.cpp:83,84
	7'h79 :
		M_03_t128_t1 = ~|RG_rl_121 ;	// line#=../rle.cpp:83,84
	7'h7a :
		M_03_t128_t1 = ~|RG_rl_122 ;	// line#=../rle.cpp:83,84
	7'h7b :
		M_03_t128_t1 = ~|RG_rl_123 ;	// line#=../rle.cpp:83,84
	7'h7c :
		M_03_t128_t1 = ~|RG_rl_124 ;	// line#=../rle.cpp:83,84
	7'h7d :
		M_03_t128_t1 = ~|RG_rl_125 ;	// line#=../rle.cpp:83,84
	7'h7e :
		M_03_t128_t1 = ~|RG_rl_126 ;	// line#=../rle.cpp:83,84
	7'h7f :
		M_03_t128_t1 = ~|RG_rl_127 ;	// line#=../rle.cpp:83,84
	default :
		M_03_t128_t1 = 1'hx ;
	endcase
always @ ( M_03_t128_t1 or M_15_t128 )	// line#=../rle.cpp:83,84
	M_03_t128 = ( { 1{ M_15_t128 } } & M_03_t128_t1 )	// line#=../rle.cpp:83,84
		 ;	// line#=../rle.cpp:83,84
assign	JF_06 = ~M_03_t128 ;
assign	jpeg_out_a00_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a00_r_en )
		jpeg_out_a00_r <= RG_rl ;
assign	jpeg_out_a01_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a01_r_en )
		jpeg_out_a01_r <= RG_rl_1 ;
assign	jpeg_out_a02_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a02_r_en )
		jpeg_out_a02_r <= RG_rl_2 ;
assign	jpeg_out_a03_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a03_r_en )
		jpeg_out_a03_r <= RG_rl_3 ;
assign	jpeg_out_a04_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a04_r_en )
		jpeg_out_a04_r <= RG_rl_4 ;
assign	jpeg_out_a05_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a05_r_en )
		jpeg_out_a05_r <= RG_rl_5 ;
assign	jpeg_out_a06_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a06_r_en )
		jpeg_out_a06_r <= RG_rl_6 ;
assign	jpeg_out_a07_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a07_r_en )
		jpeg_out_a07_r <= RG_rl_7 ;
assign	jpeg_out_a08_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a08_r_en )
		jpeg_out_a08_r <= RG_rl_8 ;
assign	jpeg_out_a09_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a09_r_en )
		jpeg_out_a09_r <= RG_rl_9 ;
assign	jpeg_out_a10_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a10_r_en )
		jpeg_out_a10_r <= RG_rl_10 ;
assign	jpeg_out_a11_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a11_r_en )
		jpeg_out_a11_r <= RG_rl_11 ;
assign	jpeg_out_a12_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a12_r_en )
		jpeg_out_a12_r <= RG_rl_12 ;
assign	jpeg_out_a13_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a13_r_en )
		jpeg_out_a13_r <= RG_rl_13 ;
assign	jpeg_out_a14_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a14_r_en )
		jpeg_out_a14_r <= RG_rl_14 ;
assign	jpeg_out_a15_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a15_r_en )
		jpeg_out_a15_r <= RG_rl_15 ;
assign	jpeg_out_a16_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a16_r_en )
		jpeg_out_a16_r <= RG_rl_16 ;
assign	jpeg_out_a17_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a17_r_en )
		jpeg_out_a17_r <= RG_rl_17 ;
assign	jpeg_out_a18_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a18_r_en )
		jpeg_out_a18_r <= RG_rl_18 ;
assign	jpeg_out_a19_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a19_r_en )
		jpeg_out_a19_r <= RG_rl_19 ;
assign	jpeg_out_a20_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a20_r_en )
		jpeg_out_a20_r <= RG_rl_20 ;
assign	jpeg_out_a21_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a21_r_en )
		jpeg_out_a21_r <= RG_rl_21 ;
assign	jpeg_out_a22_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a22_r_en )
		jpeg_out_a22_r <= RG_rl_22 ;
assign	jpeg_out_a23_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a23_r_en )
		jpeg_out_a23_r <= RG_rl_23 ;
assign	jpeg_out_a24_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a24_r_en )
		jpeg_out_a24_r <= RG_rl_24 ;
assign	jpeg_out_a25_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a25_r_en )
		jpeg_out_a25_r <= RG_rl_25 ;
assign	jpeg_out_a26_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a26_r_en )
		jpeg_out_a26_r <= RG_rl_26 ;
assign	jpeg_out_a27_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a27_r_en )
		jpeg_out_a27_r <= RG_rl_27 ;
assign	jpeg_out_a28_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a28_r_en )
		jpeg_out_a28_r <= RG_rl_28 ;
assign	jpeg_out_a29_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a29_r_en )
		jpeg_out_a29_r <= RG_rl_29 ;
assign	jpeg_out_a30_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a30_r_en )
		jpeg_out_a30_r <= RG_rl_30 ;
assign	jpeg_out_a31_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a31_r_en )
		jpeg_out_a31_r <= RG_rl_31 ;
assign	jpeg_out_a32_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a32_r_en )
		jpeg_out_a32_r <= RG_rl_32 ;
assign	jpeg_out_a33_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a33_r_en )
		jpeg_out_a33_r <= RG_rl_33 ;
assign	jpeg_out_a34_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a34_r_en )
		jpeg_out_a34_r <= RG_rl_34 ;
assign	jpeg_out_a35_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a35_r_en )
		jpeg_out_a35_r <= RG_rl_35 ;
assign	jpeg_out_a36_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a36_r_en )
		jpeg_out_a36_r <= RG_rl_36 ;
assign	jpeg_out_a37_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a37_r_en )
		jpeg_out_a37_r <= RG_rl_37 ;
assign	jpeg_out_a38_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a38_r_en )
		jpeg_out_a38_r <= RG_rl_38 ;
assign	jpeg_out_a39_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a39_r_en )
		jpeg_out_a39_r <= RG_rl_39 ;
assign	jpeg_out_a40_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a40_r_en )
		jpeg_out_a40_r <= RG_rl_40 ;
assign	jpeg_out_a41_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a41_r_en )
		jpeg_out_a41_r <= RG_rl_41 ;
assign	jpeg_out_a42_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a42_r_en )
		jpeg_out_a42_r <= RG_rl_42 ;
assign	jpeg_out_a43_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a43_r_en )
		jpeg_out_a43_r <= RG_rl_43 ;
assign	jpeg_out_a44_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a44_r_en )
		jpeg_out_a44_r <= RG_rl_44 ;
assign	jpeg_out_a45_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a45_r_en )
		jpeg_out_a45_r <= RG_rl_45 ;
assign	jpeg_out_a46_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a46_r_en )
		jpeg_out_a46_r <= RG_rl_46 ;
assign	jpeg_out_a47_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a47_r_en )
		jpeg_out_a47_r <= RG_rl_47 ;
assign	jpeg_out_a48_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a48_r_en )
		jpeg_out_a48_r <= RG_rl_48 ;
assign	jpeg_out_a49_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a49_r_en )
		jpeg_out_a49_r <= RG_rl_49 ;
assign	jpeg_out_a50_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a50_r_en )
		jpeg_out_a50_r <= RG_rl_50 ;
assign	jpeg_out_a51_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a51_r_en )
		jpeg_out_a51_r <= RG_rl_51 ;
assign	jpeg_out_a52_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a52_r_en )
		jpeg_out_a52_r <= RG_rl_52 ;
assign	jpeg_out_a53_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a53_r_en )
		jpeg_out_a53_r <= RG_rl_53 ;
assign	jpeg_out_a54_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a54_r_en )
		jpeg_out_a54_r <= RG_rl_54 ;
assign	jpeg_out_a55_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a55_r_en )
		jpeg_out_a55_r <= RG_rl_55 ;
assign	jpeg_out_a56_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a56_r_en )
		jpeg_out_a56_r <= RG_rl_56 ;
assign	jpeg_out_a57_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a57_r_en )
		jpeg_out_a57_r <= RG_rl_57 ;
assign	jpeg_out_a58_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a58_r_en )
		jpeg_out_a58_r <= RG_rl_58 ;
assign	jpeg_out_a59_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a59_r_en )
		jpeg_out_a59_r <= RG_rl_59 ;
assign	jpeg_out_a60_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a60_r_en )
		jpeg_out_a60_r <= RG_rl_60 ;
assign	jpeg_out_a61_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a61_r_en )
		jpeg_out_a61_r <= RG_rl_61 ;
assign	jpeg_out_a62_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a62_r_en )
		jpeg_out_a62_r <= RG_rl_62 ;
assign	jpeg_out_a63_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a63_r_en )
		jpeg_out_a63_r <= RG_rl_63 ;
assign	jpeg_out_a64_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a64_r_en )
		jpeg_out_a64_r <= RG_rl_64 ;
assign	jpeg_out_a65_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a65_r_en )
		jpeg_out_a65_r <= RG_rl_65 ;
assign	jpeg_out_a66_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a66_r_en )
		jpeg_out_a66_r <= RG_rl_66 ;
assign	jpeg_out_a67_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a67_r_en )
		jpeg_out_a67_r <= RG_rl_67 ;
assign	jpeg_out_a68_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a68_r_en )
		jpeg_out_a68_r <= RG_rl_68 ;
assign	jpeg_out_a69_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a69_r_en )
		jpeg_out_a69_r <= RG_rl_69 ;
assign	jpeg_out_a70_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a70_r_en )
		jpeg_out_a70_r <= RG_rl_70 ;
assign	jpeg_out_a71_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a71_r_en )
		jpeg_out_a71_r <= RG_rl_71 ;
assign	jpeg_out_a72_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a72_r_en )
		jpeg_out_a72_r <= RG_rl_72 ;
assign	jpeg_out_a73_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a73_r_en )
		jpeg_out_a73_r <= RG_rl_73 ;
assign	jpeg_out_a74_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a74_r_en )
		jpeg_out_a74_r <= RG_rl_74 ;
assign	jpeg_out_a75_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a75_r_en )
		jpeg_out_a75_r <= RG_rl_75 ;
assign	jpeg_out_a76_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a76_r_en )
		jpeg_out_a76_r <= RG_rl_76 ;
assign	jpeg_out_a77_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a77_r_en )
		jpeg_out_a77_r <= RG_rl_77 ;
assign	jpeg_out_a78_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a78_r_en )
		jpeg_out_a78_r <= RG_rl_78 ;
assign	jpeg_out_a79_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a79_r_en )
		jpeg_out_a79_r <= RG_rl_79 ;
assign	jpeg_out_a80_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a80_r_en )
		jpeg_out_a80_r <= RG_rl_80 ;
assign	jpeg_out_a81_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a81_r_en )
		jpeg_out_a81_r <= RG_rl_81 ;
assign	jpeg_out_a82_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a82_r_en )
		jpeg_out_a82_r <= RG_rl_82 ;
assign	jpeg_out_a83_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a83_r_en )
		jpeg_out_a83_r <= RG_rl_83 ;
assign	jpeg_out_a84_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a84_r_en )
		jpeg_out_a84_r <= RG_rl_84 ;
assign	jpeg_out_a85_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a85_r_en )
		jpeg_out_a85_r <= RG_rl_85 ;
assign	jpeg_out_a86_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a86_r_en )
		jpeg_out_a86_r <= RG_rl_86 ;
assign	jpeg_out_a87_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a87_r_en )
		jpeg_out_a87_r <= RG_rl_87 ;
assign	jpeg_out_a88_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a88_r_en )
		jpeg_out_a88_r <= RG_rl_88 ;
assign	jpeg_out_a89_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a89_r_en )
		jpeg_out_a89_r <= RG_rl_89 ;
assign	jpeg_out_a90_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a90_r_en )
		jpeg_out_a90_r <= RG_rl_90 ;
assign	jpeg_out_a91_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a91_r_en )
		jpeg_out_a91_r <= RG_rl_91 ;
assign	jpeg_out_a92_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a92_r_en )
		jpeg_out_a92_r <= RG_rl_92 ;
assign	jpeg_out_a93_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a93_r_en )
		jpeg_out_a93_r <= RG_rl_93 ;
assign	jpeg_out_a94_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a94_r_en )
		jpeg_out_a94_r <= RG_rl_94 ;
assign	jpeg_out_a95_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a95_r_en )
		jpeg_out_a95_r <= RG_rl_95 ;
assign	jpeg_out_a96_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a96_r_en )
		jpeg_out_a96_r <= RG_rl_96 ;
assign	jpeg_out_a97_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a97_r_en )
		jpeg_out_a97_r <= RG_rl_97 ;
assign	jpeg_out_a98_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a98_r_en )
		jpeg_out_a98_r <= RG_rl_98 ;
assign	jpeg_out_a99_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a99_r_en )
		jpeg_out_a99_r <= RG_rl_99 ;
assign	jpeg_out_a100_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a100_r_en )
		jpeg_out_a100_r <= RG_rl_100 ;
assign	jpeg_out_a101_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a101_r_en )
		jpeg_out_a101_r <= RG_rl_101 ;
assign	jpeg_out_a102_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a102_r_en )
		jpeg_out_a102_r <= RG_rl_102 ;
assign	jpeg_out_a103_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a103_r_en )
		jpeg_out_a103_r <= RG_rl_103 ;
assign	jpeg_out_a104_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a104_r_en )
		jpeg_out_a104_r <= RG_rl_104 ;
assign	jpeg_out_a105_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a105_r_en )
		jpeg_out_a105_r <= RG_rl_105 ;
assign	jpeg_out_a106_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a106_r_en )
		jpeg_out_a106_r <= RG_rl_106 ;
assign	jpeg_out_a107_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a107_r_en )
		jpeg_out_a107_r <= RG_rl_107 ;
assign	jpeg_out_a108_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a108_r_en )
		jpeg_out_a108_r <= RG_rl_108 ;
assign	jpeg_out_a109_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a109_r_en )
		jpeg_out_a109_r <= RG_rl_109 ;
assign	jpeg_out_a110_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a110_r_en )
		jpeg_out_a110_r <= RG_rl_110 ;
assign	jpeg_out_a111_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a111_r_en )
		jpeg_out_a111_r <= RG_rl_111 ;
assign	jpeg_out_a112_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a112_r_en )
		jpeg_out_a112_r <= RG_rl_112 ;
assign	jpeg_out_a113_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a113_r_en )
		jpeg_out_a113_r <= RG_rl_113 ;
assign	jpeg_out_a114_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a114_r_en )
		jpeg_out_a114_r <= RG_rl_114 ;
assign	jpeg_out_a115_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a115_r_en )
		jpeg_out_a115_r <= RG_rl_115 ;
assign	jpeg_out_a116_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a116_r_en )
		jpeg_out_a116_r <= RG_rl_116 ;
assign	jpeg_out_a117_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a117_r_en )
		jpeg_out_a117_r <= RG_rl_117 ;
assign	jpeg_out_a118_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a118_r_en )
		jpeg_out_a118_r <= RG_rl_118 ;
assign	jpeg_out_a119_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a119_r_en )
		jpeg_out_a119_r <= RG_rl_119 ;
assign	jpeg_out_a120_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a120_r_en )
		jpeg_out_a120_r <= RG_rl_120 ;
assign	jpeg_out_a121_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a121_r_en )
		jpeg_out_a121_r <= RG_rl_121 ;
assign	jpeg_out_a122_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a122_r_en )
		jpeg_out_a122_r <= RG_rl_122 ;
assign	jpeg_out_a123_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a123_r_en )
		jpeg_out_a123_r <= RG_rl_123 ;
assign	jpeg_out_a124_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a124_r_en )
		jpeg_out_a124_r <= RG_rl_124 ;
assign	jpeg_out_a125_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a125_r_en )
		jpeg_out_a125_r <= RG_rl_125 ;
assign	jpeg_out_a126_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a126_r_en )
		jpeg_out_a126_r <= RG_rl_126 ;
assign	jpeg_out_a127_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a127_r_en )
		jpeg_out_a127_r <= RG_rl_127 ;
assign	jpeg_len_out_r_en = U_184 ;
always @ ( posedge clk )	// line#=../rle.cpp:93
	if ( jpeg_len_out_r_en )
		jpeg_len_out_r <= { 4'h0 , RG_len_1 } ;
always @ ( U_184 )
	valid_r_t = ( { 1{ U_184 } } & 1'h1 )	// line#=../rle.cpp:95
		 ;	// line#=../rle.cpp:30
assign	valid_r_en = ( ST1_01d | U_184 ) ;
always @ ( posedge clk )
	if ( valid_r_en )
		valid_r <= valid_r_t ;	// line#=../rle.cpp:30,95
assign	incr8u1i1 = RG_len ;	// line#=../rle.cpp:68,79
always @ ( RG_k_1 or U_87 or RG_k or U_05 )
	TR_03 = ( ( { 6{ U_05 } } & RG_k )		// line#=../rle.cpp:111
		| ( { 6{ U_87 } } & RG_k_1 [5:0] )	// line#=../rle.cpp:142
		) ;
always @ ( TR_03 or U_87 or U_05 or incr8u2ot or U_318 )
	begin
	incr8u3i1_c1 = ( U_05 | U_87 ) ;	// line#=../rle.cpp:111,142
	incr8u3i1 = ( ( { 8{ U_318 } } & incr8u2ot )		// line#=../rle.cpp:73,74
		| ( { 8{ incr8u3i1_c1 } } & { 2'h0 , TR_03 } )	// line#=../rle.cpp:111,142
		) ;
	end
assign	incr8u4i1 = incr8u1ot ;	// line#=../rle.cpp:68,69,79,80
assign	incr32s1i1 = RG_i_j_01 ;	// line#=../rle.cpp:61,62,63,74,114,125
					// ,145,156
assign	incr32s2i1 = RG_i_k_01 ;	// line#=../rle.cpp:61,62,64,119,129,150
					// ,160
assign	decr32s1i1 = RG_i_k_01 ;	// line#=../rle.cpp:124,155
assign	decr32s2i1 = RG_i_j_01 ;	// line#=../rle.cpp:130,161
always @ ( RG_len_1 or ST1_07d or RG_len or ST1_05d )
	sub8u_7_11i1 = ( ( { 7{ ST1_05d } } & RG_len [6:0] )	// line#=../rle.cpp:77,78
		| ( { 7{ ST1_07d } } & RG_len_1 [6:0] )		// line#=../rle.cpp:83,84
		) ;
assign	sub8u_7_11i2 = { 1'h1 , ST1_07d } ;	// line#=../rle.cpp:77,78,83,84

endmodule

module jpeg_sub8u_7_1 ( i1 ,i2 ,o1 );
input	[6:0]	i1 ;
input	[1:0]	i2 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - { 5'h00 , i2 } ) ;

endmodule

module jpeg_sub8u_7 ( i1 ,i2 ,o1 );
input	[6:0]	i1 ;
input	[2:0]	i2 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - { 4'h0 , i2 } ) ;

endmodule

module jpeg_decr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_decr8u_7 ( i1 ,o1 );
input	[6:0]	i1 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_incr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr8u ( i1 ,o1 );
input	[7:0]	i1 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr4s ( i1 ,o1 );
input	[3:0]	i1 ;
output	[3:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_lop8u_1 ( i1 ,i2 ,o1 );
input	[5:0]	i1 ;
input	[5:0]	i2 ;
output		o1 ;
wire		M_01 ;

assign	M_01 = ( i1 < i2 ) ;
assign	o1 = M_01 ;

endmodule

module jpeg_sub12s_9 ( i1 ,i2 ,o1 );
input	[8:0]	i1 ;
input	[8:0]	i2 ;
output	[8:0]	o1 ;

assign	o1 = ( i1 - i2 ) ;

endmodule

module jpeg_sub8u ( i1 ,i2 ,o1 );
input	[7:0]	i1 ;
input	[1:0]	i2 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 - { 6'h00 , i2 } ) ;

endmodule
