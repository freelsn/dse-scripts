// verilog_out version 6.79.2
// options:  veriloggen jpeg_E.IFF
// bdlpars options:  -DDSE ../rle.cpp
// bdltran options:  -c1000 -s -Zresource_fcnt=GENERATE -Zresource_mcnt=GENERATE -lb /home/shuangnan/share/packages/zynq-1.BLIB -lfl /home/shuangnan/share/packages/zynq-1.FLIB jpeg.IFF -OX -a8196 -Zfu_cnt_incr_rate=0 -tcio 
// timestamp_0: 20180213182124_01267_91723
// timestamp_5: 20180213182128_02690_60421
// timestamp_9: 20180213182135_02690_27152
// timestamp_C: 20180213182134_02690_06731
// timestamp_E: 20180213182135_02690_97865
// timestamp_V: 20180213182138_04883_47886

module jpeg ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,jpeg_in_a04 ,
	jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,jpeg_in_a10 ,
	jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,jpeg_in_a16 ,
	jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,jpeg_in_a22 ,
	jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,jpeg_in_a28 ,
	jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,jpeg_in_a34 ,
	jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,jpeg_in_a40 ,
	jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,jpeg_in_a46 ,
	jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,jpeg_in_a52 ,
	jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,jpeg_in_a58 ,
	jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,jpeg_in_a64 ,
	jpeg_in_a65 ,jpeg_in_a66 ,jpeg_in_a67 ,jpeg_in_a68 ,jpeg_in_a69 ,jpeg_in_a70 ,
	jpeg_in_a71 ,jpeg_in_a72 ,jpeg_in_a73 ,jpeg_in_a74 ,jpeg_in_a75 ,jpeg_in_a76 ,
	jpeg_in_a77 ,jpeg_in_a78 ,jpeg_in_a79 ,jpeg_in_a80 ,jpeg_in_a81 ,jpeg_in_a82 ,
	jpeg_in_a83 ,jpeg_in_a84 ,jpeg_in_a85 ,jpeg_in_a86 ,jpeg_in_a87 ,jpeg_in_a88 ,
	jpeg_in_a89 ,jpeg_in_a90 ,jpeg_in_a91 ,jpeg_in_a92 ,jpeg_in_a93 ,jpeg_in_a94 ,
	jpeg_in_a95 ,jpeg_in_a96 ,jpeg_in_a97 ,jpeg_in_a98 ,jpeg_in_a99 ,jpeg_in_a100 ,
	jpeg_in_a101 ,jpeg_in_a102 ,jpeg_in_a103 ,jpeg_in_a104 ,jpeg_in_a105 ,jpeg_in_a106 ,
	jpeg_in_a107 ,jpeg_in_a108 ,jpeg_in_a109 ,jpeg_in_a110 ,jpeg_in_a111 ,jpeg_in_a112 ,
	jpeg_in_a113 ,jpeg_in_a114 ,jpeg_in_a115 ,jpeg_in_a116 ,jpeg_in_a117 ,jpeg_in_a118 ,
	jpeg_in_a119 ,jpeg_in_a120 ,jpeg_in_a121 ,jpeg_in_a122 ,jpeg_in_a123 ,jpeg_in_a124 ,
	jpeg_in_a125 ,jpeg_in_a126 ,jpeg_in_a127 ,jpeg_len_in ,jpeg_out_a00 ,jpeg_out_a01 ,
	jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,jpeg_out_a06 ,jpeg_out_a07 ,
	jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,jpeg_out_a12 ,jpeg_out_a13 ,
	jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,jpeg_out_a18 ,jpeg_out_a19 ,
	jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,jpeg_out_a24 ,jpeg_out_a25 ,
	jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,jpeg_out_a30 ,jpeg_out_a31 ,
	jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,jpeg_out_a36 ,jpeg_out_a37 ,
	jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,jpeg_out_a42 ,jpeg_out_a43 ,
	jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,jpeg_out_a48 ,jpeg_out_a49 ,
	jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,jpeg_out_a54 ,jpeg_out_a55 ,
	jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,jpeg_out_a60 ,jpeg_out_a61 ,
	jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,jpeg_out_a66 ,jpeg_out_a67 ,
	jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,jpeg_out_a72 ,jpeg_out_a73 ,
	jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,jpeg_out_a78 ,jpeg_out_a79 ,
	jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,jpeg_out_a84 ,jpeg_out_a85 ,
	jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,jpeg_out_a90 ,jpeg_out_a91 ,
	jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,jpeg_out_a96 ,jpeg_out_a97 ,
	jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,jpeg_out_a102 ,
	jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,jpeg_out_a107 ,
	jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,jpeg_out_a112 ,
	jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,jpeg_out_a117 ,
	jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,jpeg_out_a122 ,
	jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,jpeg_out_a127 ,
	jpeg_len_out ,valid );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a64 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a65 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a66 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a67 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a68 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a69 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a70 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a71 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a72 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a73 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a74 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a75 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a76 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a77 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a78 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a79 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a80 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a81 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a82 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a83 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a84 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a85 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a86 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a87 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a88 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a89 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a90 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a91 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a92 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a93 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a94 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a95 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a96 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a97 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a98 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a99 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a100 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a101 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a102 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a103 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a104 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a105 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a106 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a107 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a108 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a109 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a110 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a111 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a112 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a113 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a114 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a115 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a116 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a117 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a118 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a119 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a120 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a121 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a122 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a123 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a124 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a125 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a126 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a127 ;	// line#=../rle.h:56
input	[11:0]	jpeg_len_in ;	// line#=../rle.h:57
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
wire		ST1_01d ;
wire		ST1_02d ;
wire		ST1_03d ;
wire		ST1_04d ;
wire		ST1_05d ;
wire		ST1_06d ;
wire		ST1_07d ;
wire		ST1_08d ;
wire		ST1_09d ;
wire		ST1_10d ;
wire		ST1_11d ;
wire		ST1_12d ;
wire		JF_01 ;
wire		lop8u_11ot ;
wire		JF_03 ;
wire		FL01_01_Leos_all ;
wire		JF_06 ;
wire		JF_07 ;
wire		JF_08 ;

jpeg_fsm INST_fsm ( .clk(clk) ,.rst(rst) ,.ST1_12d(ST1_12d) ,.ST1_11d(ST1_11d) ,
	.ST1_10d(ST1_10d) ,.ST1_09d(ST1_09d) ,.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,
	.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,
	.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,.JF_01(JF_01) ,.lop8u_11ot(lop8u_11ot) ,
	.JF_03(JF_03) ,.FL01_01_Leos_all(FL01_01_Leos_all) ,.JF_06(JF_06) ,.JF_07(JF_07) ,
	.JF_08(JF_08) );
jpeg_dat INST_dat ( .clk(clk) ,.rst(rst) ,.jpeg_in_a00(jpeg_in_a00) ,.jpeg_in_a01(jpeg_in_a01) ,
	.jpeg_in_a02(jpeg_in_a02) ,.jpeg_in_a03(jpeg_in_a03) ,.jpeg_in_a04(jpeg_in_a04) ,
	.jpeg_in_a05(jpeg_in_a05) ,.jpeg_in_a06(jpeg_in_a06) ,.jpeg_in_a07(jpeg_in_a07) ,
	.jpeg_in_a08(jpeg_in_a08) ,.jpeg_in_a09(jpeg_in_a09) ,.jpeg_in_a10(jpeg_in_a10) ,
	.jpeg_in_a11(jpeg_in_a11) ,.jpeg_in_a12(jpeg_in_a12) ,.jpeg_in_a13(jpeg_in_a13) ,
	.jpeg_in_a14(jpeg_in_a14) ,.jpeg_in_a15(jpeg_in_a15) ,.jpeg_in_a16(jpeg_in_a16) ,
	.jpeg_in_a17(jpeg_in_a17) ,.jpeg_in_a18(jpeg_in_a18) ,.jpeg_in_a19(jpeg_in_a19) ,
	.jpeg_in_a20(jpeg_in_a20) ,.jpeg_in_a21(jpeg_in_a21) ,.jpeg_in_a22(jpeg_in_a22) ,
	.jpeg_in_a23(jpeg_in_a23) ,.jpeg_in_a24(jpeg_in_a24) ,.jpeg_in_a25(jpeg_in_a25) ,
	.jpeg_in_a26(jpeg_in_a26) ,.jpeg_in_a27(jpeg_in_a27) ,.jpeg_in_a28(jpeg_in_a28) ,
	.jpeg_in_a29(jpeg_in_a29) ,.jpeg_in_a30(jpeg_in_a30) ,.jpeg_in_a31(jpeg_in_a31) ,
	.jpeg_in_a32(jpeg_in_a32) ,.jpeg_in_a33(jpeg_in_a33) ,.jpeg_in_a34(jpeg_in_a34) ,
	.jpeg_in_a35(jpeg_in_a35) ,.jpeg_in_a36(jpeg_in_a36) ,.jpeg_in_a37(jpeg_in_a37) ,
	.jpeg_in_a38(jpeg_in_a38) ,.jpeg_in_a39(jpeg_in_a39) ,.jpeg_in_a40(jpeg_in_a40) ,
	.jpeg_in_a41(jpeg_in_a41) ,.jpeg_in_a42(jpeg_in_a42) ,.jpeg_in_a43(jpeg_in_a43) ,
	.jpeg_in_a44(jpeg_in_a44) ,.jpeg_in_a45(jpeg_in_a45) ,.jpeg_in_a46(jpeg_in_a46) ,
	.jpeg_in_a47(jpeg_in_a47) ,.jpeg_in_a48(jpeg_in_a48) ,.jpeg_in_a49(jpeg_in_a49) ,
	.jpeg_in_a50(jpeg_in_a50) ,.jpeg_in_a51(jpeg_in_a51) ,.jpeg_in_a52(jpeg_in_a52) ,
	.jpeg_in_a53(jpeg_in_a53) ,.jpeg_in_a54(jpeg_in_a54) ,.jpeg_in_a55(jpeg_in_a55) ,
	.jpeg_in_a56(jpeg_in_a56) ,.jpeg_in_a57(jpeg_in_a57) ,.jpeg_in_a58(jpeg_in_a58) ,
	.jpeg_in_a59(jpeg_in_a59) ,.jpeg_in_a60(jpeg_in_a60) ,.jpeg_in_a61(jpeg_in_a61) ,
	.jpeg_in_a62(jpeg_in_a62) ,.jpeg_in_a63(jpeg_in_a63) ,.jpeg_out_a00(jpeg_out_a00) ,
	.jpeg_out_a01(jpeg_out_a01) ,.jpeg_out_a02(jpeg_out_a02) ,.jpeg_out_a03(jpeg_out_a03) ,
	.jpeg_out_a04(jpeg_out_a04) ,.jpeg_out_a05(jpeg_out_a05) ,.jpeg_out_a06(jpeg_out_a06) ,
	.jpeg_out_a07(jpeg_out_a07) ,.jpeg_out_a08(jpeg_out_a08) ,.jpeg_out_a09(jpeg_out_a09) ,
	.jpeg_out_a10(jpeg_out_a10) ,.jpeg_out_a11(jpeg_out_a11) ,.jpeg_out_a12(jpeg_out_a12) ,
	.jpeg_out_a13(jpeg_out_a13) ,.jpeg_out_a14(jpeg_out_a14) ,.jpeg_out_a15(jpeg_out_a15) ,
	.jpeg_out_a16(jpeg_out_a16) ,.jpeg_out_a17(jpeg_out_a17) ,.jpeg_out_a18(jpeg_out_a18) ,
	.jpeg_out_a19(jpeg_out_a19) ,.jpeg_out_a20(jpeg_out_a20) ,.jpeg_out_a21(jpeg_out_a21) ,
	.jpeg_out_a22(jpeg_out_a22) ,.jpeg_out_a23(jpeg_out_a23) ,.jpeg_out_a24(jpeg_out_a24) ,
	.jpeg_out_a25(jpeg_out_a25) ,.jpeg_out_a26(jpeg_out_a26) ,.jpeg_out_a27(jpeg_out_a27) ,
	.jpeg_out_a28(jpeg_out_a28) ,.jpeg_out_a29(jpeg_out_a29) ,.jpeg_out_a30(jpeg_out_a30) ,
	.jpeg_out_a31(jpeg_out_a31) ,.jpeg_out_a32(jpeg_out_a32) ,.jpeg_out_a33(jpeg_out_a33) ,
	.jpeg_out_a34(jpeg_out_a34) ,.jpeg_out_a35(jpeg_out_a35) ,.jpeg_out_a36(jpeg_out_a36) ,
	.jpeg_out_a37(jpeg_out_a37) ,.jpeg_out_a38(jpeg_out_a38) ,.jpeg_out_a39(jpeg_out_a39) ,
	.jpeg_out_a40(jpeg_out_a40) ,.jpeg_out_a41(jpeg_out_a41) ,.jpeg_out_a42(jpeg_out_a42) ,
	.jpeg_out_a43(jpeg_out_a43) ,.jpeg_out_a44(jpeg_out_a44) ,.jpeg_out_a45(jpeg_out_a45) ,
	.jpeg_out_a46(jpeg_out_a46) ,.jpeg_out_a47(jpeg_out_a47) ,.jpeg_out_a48(jpeg_out_a48) ,
	.jpeg_out_a49(jpeg_out_a49) ,.jpeg_out_a50(jpeg_out_a50) ,.jpeg_out_a51(jpeg_out_a51) ,
	.jpeg_out_a52(jpeg_out_a52) ,.jpeg_out_a53(jpeg_out_a53) ,.jpeg_out_a54(jpeg_out_a54) ,
	.jpeg_out_a55(jpeg_out_a55) ,.jpeg_out_a56(jpeg_out_a56) ,.jpeg_out_a57(jpeg_out_a57) ,
	.jpeg_out_a58(jpeg_out_a58) ,.jpeg_out_a59(jpeg_out_a59) ,.jpeg_out_a60(jpeg_out_a60) ,
	.jpeg_out_a61(jpeg_out_a61) ,.jpeg_out_a62(jpeg_out_a62) ,.jpeg_out_a63(jpeg_out_a63) ,
	.jpeg_out_a64(jpeg_out_a64) ,.jpeg_out_a65(jpeg_out_a65) ,.jpeg_out_a66(jpeg_out_a66) ,
	.jpeg_out_a67(jpeg_out_a67) ,.jpeg_out_a68(jpeg_out_a68) ,.jpeg_out_a69(jpeg_out_a69) ,
	.jpeg_out_a70(jpeg_out_a70) ,.jpeg_out_a71(jpeg_out_a71) ,.jpeg_out_a72(jpeg_out_a72) ,
	.jpeg_out_a73(jpeg_out_a73) ,.jpeg_out_a74(jpeg_out_a74) ,.jpeg_out_a75(jpeg_out_a75) ,
	.jpeg_out_a76(jpeg_out_a76) ,.jpeg_out_a77(jpeg_out_a77) ,.jpeg_out_a78(jpeg_out_a78) ,
	.jpeg_out_a79(jpeg_out_a79) ,.jpeg_out_a80(jpeg_out_a80) ,.jpeg_out_a81(jpeg_out_a81) ,
	.jpeg_out_a82(jpeg_out_a82) ,.jpeg_out_a83(jpeg_out_a83) ,.jpeg_out_a84(jpeg_out_a84) ,
	.jpeg_out_a85(jpeg_out_a85) ,.jpeg_out_a86(jpeg_out_a86) ,.jpeg_out_a87(jpeg_out_a87) ,
	.jpeg_out_a88(jpeg_out_a88) ,.jpeg_out_a89(jpeg_out_a89) ,.jpeg_out_a90(jpeg_out_a90) ,
	.jpeg_out_a91(jpeg_out_a91) ,.jpeg_out_a92(jpeg_out_a92) ,.jpeg_out_a93(jpeg_out_a93) ,
	.jpeg_out_a94(jpeg_out_a94) ,.jpeg_out_a95(jpeg_out_a95) ,.jpeg_out_a96(jpeg_out_a96) ,
	.jpeg_out_a97(jpeg_out_a97) ,.jpeg_out_a98(jpeg_out_a98) ,.jpeg_out_a99(jpeg_out_a99) ,
	.jpeg_out_a100(jpeg_out_a100) ,.jpeg_out_a101(jpeg_out_a101) ,.jpeg_out_a102(jpeg_out_a102) ,
	.jpeg_out_a103(jpeg_out_a103) ,.jpeg_out_a104(jpeg_out_a104) ,.jpeg_out_a105(jpeg_out_a105) ,
	.jpeg_out_a106(jpeg_out_a106) ,.jpeg_out_a107(jpeg_out_a107) ,.jpeg_out_a108(jpeg_out_a108) ,
	.jpeg_out_a109(jpeg_out_a109) ,.jpeg_out_a110(jpeg_out_a110) ,.jpeg_out_a111(jpeg_out_a111) ,
	.jpeg_out_a112(jpeg_out_a112) ,.jpeg_out_a113(jpeg_out_a113) ,.jpeg_out_a114(jpeg_out_a114) ,
	.jpeg_out_a115(jpeg_out_a115) ,.jpeg_out_a116(jpeg_out_a116) ,.jpeg_out_a117(jpeg_out_a117) ,
	.jpeg_out_a118(jpeg_out_a118) ,.jpeg_out_a119(jpeg_out_a119) ,.jpeg_out_a120(jpeg_out_a120) ,
	.jpeg_out_a121(jpeg_out_a121) ,.jpeg_out_a122(jpeg_out_a122) ,.jpeg_out_a123(jpeg_out_a123) ,
	.jpeg_out_a124(jpeg_out_a124) ,.jpeg_out_a125(jpeg_out_a125) ,.jpeg_out_a126(jpeg_out_a126) ,
	.jpeg_out_a127(jpeg_out_a127) ,.jpeg_len_out(jpeg_len_out) ,.valid(valid) ,
	.ST1_12d(ST1_12d) ,.ST1_11d(ST1_11d) ,.ST1_10d(ST1_10d) ,.ST1_09d(ST1_09d) ,
	.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,
	.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,
	.JF_01(JF_01) ,.lop8u_11ot_port(lop8u_11ot) ,.JF_03_port(JF_03) ,.FL01_01_Leos_all(FL01_01_Leos_all) ,
	.JF_06(JF_06) ,.JF_07(JF_07) ,.JF_08(JF_08) );

endmodule

module jpeg_fsm ( clk ,rst ,ST1_12d ,ST1_11d ,ST1_10d ,ST1_09d ,ST1_08d ,ST1_07d ,
	ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,ST1_02d ,ST1_01d ,JF_01 ,lop8u_11ot ,
	JF_03 ,FL01_01_Leos_all ,JF_06 ,JF_07 ,JF_08 );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
output		ST1_12d ;
output		ST1_11d ;
output		ST1_10d ;
output		ST1_09d ;
output		ST1_08d ;
output		ST1_07d ;
output		ST1_06d ;
output		ST1_05d ;
output		ST1_04d ;
output		ST1_03d ;
output		ST1_02d ;
output		ST1_01d ;
input		JF_01 ;
input		lop8u_11ot ;
input		JF_03 ;
input		FL01_01_Leos_all ;
input		JF_06 ;
input		JF_07 ;
input		JF_08 ;
reg	[3:0]	B01_streg ;

parameter	ST1_01 = 4'h0 ;
parameter	ST1_02 = 4'h1 ;
parameter	ST1_03 = 4'h2 ;
parameter	ST1_04 = 4'h3 ;
parameter	ST1_05 = 4'h4 ;
parameter	ST1_06 = 4'h5 ;
parameter	ST1_07 = 4'h6 ;
parameter	ST1_08 = 4'h7 ;
parameter	ST1_09 = 4'h8 ;
parameter	ST1_10 = 4'h9 ;
parameter	ST1_11 = 4'ha ;
parameter	ST1_12 = 4'hb ;

assign	ST1_01d = ( ( B01_streg == ST1_01 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_02d = ( ( B01_streg == ST1_02 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_03d = ( ( B01_streg == ST1_03 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_04d = ( ( B01_streg == ST1_04 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_05d = ( ( B01_streg == ST1_05 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_06d = ( ( B01_streg == ST1_06 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_07d = ( ( B01_streg == ST1_07 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_08d = ( ( B01_streg == ST1_08 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_09d = ( ( B01_streg == ST1_09 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_10d = ( ( B01_streg == ST1_10 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_11d = ( ( B01_streg == ST1_11 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_12d = ( ( B01_streg == ST1_12 ) ? 1'h1 : 1'h0 ) ;
always @ ( posedge clk )
	if ( !rst )
		B01_streg <= ST1_01 ;
	else
		case ( B01_streg )
		ST1_01 :
			B01_streg <= ST1_02 ;
		ST1_02 :
			if ( ( JF_01 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_03 ;
		ST1_03 :
			if ( ( lop8u_11ot != 1'h0 ) )
				B01_streg <= ST1_03 ;
			else
				B01_streg <= ST1_04 ;
		ST1_04 :
			if ( ( JF_03 != 1'h0 ) )
				B01_streg <= ST1_04 ;
			else
				B01_streg <= ST1_05 ;
		ST1_05 :
			if ( ( FL01_01_Leos_all != 1'h0 ) )
				B01_streg <= ST1_06 ;
			else
				B01_streg <= ST1_05 ;
		ST1_06 :
			if ( ( JF_06 != 1'h0 ) )
				B01_streg <= ST1_07 ;
			else
				B01_streg <= ST1_08 ;
		ST1_07 :
			B01_streg <= ST1_08 ;
		ST1_08 :
			if ( ( JF_07 != 1'h0 ) )
				B01_streg <= ST1_09 ;
			else
				B01_streg <= ST1_10 ;
		ST1_09 :
			B01_streg <= ST1_10 ;
		ST1_10 :
			B01_streg <= ST1_11 ;
		ST1_11 :
			if ( ( JF_08 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_12 ;
		ST1_12 :
			B01_streg <= ST1_10 ;
		default :
			B01_streg <= ST1_01 ;
		endcase

endmodule

module jpeg_dat ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,
	jpeg_in_a04 ,jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,
	jpeg_in_a10 ,jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,
	jpeg_in_a16 ,jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,
	jpeg_in_a22 ,jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,
	jpeg_in_a28 ,jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,
	jpeg_in_a34 ,jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,
	jpeg_in_a40 ,jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,
	jpeg_in_a46 ,jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,
	jpeg_in_a52 ,jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,
	jpeg_in_a58 ,jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,
	jpeg_out_a00 ,jpeg_out_a01 ,jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,
	jpeg_out_a06 ,jpeg_out_a07 ,jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,
	jpeg_out_a12 ,jpeg_out_a13 ,jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,
	jpeg_out_a18 ,jpeg_out_a19 ,jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,
	jpeg_out_a24 ,jpeg_out_a25 ,jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,
	jpeg_out_a30 ,jpeg_out_a31 ,jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,
	jpeg_out_a36 ,jpeg_out_a37 ,jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,
	jpeg_out_a42 ,jpeg_out_a43 ,jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,
	jpeg_out_a48 ,jpeg_out_a49 ,jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,
	jpeg_out_a54 ,jpeg_out_a55 ,jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,
	jpeg_out_a60 ,jpeg_out_a61 ,jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,
	jpeg_out_a66 ,jpeg_out_a67 ,jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,
	jpeg_out_a72 ,jpeg_out_a73 ,jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,
	jpeg_out_a78 ,jpeg_out_a79 ,jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,
	jpeg_out_a84 ,jpeg_out_a85 ,jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,
	jpeg_out_a90 ,jpeg_out_a91 ,jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,
	jpeg_out_a96 ,jpeg_out_a97 ,jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,
	jpeg_out_a102 ,jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,
	jpeg_out_a107 ,jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,
	jpeg_out_a112 ,jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,
	jpeg_out_a117 ,jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,
	jpeg_out_a122 ,jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,
	jpeg_out_a127 ,jpeg_len_out ,valid ,ST1_12d ,ST1_11d ,ST1_10d ,ST1_09d ,
	ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,ST1_02d ,ST1_01d ,
	JF_01 ,lop8u_11ot_port ,JF_03_port ,FL01_01_Leos_all ,JF_06 ,JF_07 ,JF_08 );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
input		ST1_12d ;
input		ST1_11d ;
input		ST1_10d ;
input		ST1_09d ;
input		ST1_08d ;
input		ST1_07d ;
input		ST1_06d ;
input		ST1_05d ;
input		ST1_04d ;
input		ST1_03d ;
input		ST1_02d ;
input		ST1_01d ;
output		JF_01 ;
output		lop8u_11ot_port ;
output		JF_03_port ;
output		FL01_01_Leos_all ;
output		JF_06 ;
output		JF_07 ;
output		JF_08 ;
wire		M_139 ;
wire		M_138 ;
wire		M_137 ;
wire		M_136 ;
wire		M_135 ;
wire		M_134 ;
wire		M_132 ;
wire		M_131 ;
wire		M_129 ;
wire		M_128 ;
wire		M_127 ;
wire		M_126 ;
wire		M_125 ;
wire		M_124 ;
wire		M_123 ;
wire		M_122 ;
wire		M_120 ;
wire		M_119 ;
wire		M_118 ;
wire		M_117 ;
wire		M_116 ;
wire		M_115 ;
wire		M_113 ;
wire		M_112 ;
wire		M_108 ;
wire		M_107 ;
wire		M_105 ;
wire		M_104 ;
wire		M_103 ;
wire		M_102 ;
wire		U_264 ;
wire		U_263 ;
wire		U_258 ;
wire		U_246 ;
wire		U_242 ;
wire		U_237 ;
wire		U_236 ;
wire		U_231 ;
wire		U_230 ;
wire		U_228 ;
wire		U_225 ;
wire		U_224 ;
wire		U_221 ;
wire		U_217 ;
wire		U_216 ;
wire		U_215 ;
wire		U_212 ;
wire		U_209 ;
wire		U_208 ;
wire		U_207 ;
wire		U_206 ;
wire		U_205 ;
wire		U_204 ;
wire		U_200 ;
wire		U_198 ;
wire		C_11 ;
wire		U_195 ;
wire		U_192 ;
wire		U_190 ;
wire		U_188 ;
wire		U_187 ;
wire		U_186 ;
wire		U_185 ;
wire		U_183 ;
wire		U_182 ;
wire		U_181 ;
wire		U_180 ;
wire		U_176 ;
wire		U_173 ;
wire		C_07 ;
wire		U_170 ;
wire		U_169 ;
wire		U_168 ;
wire		U_166 ;
wire		U_165 ;
wire		U_164 ;
wire		U_163 ;
wire		U_162 ;
wire		C_05 ;
wire		U_161 ;
wire		U_96 ;
wire		U_95 ;
wire		U_94 ;
wire		U_93 ;
wire		U_92 ;
wire		U_91 ;
wire		U_90 ;
wire		U_89 ;
wire		U_88 ;
wire		U_87 ;
wire		U_84 ;
wire		U_83 ;
wire		U_82 ;
wire		U_81 ;
wire		U_80 ;
wire		C_02 ;
wire		U_79 ;
wire		U_14 ;
wire		U_13 ;
wire		U_12 ;
wire		U_11 ;
wire		U_10 ;
wire		U_09 ;
wire		U_08 ;
wire		U_07 ;
wire		U_06 ;
wire		U_05 ;
wire		rl_we02 ;	// line#=../rle.cpp:23
wire		rl_we01 ;	// line#=../rle.cpp:23
wire	[127:0]	rl_d03 ;	// line#=../rle.cpp:23
wire	[127:0]	rl_d02 ;	// line#=../rle.cpp:23
wire	[127:0]	rl_d01 ;	// line#=../rle.cpp:23
wire	[6:0]	rl_ad03 ;	// line#=../rle.cpp:23
wire	[6:0]	rl_ad02 ;	// line#=../rle.cpp:23
wire	[6:0]	rl_ad01 ;	// line#=../rle.cpp:23
wire	[5:0]	incr8u_61i1 ;
wire	[5:0]	incr8u_61ot ;
wire	[5:0]	incr8u_71i1 ;
wire	[6:0]	incr8u_71ot ;
wire	[31:0]	decr32s2i1 ;
wire	[31:0]	decr32s2ot ;
wire	[31:0]	decr32s1i1 ;
wire	[31:0]	decr32s1ot ;
wire	[6:0]	decr8u_71i1 ;
wire	[6:0]	decr8u_71ot ;
wire	[31:0]	incr32s3i1 ;
wire	[31:0]	incr32s3ot ;
wire	[31:0]	incr32s2i1 ;
wire	[31:0]	incr32s2ot ;
wire	[31:0]	incr32s1i1 ;
wire	[31:0]	incr32s1ot ;
wire	[7:0]	incr8u2i1 ;
wire	[7:0]	incr8u2ot ;
wire	[7:0]	incr8u1i1 ;
wire	[7:0]	incr8u1ot ;
wire	[3:0]	incr4s1i1 ;
wire	[3:0]	incr4s1ot ;
wire	[5:0]	lop8u_11i2 ;
wire	[5:0]	lop8u_11i1 ;
wire		lop8u_11ot ;
wire	[8:0]	sub12s_91i2 ;
wire	[8:0]	sub12s_91i1 ;
wire	[8:0]	sub12s_91ot ;
wire	[7:0]	sub8u1i1 ;
wire	[7:0]	sub8u1ot ;
wire		FL01_05_ndat ;
wire		FL01_04_ndat ;
wire		FL01_04_rdy ;
wire		FL01_02_Lndat ;
wire		FL01_02_Lrdy ;
wire		FL01_02_ndat ;
wire		FL01_02_rdy ;
wire		FL01_01_ndat ;
wire		FL01_06_eos ;
wire		FL01_05_eos ;
wire		FL01_04_eos ;
wire		FL01_03_eos ;
wire		FL01_02_eos ;
wire		FL01_01_eos ;
wire		FL01_02_Leos_all ;
wire		FL01_02_Leos ;
wire		FL01_01_Leos_all ;
wire		FJ_07_08 ;
wire		FJ_05_11 ;
wire		FL01_06_01a ;
wire		FL01_05_01a ;
wire		FL01_04_01a ;
wire		FL01_03_01a ;
wire		FL01_02_01a ;
wire		FL01_01_01a ;
wire		FL01_03_break ;
wire		FL01_02_break ;
wire		FL01_01_break ;
wire		JF_08 ;
wire		JF_07 ;
wire		CT_32 ;
wire		CT_31 ;
wire		CT_26 ;
wire		JF_03 ;
wire		CT_12 ;
wire		JF_01 ;
wire		zz_WE1 ;
wire	[8:0]	zz_RD2 ;
wire	[8:0]	zz_RD1 ;
wire	[8:0]	zz_RD3 ;
wire		RG_previous_dc_en ;
wire		RG_quantized_block_en ;
wire		RG_quantized_block_1_en ;
wire		RG_quantized_block_2_en ;
wire		RG_quantized_block_3_en ;
wire		RG_quantized_block_4_en ;
wire		RG_quantized_block_5_en ;
wire		RG_quantized_block_6_en ;
wire		RG_quantized_block_7_en ;
wire		RG_quantized_block_8_en ;
wire		RG_quantized_block_9_en ;
wire		RG_quantized_block_10_en ;
wire		RG_quantized_block_11_en ;
wire		RG_quantized_block_12_en ;
wire		RG_quantized_block_13_en ;
wire		RG_quantized_block_14_en ;
wire		RG_quantized_block_15_en ;
wire		RG_quantized_block_16_en ;
wire		RG_quantized_block_17_en ;
wire		RG_quantized_block_18_en ;
wire		RG_quantized_block_19_en ;
wire		RG_quantized_block_20_en ;
wire		RG_quantized_block_21_en ;
wire		RG_quantized_block_22_en ;
wire		RG_quantized_block_23_en ;
wire		RG_quantized_block_24_en ;
wire		RG_quantized_block_25_en ;
wire		RG_quantized_block_26_en ;
wire		RG_quantized_block_27_en ;
wire		RG_quantized_block_28_en ;
wire		RG_quantized_block_29_en ;
wire		RG_quantized_block_30_en ;
wire		RG_quantized_block_31_en ;
wire		RG_quantized_block_32_en ;
wire		RG_quantized_block_33_en ;
wire		RG_quantized_block_34_en ;
wire		RG_quantized_block_35_en ;
wire		RG_quantized_block_36_en ;
wire		RG_quantized_block_37_en ;
wire		RG_quantized_block_38_en ;
wire		RG_quantized_block_39_en ;
wire		RG_quantized_block_40_en ;
wire		RG_quantized_block_41_en ;
wire		RG_quantized_block_42_en ;
wire		RG_quantized_block_43_en ;
wire		RG_quantized_block_44_en ;
wire		RG_quantized_block_45_en ;
wire		RG_quantized_block_46_en ;
wire		RG_quantized_block_47_en ;
wire		RG_quantized_block_48_en ;
wire		RG_quantized_block_49_en ;
wire		RG_quantized_block_50_en ;
wire		RG_quantized_block_51_en ;
wire		RG_quantized_block_52_en ;
wire		RG_quantized_block_53_en ;
wire		RG_quantized_block_54_en ;
wire		RG_quantized_block_55_en ;
wire		RG_quantized_block_56_en ;
wire		RG_quantized_block_57_en ;
wire		RG_quantized_block_58_en ;
wire		RG_quantized_block_59_en ;
wire		RG_zz_02_en ;
wire		FF_j_en ;
wire		RG_quantized_block_60_en ;
wire		RG_i_05_en ;
wire		RG_i_04_en ;
wire		RG_i_03_en ;
wire		RG_i_02_en ;
wire		RG_k_02_en ;
wire		jpeg_out_a00_r_en ;
wire		jpeg_out_a01_r_en ;
wire		jpeg_out_a02_r_en ;
wire		jpeg_out_a03_r_en ;
wire		jpeg_out_a04_r_en ;
wire		jpeg_out_a05_r_en ;
wire		jpeg_out_a06_r_en ;
wire		jpeg_out_a07_r_en ;
wire		jpeg_out_a08_r_en ;
wire		jpeg_out_a09_r_en ;
wire		jpeg_out_a10_r_en ;
wire		jpeg_out_a11_r_en ;
wire		jpeg_out_a12_r_en ;
wire		jpeg_out_a13_r_en ;
wire		jpeg_out_a14_r_en ;
wire		jpeg_out_a15_r_en ;
wire		jpeg_out_a16_r_en ;
wire		jpeg_out_a17_r_en ;
wire		jpeg_out_a18_r_en ;
wire		jpeg_out_a19_r_en ;
wire		jpeg_out_a20_r_en ;
wire		jpeg_out_a21_r_en ;
wire		jpeg_out_a22_r_en ;
wire		jpeg_out_a23_r_en ;
wire		jpeg_out_a24_r_en ;
wire		jpeg_out_a25_r_en ;
wire		jpeg_out_a26_r_en ;
wire		jpeg_out_a27_r_en ;
wire		jpeg_out_a28_r_en ;
wire		jpeg_out_a29_r_en ;
wire		jpeg_out_a30_r_en ;
wire		jpeg_out_a31_r_en ;
wire		jpeg_out_a32_r_en ;
wire		jpeg_out_a33_r_en ;
wire		jpeg_out_a34_r_en ;
wire		jpeg_out_a35_r_en ;
wire		jpeg_out_a36_r_en ;
wire		jpeg_out_a37_r_en ;
wire		jpeg_out_a38_r_en ;
wire		jpeg_out_a39_r_en ;
wire		jpeg_out_a40_r_en ;
wire		jpeg_out_a41_r_en ;
wire		jpeg_out_a42_r_en ;
wire		jpeg_out_a43_r_en ;
wire		jpeg_out_a44_r_en ;
wire		jpeg_out_a45_r_en ;
wire		jpeg_out_a46_r_en ;
wire		jpeg_out_a47_r_en ;
wire		jpeg_out_a48_r_en ;
wire		jpeg_out_a49_r_en ;
wire		jpeg_out_a50_r_en ;
wire		jpeg_out_a51_r_en ;
wire		jpeg_out_a52_r_en ;
wire		jpeg_out_a53_r_en ;
wire		jpeg_out_a54_r_en ;
wire		jpeg_out_a55_r_en ;
wire		jpeg_out_a56_r_en ;
wire		jpeg_out_a57_r_en ;
wire		jpeg_out_a58_r_en ;
wire		jpeg_out_a59_r_en ;
wire		jpeg_out_a60_r_en ;
wire		jpeg_out_a61_r_en ;
wire		jpeg_out_a62_r_en ;
wire		jpeg_out_a63_r_en ;
wire		jpeg_out_a64_r_en ;
wire		jpeg_out_a65_r_en ;
wire		jpeg_out_a66_r_en ;
wire		jpeg_out_a67_r_en ;
wire		jpeg_out_a68_r_en ;
wire		jpeg_out_a69_r_en ;
wire		jpeg_out_a70_r_en ;
wire		jpeg_out_a71_r_en ;
wire		jpeg_out_a72_r_en ;
wire		jpeg_out_a73_r_en ;
wire		jpeg_out_a74_r_en ;
wire		jpeg_out_a75_r_en ;
wire		jpeg_out_a76_r_en ;
wire		jpeg_out_a77_r_en ;
wire		jpeg_out_a78_r_en ;
wire		jpeg_out_a79_r_en ;
wire		jpeg_out_a80_r_en ;
wire		jpeg_out_a81_r_en ;
wire		jpeg_out_a82_r_en ;
wire		jpeg_out_a83_r_en ;
wire		jpeg_out_a84_r_en ;
wire		jpeg_out_a85_r_en ;
wire		jpeg_out_a86_r_en ;
wire		jpeg_out_a87_r_en ;
wire		jpeg_out_a88_r_en ;
wire		jpeg_out_a89_r_en ;
wire		jpeg_out_a90_r_en ;
wire		jpeg_out_a91_r_en ;
wire		jpeg_out_a92_r_en ;
wire		jpeg_out_a93_r_en ;
wire		jpeg_out_a94_r_en ;
wire		jpeg_out_a95_r_en ;
wire		jpeg_out_a96_r_en ;
wire		jpeg_out_a97_r_en ;
wire		jpeg_out_a98_r_en ;
wire		jpeg_out_a99_r_en ;
wire		jpeg_out_a100_r_en ;
wire		jpeg_out_a101_r_en ;
wire		jpeg_out_a102_r_en ;
wire		jpeg_out_a103_r_en ;
wire		jpeg_out_a104_r_en ;
wire		jpeg_out_a105_r_en ;
wire		jpeg_out_a106_r_en ;
wire		jpeg_out_a107_r_en ;
wire		jpeg_out_a108_r_en ;
wire		jpeg_out_a109_r_en ;
wire		jpeg_out_a110_r_en ;
wire		jpeg_out_a111_r_en ;
wire		jpeg_out_a112_r_en ;
wire		jpeg_out_a113_r_en ;
wire		jpeg_out_a114_r_en ;
wire		jpeg_out_a115_r_en ;
wire		jpeg_out_a116_r_en ;
wire		jpeg_out_a117_r_en ;
wire		jpeg_out_a118_r_en ;
wire		jpeg_out_a119_r_en ;
wire		jpeg_out_a120_r_en ;
wire		jpeg_out_a121_r_en ;
wire		jpeg_out_a122_r_en ;
wire		jpeg_out_a123_r_en ;
wire		jpeg_out_a124_r_en ;
wire		jpeg_out_a125_r_en ;
wire		jpeg_out_a126_r_en ;
wire		jpeg_out_a127_r_en ;
wire		jpeg_len_out_r_en ;
wire		M_01 ;
wire		rl_rg00_en ;
wire		rl_rg01_en ;
wire		rl_rg02_en ;
wire		rl_rg03_en ;
wire		rl_rg04_en ;
wire		rl_rg05_en ;
wire		rl_rg06_en ;
wire		rl_rg07_en ;
wire		rl_rg08_en ;
wire		rl_rg09_en ;
wire		rl_rg10_en ;
wire		rl_rg11_en ;
wire		rl_rg12_en ;
wire		rl_rg13_en ;
wire		rl_rg14_en ;
wire		rl_rg15_en ;
wire		rl_rg16_en ;
wire		rl_rg17_en ;
wire		rl_rg18_en ;
wire		rl_rg19_en ;
wire		rl_rg20_en ;
wire		rl_rg21_en ;
wire		rl_rg22_en ;
wire		rl_rg23_en ;
wire		rl_rg24_en ;
wire		rl_rg25_en ;
wire		rl_rg26_en ;
wire		rl_rg27_en ;
wire		rl_rg28_en ;
wire		rl_rg29_en ;
wire		rl_rg30_en ;
wire		rl_rg31_en ;
wire		rl_rg32_en ;
wire		rl_rg33_en ;
wire		rl_rg34_en ;
wire		rl_rg35_en ;
wire		rl_rg36_en ;
wire		rl_rg37_en ;
wire		rl_rg38_en ;
wire		rl_rg39_en ;
wire		rl_rg40_en ;
wire		rl_rg41_en ;
wire		rl_rg42_en ;
wire		rl_rg43_en ;
wire		rl_rg44_en ;
wire		rl_rg45_en ;
wire		rl_rg46_en ;
wire		rl_rg47_en ;
wire		rl_rg48_en ;
wire		rl_rg49_en ;
wire		rl_rg50_en ;
wire		rl_rg51_en ;
wire		rl_rg52_en ;
wire		rl_rg53_en ;
wire		rl_rg54_en ;
wire		rl_rg55_en ;
wire		rl_rg56_en ;
wire		rl_rg57_en ;
wire		rl_rg58_en ;
wire		rl_rg59_en ;
wire		rl_rg60_en ;
wire		rl_rg61_en ;
wire		rl_rg62_en ;
wire		rl_rg63_en ;
wire		rl_rg64_en ;
wire		rl_rg65_en ;
wire		rl_rg66_en ;
wire		rl_rg67_en ;
wire		rl_rg68_en ;
wire		rl_rg69_en ;
wire		rl_rg70_en ;
wire		rl_rg71_en ;
wire		rl_rg72_en ;
wire		rl_rg73_en ;
wire		rl_rg74_en ;
wire		rl_rg75_en ;
wire		rl_rg76_en ;
wire		rl_rg77_en ;
wire		rl_rg78_en ;
wire		rl_rg79_en ;
wire		rl_rg80_en ;
wire		rl_rg81_en ;
wire		rl_rg82_en ;
wire		rl_rg83_en ;
wire		rl_rg84_en ;
wire		rl_rg85_en ;
wire		rl_rg86_en ;
wire		rl_rg87_en ;
wire		rl_rg88_en ;
wire		rl_rg89_en ;
wire		rl_rg90_en ;
wire		rl_rg91_en ;
wire		rl_rg92_en ;
wire		rl_rg93_en ;
wire		rl_rg94_en ;
wire		rl_rg95_en ;
wire		rl_rg96_en ;
wire		rl_rg97_en ;
wire		rl_rg98_en ;
wire		rl_rg99_en ;
wire		rl_rg100_en ;
wire		rl_rg101_en ;
wire		rl_rg102_en ;
wire		rl_rg103_en ;
wire		rl_rg104_en ;
wire		rl_rg105_en ;
wire		rl_rg106_en ;
wire		rl_rg107_en ;
wire		rl_rg108_en ;
wire		rl_rg109_en ;
wire		rl_rg110_en ;
wire		rl_rg111_en ;
wire		rl_rg112_en ;
wire		rl_rg113_en ;
wire		rl_rg114_en ;
wire		rl_rg115_en ;
wire		rl_rg116_en ;
wire		rl_rg117_en ;
wire		rl_rg118_en ;
wire		rl_rg119_en ;
wire		rl_rg120_en ;
wire		rl_rg121_en ;
wire		rl_rg122_en ;
wire		rl_rg123_en ;
wire		rl_rg124_en ;
wire		rl_rg125_en ;
wire		rl_rg126_en ;
wire		rl_rg127_en ;
wire		RG_i_06_en ;
wire		RG_i_en ;
wire		RG_j_k_en ;
wire		RG_k_quantized_block_04_en ;
wire		RG_k_quantized_block_03_en ;
wire		RG_previous_dc_quantized_block_en ;
wire		RG_len_05_en ;
wire		FF_d_02_en ;
wire		RG_76_05_en ;
wire		RG_k_05_en ;
wire		flag_r1_en ;
wire		flag_r2_en ;
wire		flag_r3_en ;
wire		FL01_01_streg_en ;
wire		FL01_02_streg_en ;
wire		FL01_03_streg_en ;
wire		FL01_04_streg_en ;
wire		FL01_05_streg_en ;
wire		FL01_06_streg_en ;
wire		valid_r_en ;
reg	[8:0]	rl_rg127 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg126 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg125 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg124 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg123 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg122 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg121 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg120 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg119 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg118 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg117 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg116 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg115 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg114 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg113 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg112 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg111 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg110 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg109 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg108 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg107 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg106 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg105 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg104 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg103 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg102 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg101 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg100 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg99 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg98 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg97 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg96 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg95 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg94 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg93 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg92 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg91 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg90 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg89 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg88 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg87 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg86 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg85 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg84 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg83 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg82 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg81 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg80 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg79 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg78 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg77 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg76 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg75 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg74 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg73 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg72 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg71 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg70 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg69 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg68 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg67 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg66 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg65 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg64 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg63 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg62 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg61 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg60 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg59 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg58 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg57 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg56 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg55 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg54 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg53 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg52 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg51 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg50 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg49 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg48 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg47 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg46 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg45 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg44 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg43 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg42 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg41 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg40 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg39 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg38 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg37 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg36 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg35 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg34 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg33 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg32 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg31 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg30 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg29 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg28 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg27 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg26 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg25 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg24 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg23 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg22 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg21 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg20 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg19 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg18 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg17 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg16 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg15 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg14 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg13 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg12 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg11 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg10 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg09 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg08 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg07 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg06 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg05 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg04 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg03 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg02 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg01 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg00 ;	// line#=../rle.cpp:23
reg	FL01_06_streg ;
reg	FL01_05_streg ;
reg	FL01_04_streg ;
reg	FL01_03_streg ;
reg	[1:0]	FL01_02_streg ;
reg	[1:0]	FL01_01_streg ;
reg	flag_r3 ;
reg	flag_r2 ;
reg	flag_r1 ;
reg	[8:0]	RG_previous_dc ;	// line#=../rle.h:66
reg	[3:0]	RG_j ;	// line#=../rle.cpp:27
reg	[31:0]	RG_i_06 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_i ;	// line#=../rle.cpp:25,105
reg	[31:0]	RG_j_k ;	// line#=../rle.cpp:25,105
reg	[8:0]	RG_quantized_block ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_1 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_2 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_3 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_4 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_5 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_6 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_7 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_8 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_9 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_10 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_11 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_12 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_13 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_14 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_15 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_16 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_17 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_18 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_19 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_20 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_21 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_22 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_23 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_24 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_25 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_26 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_27 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_28 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_29 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_30 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_31 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_32 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_33 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_34 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_35 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_36 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_37 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_38 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_39 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_40 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_41 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_42 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_43 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_44 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_45 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_46 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_47 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_48 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_49 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_50 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_51 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_52 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_53 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_54 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_55 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_56 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_57 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_58 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_59 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_k_quantized_block_04 ;	// line#=../rle.cpp:22,25
reg	[8:0]	RG_k_quantized_block_03 ;	// line#=../rle.cpp:22,25
reg	[8:0]	RG_zz_02 ;	// line#=../rle.h:65
reg	[8:0]	RG_previous_dc_quantized_block ;	// line#=../rle.cpp:22 ../rle.h:66
reg	[7:0]	RG_len_05 ;	// line#=../rle.cpp:24
reg	[5:0]	RG_k ;	// line#=../rle.cpp:105
reg	FF_d_02 ;	// line#=../rle.cpp:105
reg	FF_j ;	// line#=../rle.cpp:27
reg	[8:0]	RG_quantized_block_60 ;	// line#=../rle.cpp:22
reg	[31:0]	RG_i_05 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_i_04 ;	// line#=../rle.cpp:25
reg	RG_76_05 ;
reg	[31:0]	RG_i_03 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_i_02 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_k_02 ;	// line#=../rle.cpp:25
reg	[6:0]	RG_k_05 ;	// line#=../rle.cpp:105
reg	[8:0]	jpeg_out_a00_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a01_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a02_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a03_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a04_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a05_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a06_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a07_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a08_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a09_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a10_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a11_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a12_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a13_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a14_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a15_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a16_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a17_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a18_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a19_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a20_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a21_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a22_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a23_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a24_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a25_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a26_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a27_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a28_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a29_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a30_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a31_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a32_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a33_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a34_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a35_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a36_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a37_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a38_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a39_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a40_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a41_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a42_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a43_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a44_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a45_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a46_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a47_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a48_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a49_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a50_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a51_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a52_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a53_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a54_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a55_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a56_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a57_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a58_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a59_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a60_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a61_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a62_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a63_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a64_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a65_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a66_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a67_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a68_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a69_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a70_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a71_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a72_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a73_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a74_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a75_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a76_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a77_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a78_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a79_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a80_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a81_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a82_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a83_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a84_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a85_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a86_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a87_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a88_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a89_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a90_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a91_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a92_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a93_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a94_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a95_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a96_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a97_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a98_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a99_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a100_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a101_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a102_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a103_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a104_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a105_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a106_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a107_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a108_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a109_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a110_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a111_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a112_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a113_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a114_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a115_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a116_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a117_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a118_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a119_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a120_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a121_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a122_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a123_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a124_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a125_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a126_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a127_r ;	// line#=../rle.h:60
reg	[11:0]	jpeg_len_out_r ;	// line#=../rle.h:61
reg	valid_r ;	// line#=../rle.h:62
reg	[8:0]	rl_rd00 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg00_t ;
reg	rl_rg00_t_c1 ;
reg	rl_rg00_t_c2 ;
reg	rl_rg00_t_c3 ;
reg	rl_rg00_t_c4 ;
reg	[8:0]	rl_rg01_t ;
reg	rl_rg01_t_c1 ;
reg	rl_rg01_t_c2 ;
reg	rl_rg01_t_c3 ;
reg	[8:0]	rl_rg02_t ;
reg	rl_rg02_t_c1 ;
reg	rl_rg02_t_c2 ;
reg	rl_rg02_t_c3 ;
reg	[8:0]	rl_rg03_t ;
reg	rl_rg03_t_c1 ;
reg	rl_rg03_t_c2 ;
reg	rl_rg03_t_c3 ;
reg	[8:0]	rl_rg04_t ;
reg	rl_rg04_t_c1 ;
reg	rl_rg04_t_c2 ;
reg	rl_rg04_t_c3 ;
reg	[8:0]	rl_rg05_t ;
reg	rl_rg05_t_c1 ;
reg	rl_rg05_t_c2 ;
reg	rl_rg05_t_c3 ;
reg	[8:0]	rl_rg06_t ;
reg	rl_rg06_t_c1 ;
reg	rl_rg06_t_c2 ;
reg	rl_rg06_t_c3 ;
reg	[8:0]	rl_rg07_t ;
reg	rl_rg07_t_c1 ;
reg	rl_rg07_t_c2 ;
reg	rl_rg07_t_c3 ;
reg	[8:0]	rl_rg08_t ;
reg	rl_rg08_t_c1 ;
reg	rl_rg08_t_c2 ;
reg	rl_rg08_t_c3 ;
reg	[8:0]	rl_rg09_t ;
reg	rl_rg09_t_c1 ;
reg	rl_rg09_t_c2 ;
reg	rl_rg09_t_c3 ;
reg	[8:0]	rl_rg10_t ;
reg	rl_rg10_t_c1 ;
reg	rl_rg10_t_c2 ;
reg	rl_rg10_t_c3 ;
reg	[8:0]	rl_rg11_t ;
reg	rl_rg11_t_c1 ;
reg	rl_rg11_t_c2 ;
reg	rl_rg11_t_c3 ;
reg	[8:0]	rl_rg12_t ;
reg	rl_rg12_t_c1 ;
reg	rl_rg12_t_c2 ;
reg	rl_rg12_t_c3 ;
reg	[8:0]	rl_rg13_t ;
reg	rl_rg13_t_c1 ;
reg	rl_rg13_t_c2 ;
reg	rl_rg13_t_c3 ;
reg	[8:0]	rl_rg14_t ;
reg	rl_rg14_t_c1 ;
reg	rl_rg14_t_c2 ;
reg	rl_rg14_t_c3 ;
reg	[8:0]	rl_rg15_t ;
reg	rl_rg15_t_c1 ;
reg	rl_rg15_t_c2 ;
reg	rl_rg15_t_c3 ;
reg	[8:0]	rl_rg16_t ;
reg	rl_rg16_t_c1 ;
reg	rl_rg16_t_c2 ;
reg	rl_rg16_t_c3 ;
reg	[8:0]	rl_rg17_t ;
reg	rl_rg17_t_c1 ;
reg	rl_rg17_t_c2 ;
reg	rl_rg17_t_c3 ;
reg	[8:0]	rl_rg18_t ;
reg	rl_rg18_t_c1 ;
reg	rl_rg18_t_c2 ;
reg	rl_rg18_t_c3 ;
reg	[8:0]	rl_rg19_t ;
reg	rl_rg19_t_c1 ;
reg	rl_rg19_t_c2 ;
reg	rl_rg19_t_c3 ;
reg	[8:0]	rl_rg20_t ;
reg	rl_rg20_t_c1 ;
reg	rl_rg20_t_c2 ;
reg	rl_rg20_t_c3 ;
reg	[8:0]	rl_rg21_t ;
reg	rl_rg21_t_c1 ;
reg	rl_rg21_t_c2 ;
reg	rl_rg21_t_c3 ;
reg	[8:0]	rl_rg22_t ;
reg	rl_rg22_t_c1 ;
reg	rl_rg22_t_c2 ;
reg	rl_rg22_t_c3 ;
reg	[8:0]	rl_rg23_t ;
reg	rl_rg23_t_c1 ;
reg	rl_rg23_t_c2 ;
reg	rl_rg23_t_c3 ;
reg	[8:0]	rl_rg24_t ;
reg	rl_rg24_t_c1 ;
reg	rl_rg24_t_c2 ;
reg	rl_rg24_t_c3 ;
reg	[8:0]	rl_rg25_t ;
reg	rl_rg25_t_c1 ;
reg	rl_rg25_t_c2 ;
reg	rl_rg25_t_c3 ;
reg	[8:0]	rl_rg26_t ;
reg	rl_rg26_t_c1 ;
reg	rl_rg26_t_c2 ;
reg	rl_rg26_t_c3 ;
reg	[8:0]	rl_rg27_t ;
reg	rl_rg27_t_c1 ;
reg	rl_rg27_t_c2 ;
reg	rl_rg27_t_c3 ;
reg	[8:0]	rl_rg28_t ;
reg	rl_rg28_t_c1 ;
reg	rl_rg28_t_c2 ;
reg	rl_rg28_t_c3 ;
reg	[8:0]	rl_rg29_t ;
reg	rl_rg29_t_c1 ;
reg	rl_rg29_t_c2 ;
reg	rl_rg29_t_c3 ;
reg	[8:0]	rl_rg30_t ;
reg	rl_rg30_t_c1 ;
reg	rl_rg30_t_c2 ;
reg	rl_rg30_t_c3 ;
reg	[8:0]	rl_rg31_t ;
reg	rl_rg31_t_c1 ;
reg	rl_rg31_t_c2 ;
reg	rl_rg31_t_c3 ;
reg	[8:0]	rl_rg32_t ;
reg	rl_rg32_t_c1 ;
reg	rl_rg32_t_c2 ;
reg	rl_rg32_t_c3 ;
reg	[8:0]	rl_rg33_t ;
reg	rl_rg33_t_c1 ;
reg	rl_rg33_t_c2 ;
reg	rl_rg33_t_c3 ;
reg	[8:0]	rl_rg34_t ;
reg	rl_rg34_t_c1 ;
reg	rl_rg34_t_c2 ;
reg	rl_rg34_t_c3 ;
reg	[8:0]	rl_rg35_t ;
reg	rl_rg35_t_c1 ;
reg	rl_rg35_t_c2 ;
reg	rl_rg35_t_c3 ;
reg	[8:0]	rl_rg36_t ;
reg	rl_rg36_t_c1 ;
reg	rl_rg36_t_c2 ;
reg	rl_rg36_t_c3 ;
reg	[8:0]	rl_rg37_t ;
reg	rl_rg37_t_c1 ;
reg	rl_rg37_t_c2 ;
reg	rl_rg37_t_c3 ;
reg	[8:0]	rl_rg38_t ;
reg	rl_rg38_t_c1 ;
reg	rl_rg38_t_c2 ;
reg	rl_rg38_t_c3 ;
reg	[8:0]	rl_rg39_t ;
reg	rl_rg39_t_c1 ;
reg	rl_rg39_t_c2 ;
reg	rl_rg39_t_c3 ;
reg	[8:0]	rl_rg40_t ;
reg	rl_rg40_t_c1 ;
reg	rl_rg40_t_c2 ;
reg	rl_rg40_t_c3 ;
reg	[8:0]	rl_rg41_t ;
reg	rl_rg41_t_c1 ;
reg	rl_rg41_t_c2 ;
reg	rl_rg41_t_c3 ;
reg	[8:0]	rl_rg42_t ;
reg	rl_rg42_t_c1 ;
reg	rl_rg42_t_c2 ;
reg	rl_rg42_t_c3 ;
reg	[8:0]	rl_rg43_t ;
reg	rl_rg43_t_c1 ;
reg	rl_rg43_t_c2 ;
reg	rl_rg43_t_c3 ;
reg	[8:0]	rl_rg44_t ;
reg	rl_rg44_t_c1 ;
reg	rl_rg44_t_c2 ;
reg	rl_rg44_t_c3 ;
reg	[8:0]	rl_rg45_t ;
reg	rl_rg45_t_c1 ;
reg	rl_rg45_t_c2 ;
reg	rl_rg45_t_c3 ;
reg	[8:0]	rl_rg46_t ;
reg	rl_rg46_t_c1 ;
reg	rl_rg46_t_c2 ;
reg	rl_rg46_t_c3 ;
reg	[8:0]	rl_rg47_t ;
reg	rl_rg47_t_c1 ;
reg	rl_rg47_t_c2 ;
reg	rl_rg47_t_c3 ;
reg	[8:0]	rl_rg48_t ;
reg	rl_rg48_t_c1 ;
reg	rl_rg48_t_c2 ;
reg	rl_rg48_t_c3 ;
reg	[8:0]	rl_rg49_t ;
reg	rl_rg49_t_c1 ;
reg	rl_rg49_t_c2 ;
reg	rl_rg49_t_c3 ;
reg	[8:0]	rl_rg50_t ;
reg	rl_rg50_t_c1 ;
reg	rl_rg50_t_c2 ;
reg	rl_rg50_t_c3 ;
reg	[8:0]	rl_rg51_t ;
reg	rl_rg51_t_c1 ;
reg	rl_rg51_t_c2 ;
reg	rl_rg51_t_c3 ;
reg	[8:0]	rl_rg52_t ;
reg	rl_rg52_t_c1 ;
reg	rl_rg52_t_c2 ;
reg	rl_rg52_t_c3 ;
reg	[8:0]	rl_rg53_t ;
reg	rl_rg53_t_c1 ;
reg	rl_rg53_t_c2 ;
reg	rl_rg53_t_c3 ;
reg	[8:0]	rl_rg54_t ;
reg	rl_rg54_t_c1 ;
reg	rl_rg54_t_c2 ;
reg	rl_rg54_t_c3 ;
reg	[8:0]	rl_rg55_t ;
reg	rl_rg55_t_c1 ;
reg	rl_rg55_t_c2 ;
reg	rl_rg55_t_c3 ;
reg	[8:0]	rl_rg56_t ;
reg	rl_rg56_t_c1 ;
reg	rl_rg56_t_c2 ;
reg	rl_rg56_t_c3 ;
reg	[8:0]	rl_rg57_t ;
reg	rl_rg57_t_c1 ;
reg	rl_rg57_t_c2 ;
reg	rl_rg57_t_c3 ;
reg	[8:0]	rl_rg58_t ;
reg	rl_rg58_t_c1 ;
reg	rl_rg58_t_c2 ;
reg	rl_rg58_t_c3 ;
reg	[8:0]	rl_rg59_t ;
reg	rl_rg59_t_c1 ;
reg	rl_rg59_t_c2 ;
reg	rl_rg59_t_c3 ;
reg	[8:0]	rl_rg60_t ;
reg	rl_rg60_t_c1 ;
reg	rl_rg60_t_c2 ;
reg	rl_rg60_t_c3 ;
reg	[8:0]	rl_rg61_t ;
reg	rl_rg61_t_c1 ;
reg	rl_rg61_t_c2 ;
reg	rl_rg61_t_c3 ;
reg	[8:0]	rl_rg62_t ;
reg	rl_rg62_t_c1 ;
reg	rl_rg62_t_c2 ;
reg	rl_rg62_t_c3 ;
reg	[8:0]	rl_rg63_t ;
reg	rl_rg63_t_c1 ;
reg	rl_rg63_t_c2 ;
reg	rl_rg63_t_c3 ;
reg	[8:0]	rl_rg64_t ;
reg	rl_rg64_t_c1 ;
reg	rl_rg64_t_c2 ;
reg	rl_rg64_t_c3 ;
reg	[8:0]	rl_rg65_t ;
reg	rl_rg65_t_c1 ;
reg	rl_rg65_t_c2 ;
reg	rl_rg65_t_c3 ;
reg	[8:0]	rl_rg66_t ;
reg	rl_rg66_t_c1 ;
reg	rl_rg66_t_c2 ;
reg	rl_rg66_t_c3 ;
reg	[8:0]	rl_rg67_t ;
reg	rl_rg67_t_c1 ;
reg	rl_rg67_t_c2 ;
reg	rl_rg67_t_c3 ;
reg	[8:0]	rl_rg68_t ;
reg	rl_rg68_t_c1 ;
reg	rl_rg68_t_c2 ;
reg	rl_rg68_t_c3 ;
reg	[8:0]	rl_rg69_t ;
reg	rl_rg69_t_c1 ;
reg	rl_rg69_t_c2 ;
reg	rl_rg69_t_c3 ;
reg	[8:0]	rl_rg70_t ;
reg	rl_rg70_t_c1 ;
reg	rl_rg70_t_c2 ;
reg	rl_rg70_t_c3 ;
reg	[8:0]	rl_rg71_t ;
reg	rl_rg71_t_c1 ;
reg	rl_rg71_t_c2 ;
reg	rl_rg71_t_c3 ;
reg	[8:0]	rl_rg72_t ;
reg	rl_rg72_t_c1 ;
reg	rl_rg72_t_c2 ;
reg	rl_rg72_t_c3 ;
reg	[8:0]	rl_rg73_t ;
reg	rl_rg73_t_c1 ;
reg	rl_rg73_t_c2 ;
reg	rl_rg73_t_c3 ;
reg	[8:0]	rl_rg74_t ;
reg	rl_rg74_t_c1 ;
reg	rl_rg74_t_c2 ;
reg	rl_rg74_t_c3 ;
reg	[8:0]	rl_rg75_t ;
reg	rl_rg75_t_c1 ;
reg	rl_rg75_t_c2 ;
reg	rl_rg75_t_c3 ;
reg	[8:0]	rl_rg76_t ;
reg	rl_rg76_t_c1 ;
reg	rl_rg76_t_c2 ;
reg	rl_rg76_t_c3 ;
reg	[8:0]	rl_rg77_t ;
reg	rl_rg77_t_c1 ;
reg	rl_rg77_t_c2 ;
reg	rl_rg77_t_c3 ;
reg	[8:0]	rl_rg78_t ;
reg	rl_rg78_t_c1 ;
reg	rl_rg78_t_c2 ;
reg	rl_rg78_t_c3 ;
reg	[8:0]	rl_rg79_t ;
reg	rl_rg79_t_c1 ;
reg	rl_rg79_t_c2 ;
reg	rl_rg79_t_c3 ;
reg	[8:0]	rl_rg80_t ;
reg	rl_rg80_t_c1 ;
reg	rl_rg80_t_c2 ;
reg	rl_rg80_t_c3 ;
reg	[8:0]	rl_rg81_t ;
reg	rl_rg81_t_c1 ;
reg	rl_rg81_t_c2 ;
reg	rl_rg81_t_c3 ;
reg	[8:0]	rl_rg82_t ;
reg	rl_rg82_t_c1 ;
reg	rl_rg82_t_c2 ;
reg	rl_rg82_t_c3 ;
reg	[8:0]	rl_rg83_t ;
reg	rl_rg83_t_c1 ;
reg	rl_rg83_t_c2 ;
reg	rl_rg83_t_c3 ;
reg	[8:0]	rl_rg84_t ;
reg	rl_rg84_t_c1 ;
reg	rl_rg84_t_c2 ;
reg	rl_rg84_t_c3 ;
reg	[8:0]	rl_rg85_t ;
reg	rl_rg85_t_c1 ;
reg	rl_rg85_t_c2 ;
reg	rl_rg85_t_c3 ;
reg	[8:0]	rl_rg86_t ;
reg	rl_rg86_t_c1 ;
reg	rl_rg86_t_c2 ;
reg	rl_rg86_t_c3 ;
reg	[8:0]	rl_rg87_t ;
reg	rl_rg87_t_c1 ;
reg	rl_rg87_t_c2 ;
reg	rl_rg87_t_c3 ;
reg	[8:0]	rl_rg88_t ;
reg	rl_rg88_t_c1 ;
reg	rl_rg88_t_c2 ;
reg	rl_rg88_t_c3 ;
reg	[8:0]	rl_rg89_t ;
reg	rl_rg89_t_c1 ;
reg	rl_rg89_t_c2 ;
reg	rl_rg89_t_c3 ;
reg	[8:0]	rl_rg90_t ;
reg	rl_rg90_t_c1 ;
reg	rl_rg90_t_c2 ;
reg	rl_rg90_t_c3 ;
reg	[8:0]	rl_rg91_t ;
reg	rl_rg91_t_c1 ;
reg	rl_rg91_t_c2 ;
reg	rl_rg91_t_c3 ;
reg	[8:0]	rl_rg92_t ;
reg	rl_rg92_t_c1 ;
reg	rl_rg92_t_c2 ;
reg	rl_rg92_t_c3 ;
reg	[8:0]	rl_rg93_t ;
reg	rl_rg93_t_c1 ;
reg	rl_rg93_t_c2 ;
reg	rl_rg93_t_c3 ;
reg	[8:0]	rl_rg94_t ;
reg	rl_rg94_t_c1 ;
reg	rl_rg94_t_c2 ;
reg	rl_rg94_t_c3 ;
reg	[8:0]	rl_rg95_t ;
reg	rl_rg95_t_c1 ;
reg	rl_rg95_t_c2 ;
reg	rl_rg95_t_c3 ;
reg	[8:0]	rl_rg96_t ;
reg	rl_rg96_t_c1 ;
reg	rl_rg96_t_c2 ;
reg	rl_rg96_t_c3 ;
reg	[8:0]	rl_rg97_t ;
reg	rl_rg97_t_c1 ;
reg	rl_rg97_t_c2 ;
reg	rl_rg97_t_c3 ;
reg	[8:0]	rl_rg98_t ;
reg	rl_rg98_t_c1 ;
reg	rl_rg98_t_c2 ;
reg	rl_rg98_t_c3 ;
reg	[8:0]	rl_rg99_t ;
reg	rl_rg99_t_c1 ;
reg	rl_rg99_t_c2 ;
reg	rl_rg99_t_c3 ;
reg	[8:0]	rl_rg100_t ;
reg	rl_rg100_t_c1 ;
reg	rl_rg100_t_c2 ;
reg	rl_rg100_t_c3 ;
reg	[8:0]	rl_rg101_t ;
reg	rl_rg101_t_c1 ;
reg	rl_rg101_t_c2 ;
reg	rl_rg101_t_c3 ;
reg	[8:0]	rl_rg102_t ;
reg	rl_rg102_t_c1 ;
reg	rl_rg102_t_c2 ;
reg	rl_rg102_t_c3 ;
reg	[8:0]	rl_rg103_t ;
reg	rl_rg103_t_c1 ;
reg	rl_rg103_t_c2 ;
reg	rl_rg103_t_c3 ;
reg	[8:0]	rl_rg104_t ;
reg	rl_rg104_t_c1 ;
reg	rl_rg104_t_c2 ;
reg	rl_rg104_t_c3 ;
reg	[8:0]	rl_rg105_t ;
reg	rl_rg105_t_c1 ;
reg	rl_rg105_t_c2 ;
reg	rl_rg105_t_c3 ;
reg	[8:0]	rl_rg106_t ;
reg	rl_rg106_t_c1 ;
reg	rl_rg106_t_c2 ;
reg	rl_rg106_t_c3 ;
reg	[8:0]	rl_rg107_t ;
reg	rl_rg107_t_c1 ;
reg	rl_rg107_t_c2 ;
reg	rl_rg107_t_c3 ;
reg	[8:0]	rl_rg108_t ;
reg	rl_rg108_t_c1 ;
reg	rl_rg108_t_c2 ;
reg	rl_rg108_t_c3 ;
reg	[8:0]	rl_rg109_t ;
reg	rl_rg109_t_c1 ;
reg	rl_rg109_t_c2 ;
reg	rl_rg109_t_c3 ;
reg	[8:0]	rl_rg110_t ;
reg	rl_rg110_t_c1 ;
reg	rl_rg110_t_c2 ;
reg	rl_rg110_t_c3 ;
reg	[8:0]	rl_rg111_t ;
reg	rl_rg111_t_c1 ;
reg	rl_rg111_t_c2 ;
reg	rl_rg111_t_c3 ;
reg	[8:0]	rl_rg112_t ;
reg	rl_rg112_t_c1 ;
reg	rl_rg112_t_c2 ;
reg	rl_rg112_t_c3 ;
reg	[8:0]	rl_rg113_t ;
reg	rl_rg113_t_c1 ;
reg	rl_rg113_t_c2 ;
reg	rl_rg113_t_c3 ;
reg	[8:0]	rl_rg114_t ;
reg	rl_rg114_t_c1 ;
reg	rl_rg114_t_c2 ;
reg	rl_rg114_t_c3 ;
reg	[8:0]	rl_rg115_t ;
reg	rl_rg115_t_c1 ;
reg	rl_rg115_t_c2 ;
reg	rl_rg115_t_c3 ;
reg	[8:0]	rl_rg116_t ;
reg	rl_rg116_t_c1 ;
reg	rl_rg116_t_c2 ;
reg	rl_rg116_t_c3 ;
reg	[8:0]	rl_rg117_t ;
reg	rl_rg117_t_c1 ;
reg	rl_rg117_t_c2 ;
reg	rl_rg117_t_c3 ;
reg	[8:0]	rl_rg118_t ;
reg	rl_rg118_t_c1 ;
reg	rl_rg118_t_c2 ;
reg	rl_rg118_t_c3 ;
reg	[8:0]	rl_rg119_t ;
reg	rl_rg119_t_c1 ;
reg	rl_rg119_t_c2 ;
reg	rl_rg119_t_c3 ;
reg	[8:0]	rl_rg120_t ;
reg	rl_rg120_t_c1 ;
reg	rl_rg120_t_c2 ;
reg	rl_rg120_t_c3 ;
reg	[8:0]	rl_rg121_t ;
reg	rl_rg121_t_c1 ;
reg	rl_rg121_t_c2 ;
reg	rl_rg121_t_c3 ;
reg	[8:0]	rl_rg122_t ;
reg	rl_rg122_t_c1 ;
reg	rl_rg122_t_c2 ;
reg	rl_rg122_t_c3 ;
reg	[8:0]	rl_rg123_t ;
reg	rl_rg123_t_c1 ;
reg	rl_rg123_t_c2 ;
reg	rl_rg123_t_c3 ;
reg	[8:0]	rl_rg124_t ;
reg	rl_rg124_t_c1 ;
reg	rl_rg124_t_c2 ;
reg	rl_rg124_t_c3 ;
reg	[8:0]	rl_rg125_t ;
reg	rl_rg125_t_c1 ;
reg	rl_rg125_t_c2 ;
reg	rl_rg125_t_c3 ;
reg	[8:0]	rl_rg126_t ;
reg	rl_rg126_t_c1 ;
reg	rl_rg126_t_c2 ;
reg	rl_rg126_t_c3 ;
reg	[8:0]	rl_rg127_t ;
reg	rl_rg127_t_c1 ;
reg	rl_rg127_t_c2 ;
reg	rl_rg127_t_c3 ;
reg	M_01_t1 ;
reg	JF_06 ;
reg	CT_35 ;
reg	[3:0]	RG_j_t ;
reg	[31:0]	RG_i_06_t ;
reg	RG_i_06_t_c1 ;
reg	RG_i_06_t_c2 ;
reg	[2:0]	TR_01 ;
reg	[31:0]	RG_i_t ;
reg	RG_i_t_c1 ;
reg	RG_i_t_c2 ;
reg	[31:0]	RG_j_k_t ;
reg	RG_j_k_t_c1 ;
reg	RG_j_k_t_c2 ;
reg	RG_j_k_t_c3 ;
reg	[8:0]	RG_k_quantized_block_04_t ;
reg	[8:0]	RG_k_quantized_block_03_t ;
reg	[8:0]	RG_previous_dc_quantized_block_t ;
reg	[7:0]	RG_len_05_t ;
reg	RG_len_05_t_c1 ;
reg	[5:0]	RG_k_t ;
reg	FF_d_02_t ;
reg	FF_d_02_t_c1 ;
reg	FF_d_02_t_c2 ;
reg	RG_76_05_t ;
reg	[6:0]	RG_k_05_t ;
reg	flag_r1_t ;
reg	flag_r1_t_c1 ;
reg	flag_r2_t ;
reg	flag_r2_t_c1 ;
reg	flag_r3_t ;
reg	flag_r3_t_c1 ;
reg	[1:0]	FL01_01_streg_t ;
reg	FL01_01_streg_t_c1 ;
reg	FL01_01_streg_t_c2 ;
reg	[1:0]	FL01_02_streg_t ;
reg	FL01_02_streg_t_c1 ;
reg	FL01_02_streg_t_c2 ;
reg	[1:0]	FL01_02_streg_t1 ;
reg	FL01_02_streg_t1_c1 ;
reg	FL01_02_streg_t1_c2 ;
reg	FL01_02_streg_t1_c3 ;
reg	FL01_03_streg_t ;
reg	FL01_03_streg_t_c1 ;
reg	FL01_03_streg_t_c2 ;
reg	FL01_04_streg_t ;
reg	FL01_04_streg_t_c1 ;
reg	FL01_04_streg_t_c2 ;
reg	FL01_05_streg_t ;
reg	FL01_05_streg_t_c1 ;
reg	FL01_05_streg_t_c2 ;
reg	FL01_06_streg_t ;
reg	FL01_06_streg_t_c1 ;
reg	FL01_06_streg_t_c2 ;
reg	valid_r_t ;
reg	[2:0]	sub8u1i2 ;
reg	sub8u1i2_c1 ;
reg	[5:0]	zz_AD1 ;
reg	zz_AD1_c1 ;
reg	zz_AD1_c2 ;
reg	[8:0]	TR_06 ;
reg	[8:0]	TR_07 ;
reg	[8:0]	TR_08 ;
reg	[8:0]	TR_09 ;
reg	[8:0]	TR_10 ;
reg	[8:0]	TR_11 ;
reg	[8:0]	TR_12 ;
reg	[8:0]	TR_13 ;
reg	[8:0]	zz_WD1 ;
reg	[6:0]	rl_ad00 ;	// line#=../rle.cpp:23
reg	rl_ad00_c1 ;
reg	[8:0]	rl_wd02 ;	// line#=../rle.cpp:23

jpeg_incr8u_6 INST_incr8u_6_1 ( .i1(incr8u_61i1) ,.o1(incr8u_61ot) );	// line#=../rle.cpp:111
jpeg_incr8u_7 INST_incr8u_7_1 ( .i1(incr8u_71i1) ,.o1(incr8u_71ot) );	// line#=../rle.cpp:142
jpeg_decr32s INST_decr32s_1 ( .i1(decr32s1i1) ,.o1(decr32s1ot) );	// line#=../rle.cpp:124,155
jpeg_decr32s INST_decr32s_2 ( .i1(decr32s2i1) ,.o1(decr32s2ot) );	// line#=../rle.cpp:130,161
jpeg_decr8u_7 INST_decr8u_7_1 ( .i1(decr8u_71i1) ,.o1(decr8u_71ot) );	// line#=../rle.cpp:77,78
jpeg_incr32s INST_incr32s_1 ( .i1(incr32s1i1) ,.o1(incr32s1ot) );	// line#=../rle.cpp:64,114,125,145,156
jpeg_incr32s INST_incr32s_2 ( .i1(incr32s2i1) ,.o1(incr32s2ot) );	// line#=../rle.cpp:61,62,63,119,129,150
									// ,160
jpeg_incr32s INST_incr32s_3 ( .i1(incr32s3i1) ,.o1(incr32s3ot) );	// line#=../rle.cpp:74
jpeg_incr8u INST_incr8u_1 ( .i1(incr8u1i1) ,.o1(incr8u1ot) );	// line#=../rle.cpp:68,73,79,80
jpeg_incr8u INST_incr8u_2 ( .i1(incr8u2i1) ,.o1(incr8u2ot) );	// line#=../rle.cpp:69,74
jpeg_incr4s INST_incr4s_1 ( .i1(incr4s1i1) ,.o1(incr4s1ot) );	// line#=../rle.cpp:34
jpeg_lop8u_1 INST_lop8u_1_1 ( .i1(lop8u_11i1) ,.i2(lop8u_11i2) ,.o1(lop8u_11ot) );	// line#=../rle.cpp:109,110
assign	lop8u_11ot_port = lop8u_11ot ;
jpeg_sub12s_9 INST_sub12s_9_1 ( .i1(sub12s_91i1) ,.i2(sub12s_91i2) ,.o1(sub12s_91ot) );	// line#=../rle.cpp:52
jpeg_sub8u INST_sub8u_1 ( .i1(sub8u1i1) ,.i2(sub8u1i2) ,.o1(sub8u1ot) );	// line#=../rle.cpp:77,78,83,84,86
assign	jpeg_out_a00 = jpeg_out_a00_r ;	// line#=../rle.h:60
assign	jpeg_out_a01 = jpeg_out_a01_r ;	// line#=../rle.h:60
assign	jpeg_out_a02 = jpeg_out_a02_r ;	// line#=../rle.h:60
assign	jpeg_out_a03 = jpeg_out_a03_r ;	// line#=../rle.h:60
assign	jpeg_out_a04 = jpeg_out_a04_r ;	// line#=../rle.h:60
assign	jpeg_out_a05 = jpeg_out_a05_r ;	// line#=../rle.h:60
assign	jpeg_out_a06 = jpeg_out_a06_r ;	// line#=../rle.h:60
assign	jpeg_out_a07 = jpeg_out_a07_r ;	// line#=../rle.h:60
assign	jpeg_out_a08 = jpeg_out_a08_r ;	// line#=../rle.h:60
assign	jpeg_out_a09 = jpeg_out_a09_r ;	// line#=../rle.h:60
assign	jpeg_out_a10 = jpeg_out_a10_r ;	// line#=../rle.h:60
assign	jpeg_out_a11 = jpeg_out_a11_r ;	// line#=../rle.h:60
assign	jpeg_out_a12 = jpeg_out_a12_r ;	// line#=../rle.h:60
assign	jpeg_out_a13 = jpeg_out_a13_r ;	// line#=../rle.h:60
assign	jpeg_out_a14 = jpeg_out_a14_r ;	// line#=../rle.h:60
assign	jpeg_out_a15 = jpeg_out_a15_r ;	// line#=../rle.h:60
assign	jpeg_out_a16 = jpeg_out_a16_r ;	// line#=../rle.h:60
assign	jpeg_out_a17 = jpeg_out_a17_r ;	// line#=../rle.h:60
assign	jpeg_out_a18 = jpeg_out_a18_r ;	// line#=../rle.h:60
assign	jpeg_out_a19 = jpeg_out_a19_r ;	// line#=../rle.h:60
assign	jpeg_out_a20 = jpeg_out_a20_r ;	// line#=../rle.h:60
assign	jpeg_out_a21 = jpeg_out_a21_r ;	// line#=../rle.h:60
assign	jpeg_out_a22 = jpeg_out_a22_r ;	// line#=../rle.h:60
assign	jpeg_out_a23 = jpeg_out_a23_r ;	// line#=../rle.h:60
assign	jpeg_out_a24 = jpeg_out_a24_r ;	// line#=../rle.h:60
assign	jpeg_out_a25 = jpeg_out_a25_r ;	// line#=../rle.h:60
assign	jpeg_out_a26 = jpeg_out_a26_r ;	// line#=../rle.h:60
assign	jpeg_out_a27 = jpeg_out_a27_r ;	// line#=../rle.h:60
assign	jpeg_out_a28 = jpeg_out_a28_r ;	// line#=../rle.h:60
assign	jpeg_out_a29 = jpeg_out_a29_r ;	// line#=../rle.h:60
assign	jpeg_out_a30 = jpeg_out_a30_r ;	// line#=../rle.h:60
assign	jpeg_out_a31 = jpeg_out_a31_r ;	// line#=../rle.h:60
assign	jpeg_out_a32 = jpeg_out_a32_r ;	// line#=../rle.h:60
assign	jpeg_out_a33 = jpeg_out_a33_r ;	// line#=../rle.h:60
assign	jpeg_out_a34 = jpeg_out_a34_r ;	// line#=../rle.h:60
assign	jpeg_out_a35 = jpeg_out_a35_r ;	// line#=../rle.h:60
assign	jpeg_out_a36 = jpeg_out_a36_r ;	// line#=../rle.h:60
assign	jpeg_out_a37 = jpeg_out_a37_r ;	// line#=../rle.h:60
assign	jpeg_out_a38 = jpeg_out_a38_r ;	// line#=../rle.h:60
assign	jpeg_out_a39 = jpeg_out_a39_r ;	// line#=../rle.h:60
assign	jpeg_out_a40 = jpeg_out_a40_r ;	// line#=../rle.h:60
assign	jpeg_out_a41 = jpeg_out_a41_r ;	// line#=../rle.h:60
assign	jpeg_out_a42 = jpeg_out_a42_r ;	// line#=../rle.h:60
assign	jpeg_out_a43 = jpeg_out_a43_r ;	// line#=../rle.h:60
assign	jpeg_out_a44 = jpeg_out_a44_r ;	// line#=../rle.h:60
assign	jpeg_out_a45 = jpeg_out_a45_r ;	// line#=../rle.h:60
assign	jpeg_out_a46 = jpeg_out_a46_r ;	// line#=../rle.h:60
assign	jpeg_out_a47 = jpeg_out_a47_r ;	// line#=../rle.h:60
assign	jpeg_out_a48 = jpeg_out_a48_r ;	// line#=../rle.h:60
assign	jpeg_out_a49 = jpeg_out_a49_r ;	// line#=../rle.h:60
assign	jpeg_out_a50 = jpeg_out_a50_r ;	// line#=../rle.h:60
assign	jpeg_out_a51 = jpeg_out_a51_r ;	// line#=../rle.h:60
assign	jpeg_out_a52 = jpeg_out_a52_r ;	// line#=../rle.h:60
assign	jpeg_out_a53 = jpeg_out_a53_r ;	// line#=../rle.h:60
assign	jpeg_out_a54 = jpeg_out_a54_r ;	// line#=../rle.h:60
assign	jpeg_out_a55 = jpeg_out_a55_r ;	// line#=../rle.h:60
assign	jpeg_out_a56 = jpeg_out_a56_r ;	// line#=../rle.h:60
assign	jpeg_out_a57 = jpeg_out_a57_r ;	// line#=../rle.h:60
assign	jpeg_out_a58 = jpeg_out_a58_r ;	// line#=../rle.h:60
assign	jpeg_out_a59 = jpeg_out_a59_r ;	// line#=../rle.h:60
assign	jpeg_out_a60 = jpeg_out_a60_r ;	// line#=../rle.h:60
assign	jpeg_out_a61 = jpeg_out_a61_r ;	// line#=../rle.h:60
assign	jpeg_out_a62 = jpeg_out_a62_r ;	// line#=../rle.h:60
assign	jpeg_out_a63 = jpeg_out_a63_r ;	// line#=../rle.h:60
assign	jpeg_out_a64 = jpeg_out_a64_r ;	// line#=../rle.h:60
assign	jpeg_out_a65 = jpeg_out_a65_r ;	// line#=../rle.h:60
assign	jpeg_out_a66 = jpeg_out_a66_r ;	// line#=../rle.h:60
assign	jpeg_out_a67 = jpeg_out_a67_r ;	// line#=../rle.h:60
assign	jpeg_out_a68 = jpeg_out_a68_r ;	// line#=../rle.h:60
assign	jpeg_out_a69 = jpeg_out_a69_r ;	// line#=../rle.h:60
assign	jpeg_out_a70 = jpeg_out_a70_r ;	// line#=../rle.h:60
assign	jpeg_out_a71 = jpeg_out_a71_r ;	// line#=../rle.h:60
assign	jpeg_out_a72 = jpeg_out_a72_r ;	// line#=../rle.h:60
assign	jpeg_out_a73 = jpeg_out_a73_r ;	// line#=../rle.h:60
assign	jpeg_out_a74 = jpeg_out_a74_r ;	// line#=../rle.h:60
assign	jpeg_out_a75 = jpeg_out_a75_r ;	// line#=../rle.h:60
assign	jpeg_out_a76 = jpeg_out_a76_r ;	// line#=../rle.h:60
assign	jpeg_out_a77 = jpeg_out_a77_r ;	// line#=../rle.h:60
assign	jpeg_out_a78 = jpeg_out_a78_r ;	// line#=../rle.h:60
assign	jpeg_out_a79 = jpeg_out_a79_r ;	// line#=../rle.h:60
assign	jpeg_out_a80 = jpeg_out_a80_r ;	// line#=../rle.h:60
assign	jpeg_out_a81 = jpeg_out_a81_r ;	// line#=../rle.h:60
assign	jpeg_out_a82 = jpeg_out_a82_r ;	// line#=../rle.h:60
assign	jpeg_out_a83 = jpeg_out_a83_r ;	// line#=../rle.h:60
assign	jpeg_out_a84 = jpeg_out_a84_r ;	// line#=../rle.h:60
assign	jpeg_out_a85 = jpeg_out_a85_r ;	// line#=../rle.h:60
assign	jpeg_out_a86 = jpeg_out_a86_r ;	// line#=../rle.h:60
assign	jpeg_out_a87 = jpeg_out_a87_r ;	// line#=../rle.h:60
assign	jpeg_out_a88 = jpeg_out_a88_r ;	// line#=../rle.h:60
assign	jpeg_out_a89 = jpeg_out_a89_r ;	// line#=../rle.h:60
assign	jpeg_out_a90 = jpeg_out_a90_r ;	// line#=../rle.h:60
assign	jpeg_out_a91 = jpeg_out_a91_r ;	// line#=../rle.h:60
assign	jpeg_out_a92 = jpeg_out_a92_r ;	// line#=../rle.h:60
assign	jpeg_out_a93 = jpeg_out_a93_r ;	// line#=../rle.h:60
assign	jpeg_out_a94 = jpeg_out_a94_r ;	// line#=../rle.h:60
assign	jpeg_out_a95 = jpeg_out_a95_r ;	// line#=../rle.h:60
assign	jpeg_out_a96 = jpeg_out_a96_r ;	// line#=../rle.h:60
assign	jpeg_out_a97 = jpeg_out_a97_r ;	// line#=../rle.h:60
assign	jpeg_out_a98 = jpeg_out_a98_r ;	// line#=../rle.h:60
assign	jpeg_out_a99 = jpeg_out_a99_r ;	// line#=../rle.h:60
assign	jpeg_out_a100 = jpeg_out_a100_r ;	// line#=../rle.h:60
assign	jpeg_out_a101 = jpeg_out_a101_r ;	// line#=../rle.h:60
assign	jpeg_out_a102 = jpeg_out_a102_r ;	// line#=../rle.h:60
assign	jpeg_out_a103 = jpeg_out_a103_r ;	// line#=../rle.h:60
assign	jpeg_out_a104 = jpeg_out_a104_r ;	// line#=../rle.h:60
assign	jpeg_out_a105 = jpeg_out_a105_r ;	// line#=../rle.h:60
assign	jpeg_out_a106 = jpeg_out_a106_r ;	// line#=../rle.h:60
assign	jpeg_out_a107 = jpeg_out_a107_r ;	// line#=../rle.h:60
assign	jpeg_out_a108 = jpeg_out_a108_r ;	// line#=../rle.h:60
assign	jpeg_out_a109 = jpeg_out_a109_r ;	// line#=../rle.h:60
assign	jpeg_out_a110 = jpeg_out_a110_r ;	// line#=../rle.h:60
assign	jpeg_out_a111 = jpeg_out_a111_r ;	// line#=../rle.h:60
assign	jpeg_out_a112 = jpeg_out_a112_r ;	// line#=../rle.h:60
assign	jpeg_out_a113 = jpeg_out_a113_r ;	// line#=../rle.h:60
assign	jpeg_out_a114 = jpeg_out_a114_r ;	// line#=../rle.h:60
assign	jpeg_out_a115 = jpeg_out_a115_r ;	// line#=../rle.h:60
assign	jpeg_out_a116 = jpeg_out_a116_r ;	// line#=../rle.h:60
assign	jpeg_out_a117 = jpeg_out_a117_r ;	// line#=../rle.h:60
assign	jpeg_out_a118 = jpeg_out_a118_r ;	// line#=../rle.h:60
assign	jpeg_out_a119 = jpeg_out_a119_r ;	// line#=../rle.h:60
assign	jpeg_out_a120 = jpeg_out_a120_r ;	// line#=../rle.h:60
assign	jpeg_out_a121 = jpeg_out_a121_r ;	// line#=../rle.h:60
assign	jpeg_out_a122 = jpeg_out_a122_r ;	// line#=../rle.h:60
assign	jpeg_out_a123 = jpeg_out_a123_r ;	// line#=../rle.h:60
assign	jpeg_out_a124 = jpeg_out_a124_r ;	// line#=../rle.h:60
assign	jpeg_out_a125 = jpeg_out_a125_r ;	// line#=../rle.h:60
assign	jpeg_out_a126 = jpeg_out_a126_r ;	// line#=../rle.h:60
assign	jpeg_out_a127 = jpeg_out_a127_r ;	// line#=../rle.h:60
assign	jpeg_len_out = jpeg_len_out_r ;	// line#=../rle.h:61
assign	valid = valid_r ;	// line#=../rle.h:62
jpeg_decoder_7to128 INST_decoder_7to128_1 ( .DECODER_in(rl_ad01) ,.DECODER_out(rl_d01) );	// line#=../rle.cpp:23
jpeg_decoder_7to128 INST_decoder_7to128_2 ( .DECODER_in(rl_ad02) ,.DECODER_out(rl_d02) );	// line#=../rle.cpp:23
jpeg_decoder_7to128 INST_decoder_7to128_3 ( .DECODER_in(rl_ad03) ,.DECODER_out(rl_d03) );	// line#=../rle.cpp:23
always @ ( rl_rg127 or rl_rg126 or rl_rg125 or rl_rg124 or rl_rg123 or rl_rg122 or 
	rl_rg121 or rl_rg120 or rl_rg119 or rl_rg118 or rl_rg117 or rl_rg116 or 
	rl_rg115 or rl_rg114 or rl_rg113 or rl_rg112 or rl_rg111 or rl_rg110 or 
	rl_rg109 or rl_rg108 or rl_rg107 or rl_rg106 or rl_rg105 or rl_rg104 or 
	rl_rg103 or rl_rg102 or rl_rg101 or rl_rg100 or rl_rg99 or rl_rg98 or rl_rg97 or 
	rl_rg96 or rl_rg95 or rl_rg94 or rl_rg93 or rl_rg92 or rl_rg91 or rl_rg90 or 
	rl_rg89 or rl_rg88 or rl_rg87 or rl_rg86 or rl_rg85 or rl_rg84 or rl_rg83 or 
	rl_rg82 or rl_rg81 or rl_rg80 or rl_rg79 or rl_rg78 or rl_rg77 or rl_rg76 or 
	rl_rg75 or rl_rg74 or rl_rg73 or rl_rg72 or rl_rg71 or rl_rg70 or rl_rg69 or 
	rl_rg68 or rl_rg67 or rl_rg66 or rl_rg65 or rl_rg64 or rl_rg63 or rl_rg62 or 
	rl_rg61 or rl_rg60 or rl_rg59 or rl_rg58 or rl_rg57 or rl_rg56 or rl_rg55 or 
	rl_rg54 or rl_rg53 or rl_rg52 or rl_rg51 or rl_rg50 or rl_rg49 or rl_rg48 or 
	rl_rg47 or rl_rg46 or rl_rg45 or rl_rg44 or rl_rg43 or rl_rg42 or rl_rg41 or 
	rl_rg40 or rl_rg39 or rl_rg38 or rl_rg37 or rl_rg36 or rl_rg35 or rl_rg34 or 
	rl_rg33 or rl_rg32 or rl_rg31 or rl_rg30 or rl_rg29 or rl_rg28 or rl_rg27 or 
	rl_rg26 or rl_rg25 or rl_rg24 or rl_rg23 or rl_rg22 or rl_rg21 or rl_rg20 or 
	rl_rg19 or rl_rg18 or rl_rg17 or rl_rg16 or rl_rg15 or rl_rg14 or rl_rg13 or 
	rl_rg12 or rl_rg11 or rl_rg10 or rl_rg09 or rl_rg08 or rl_rg07 or rl_rg06 or 
	rl_rg05 or rl_rg04 or rl_rg03 or rl_rg02 or rl_rg01 or rl_rg00 or rl_ad00 )	// line#=../rle.cpp:23
	case ( rl_ad00 )
	7'h00 :
		rl_rd00 = rl_rg00 ;
	7'h01 :
		rl_rd00 = rl_rg01 ;
	7'h02 :
		rl_rd00 = rl_rg02 ;
	7'h03 :
		rl_rd00 = rl_rg03 ;
	7'h04 :
		rl_rd00 = rl_rg04 ;
	7'h05 :
		rl_rd00 = rl_rg05 ;
	7'h06 :
		rl_rd00 = rl_rg06 ;
	7'h07 :
		rl_rd00 = rl_rg07 ;
	7'h08 :
		rl_rd00 = rl_rg08 ;
	7'h09 :
		rl_rd00 = rl_rg09 ;
	7'h0a :
		rl_rd00 = rl_rg10 ;
	7'h0b :
		rl_rd00 = rl_rg11 ;
	7'h0c :
		rl_rd00 = rl_rg12 ;
	7'h0d :
		rl_rd00 = rl_rg13 ;
	7'h0e :
		rl_rd00 = rl_rg14 ;
	7'h0f :
		rl_rd00 = rl_rg15 ;
	7'h10 :
		rl_rd00 = rl_rg16 ;
	7'h11 :
		rl_rd00 = rl_rg17 ;
	7'h12 :
		rl_rd00 = rl_rg18 ;
	7'h13 :
		rl_rd00 = rl_rg19 ;
	7'h14 :
		rl_rd00 = rl_rg20 ;
	7'h15 :
		rl_rd00 = rl_rg21 ;
	7'h16 :
		rl_rd00 = rl_rg22 ;
	7'h17 :
		rl_rd00 = rl_rg23 ;
	7'h18 :
		rl_rd00 = rl_rg24 ;
	7'h19 :
		rl_rd00 = rl_rg25 ;
	7'h1a :
		rl_rd00 = rl_rg26 ;
	7'h1b :
		rl_rd00 = rl_rg27 ;
	7'h1c :
		rl_rd00 = rl_rg28 ;
	7'h1d :
		rl_rd00 = rl_rg29 ;
	7'h1e :
		rl_rd00 = rl_rg30 ;
	7'h1f :
		rl_rd00 = rl_rg31 ;
	7'h20 :
		rl_rd00 = rl_rg32 ;
	7'h21 :
		rl_rd00 = rl_rg33 ;
	7'h22 :
		rl_rd00 = rl_rg34 ;
	7'h23 :
		rl_rd00 = rl_rg35 ;
	7'h24 :
		rl_rd00 = rl_rg36 ;
	7'h25 :
		rl_rd00 = rl_rg37 ;
	7'h26 :
		rl_rd00 = rl_rg38 ;
	7'h27 :
		rl_rd00 = rl_rg39 ;
	7'h28 :
		rl_rd00 = rl_rg40 ;
	7'h29 :
		rl_rd00 = rl_rg41 ;
	7'h2a :
		rl_rd00 = rl_rg42 ;
	7'h2b :
		rl_rd00 = rl_rg43 ;
	7'h2c :
		rl_rd00 = rl_rg44 ;
	7'h2d :
		rl_rd00 = rl_rg45 ;
	7'h2e :
		rl_rd00 = rl_rg46 ;
	7'h2f :
		rl_rd00 = rl_rg47 ;
	7'h30 :
		rl_rd00 = rl_rg48 ;
	7'h31 :
		rl_rd00 = rl_rg49 ;
	7'h32 :
		rl_rd00 = rl_rg50 ;
	7'h33 :
		rl_rd00 = rl_rg51 ;
	7'h34 :
		rl_rd00 = rl_rg52 ;
	7'h35 :
		rl_rd00 = rl_rg53 ;
	7'h36 :
		rl_rd00 = rl_rg54 ;
	7'h37 :
		rl_rd00 = rl_rg55 ;
	7'h38 :
		rl_rd00 = rl_rg56 ;
	7'h39 :
		rl_rd00 = rl_rg57 ;
	7'h3a :
		rl_rd00 = rl_rg58 ;
	7'h3b :
		rl_rd00 = rl_rg59 ;
	7'h3c :
		rl_rd00 = rl_rg60 ;
	7'h3d :
		rl_rd00 = rl_rg61 ;
	7'h3e :
		rl_rd00 = rl_rg62 ;
	7'h3f :
		rl_rd00 = rl_rg63 ;
	7'h40 :
		rl_rd00 = rl_rg64 ;
	7'h41 :
		rl_rd00 = rl_rg65 ;
	7'h42 :
		rl_rd00 = rl_rg66 ;
	7'h43 :
		rl_rd00 = rl_rg67 ;
	7'h44 :
		rl_rd00 = rl_rg68 ;
	7'h45 :
		rl_rd00 = rl_rg69 ;
	7'h46 :
		rl_rd00 = rl_rg70 ;
	7'h47 :
		rl_rd00 = rl_rg71 ;
	7'h48 :
		rl_rd00 = rl_rg72 ;
	7'h49 :
		rl_rd00 = rl_rg73 ;
	7'h4a :
		rl_rd00 = rl_rg74 ;
	7'h4b :
		rl_rd00 = rl_rg75 ;
	7'h4c :
		rl_rd00 = rl_rg76 ;
	7'h4d :
		rl_rd00 = rl_rg77 ;
	7'h4e :
		rl_rd00 = rl_rg78 ;
	7'h4f :
		rl_rd00 = rl_rg79 ;
	7'h50 :
		rl_rd00 = rl_rg80 ;
	7'h51 :
		rl_rd00 = rl_rg81 ;
	7'h52 :
		rl_rd00 = rl_rg82 ;
	7'h53 :
		rl_rd00 = rl_rg83 ;
	7'h54 :
		rl_rd00 = rl_rg84 ;
	7'h55 :
		rl_rd00 = rl_rg85 ;
	7'h56 :
		rl_rd00 = rl_rg86 ;
	7'h57 :
		rl_rd00 = rl_rg87 ;
	7'h58 :
		rl_rd00 = rl_rg88 ;
	7'h59 :
		rl_rd00 = rl_rg89 ;
	7'h5a :
		rl_rd00 = rl_rg90 ;
	7'h5b :
		rl_rd00 = rl_rg91 ;
	7'h5c :
		rl_rd00 = rl_rg92 ;
	7'h5d :
		rl_rd00 = rl_rg93 ;
	7'h5e :
		rl_rd00 = rl_rg94 ;
	7'h5f :
		rl_rd00 = rl_rg95 ;
	7'h60 :
		rl_rd00 = rl_rg96 ;
	7'h61 :
		rl_rd00 = rl_rg97 ;
	7'h62 :
		rl_rd00 = rl_rg98 ;
	7'h63 :
		rl_rd00 = rl_rg99 ;
	7'h64 :
		rl_rd00 = rl_rg100 ;
	7'h65 :
		rl_rd00 = rl_rg101 ;
	7'h66 :
		rl_rd00 = rl_rg102 ;
	7'h67 :
		rl_rd00 = rl_rg103 ;
	7'h68 :
		rl_rd00 = rl_rg104 ;
	7'h69 :
		rl_rd00 = rl_rg105 ;
	7'h6a :
		rl_rd00 = rl_rg106 ;
	7'h6b :
		rl_rd00 = rl_rg107 ;
	7'h6c :
		rl_rd00 = rl_rg108 ;
	7'h6d :
		rl_rd00 = rl_rg109 ;
	7'h6e :
		rl_rd00 = rl_rg110 ;
	7'h6f :
		rl_rd00 = rl_rg111 ;
	7'h70 :
		rl_rd00 = rl_rg112 ;
	7'h71 :
		rl_rd00 = rl_rg113 ;
	7'h72 :
		rl_rd00 = rl_rg114 ;
	7'h73 :
		rl_rd00 = rl_rg115 ;
	7'h74 :
		rl_rd00 = rl_rg116 ;
	7'h75 :
		rl_rd00 = rl_rg117 ;
	7'h76 :
		rl_rd00 = rl_rg118 ;
	7'h77 :
		rl_rd00 = rl_rg119 ;
	7'h78 :
		rl_rd00 = rl_rg120 ;
	7'h79 :
		rl_rd00 = rl_rg121 ;
	7'h7a :
		rl_rd00 = rl_rg122 ;
	7'h7b :
		rl_rd00 = rl_rg123 ;
	7'h7c :
		rl_rd00 = rl_rg124 ;
	7'h7d :
		rl_rd00 = rl_rg125 ;
	7'h7e :
		rl_rd00 = rl_rg126 ;
	7'h7f :
		rl_rd00 = rl_rg127 ;
	default :
		rl_rd00 = 9'hx ;
	endcase
jpeg_MEM_zz zz ( .AD1(zz_AD1) ,.RD1(zz_RD1) ,.WD1(zz_WD1) ,.WE1(zz_WE1) ,.CLK1(clk) ,
	.RA2(RG_i[5:0]) ,.RD2(zz_RD2) ,.RA3(6'h00) ,.RD3(zz_RD3) );	// line#=../rle.h:65
assign	M_01 = ~( ( ( rl_we01 & rl_d01 [127] ) | ( rl_we02 & rl_d02 [127] ) ) | ( 
	U_187 & rl_d03 [127] ) ) ;
always @ ( sub12s_91ot or M_01 or U_88 or zz_RD1 or rl_d03 or U_187 or rl_wd02 or 
	rl_d02 or rl_we02 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg00_t_c1 = ( rl_we01 & rl_d01 [127] ) ;	// line#=../rle.cpp:69,85
	rl_rg00_t_c2 = ( rl_we02 & rl_d02 [127] ) ;
	rl_rg00_t_c3 = ( U_187 & rl_d03 [127] ) ;	// line#=../rle.cpp:74
	rl_rg00_t_c4 = ( U_88 & M_01 ) ;	// line#=../rle.cpp:52
	rl_rg00_t = ( ( { 9{ rl_rg00_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg00_t_c3 } } & zz_RD1 )		// line#=../rle.cpp:74
		| ( { 9{ rl_rg00_t_c4 } } & sub12s_91ot )	// line#=../rle.cpp:52
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg00_en = ( rl_rg00_t_c1 | rl_rg00_t_c2 | rl_rg00_t_c3 | rl_rg00_t_c4 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg00 <= 9'h000 ;
	else if ( rl_rg00_en )
		rl_rg00 <= rl_rg00_t ;	// line#=../rle.cpp:23,52,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg01_t_c1 = ( rl_we01 & rl_d01 [126] ) ;	// line#=../rle.cpp:69,85
	rl_rg01_t_c2 = ( rl_we02 & rl_d02 [126] ) ;
	rl_rg01_t_c3 = ( U_187 & rl_d03 [126] ) ;	// line#=../rle.cpp:74
	rl_rg01_t = ( ( { 9{ rl_rg01_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg01_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg01_en = ( rl_rg01_t_c1 | rl_rg01_t_c2 | rl_rg01_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg01 <= 9'h000 ;
	else if ( rl_rg01_en )
		rl_rg01 <= rl_rg01_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg02_t_c1 = ( rl_we01 & rl_d01 [125] ) ;	// line#=../rle.cpp:69,85
	rl_rg02_t_c2 = ( rl_we02 & rl_d02 [125] ) ;
	rl_rg02_t_c3 = ( U_187 & rl_d03 [125] ) ;	// line#=../rle.cpp:74
	rl_rg02_t = ( ( { 9{ rl_rg02_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg02_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg02_en = ( rl_rg02_t_c1 | rl_rg02_t_c2 | rl_rg02_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg02 <= 9'h000 ;
	else if ( rl_rg02_en )
		rl_rg02 <= rl_rg02_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg03_t_c1 = ( rl_we01 & rl_d01 [124] ) ;	// line#=../rle.cpp:69,85
	rl_rg03_t_c2 = ( rl_we02 & rl_d02 [124] ) ;
	rl_rg03_t_c3 = ( U_187 & rl_d03 [124] ) ;	// line#=../rle.cpp:74
	rl_rg03_t = ( ( { 9{ rl_rg03_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg03_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg03_en = ( rl_rg03_t_c1 | rl_rg03_t_c2 | rl_rg03_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg03 <= 9'h000 ;
	else if ( rl_rg03_en )
		rl_rg03 <= rl_rg03_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg04_t_c1 = ( rl_we01 & rl_d01 [123] ) ;	// line#=../rle.cpp:69,85
	rl_rg04_t_c2 = ( rl_we02 & rl_d02 [123] ) ;
	rl_rg04_t_c3 = ( U_187 & rl_d03 [123] ) ;	// line#=../rle.cpp:74
	rl_rg04_t = ( ( { 9{ rl_rg04_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg04_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg04_en = ( rl_rg04_t_c1 | rl_rg04_t_c2 | rl_rg04_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg04 <= 9'h000 ;
	else if ( rl_rg04_en )
		rl_rg04 <= rl_rg04_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg05_t_c1 = ( rl_we01 & rl_d01 [122] ) ;	// line#=../rle.cpp:69,85
	rl_rg05_t_c2 = ( rl_we02 & rl_d02 [122] ) ;
	rl_rg05_t_c3 = ( U_187 & rl_d03 [122] ) ;	// line#=../rle.cpp:74
	rl_rg05_t = ( ( { 9{ rl_rg05_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg05_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg05_en = ( rl_rg05_t_c1 | rl_rg05_t_c2 | rl_rg05_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg05 <= 9'h000 ;
	else if ( rl_rg05_en )
		rl_rg05 <= rl_rg05_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg06_t_c1 = ( rl_we01 & rl_d01 [121] ) ;	// line#=../rle.cpp:69,85
	rl_rg06_t_c2 = ( rl_we02 & rl_d02 [121] ) ;
	rl_rg06_t_c3 = ( U_187 & rl_d03 [121] ) ;	// line#=../rle.cpp:74
	rl_rg06_t = ( ( { 9{ rl_rg06_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg06_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg06_en = ( rl_rg06_t_c1 | rl_rg06_t_c2 | rl_rg06_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg06 <= 9'h000 ;
	else if ( rl_rg06_en )
		rl_rg06 <= rl_rg06_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg07_t_c1 = ( rl_we01 & rl_d01 [120] ) ;	// line#=../rle.cpp:69,85
	rl_rg07_t_c2 = ( rl_we02 & rl_d02 [120] ) ;
	rl_rg07_t_c3 = ( U_187 & rl_d03 [120] ) ;	// line#=../rle.cpp:74
	rl_rg07_t = ( ( { 9{ rl_rg07_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg07_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg07_en = ( rl_rg07_t_c1 | rl_rg07_t_c2 | rl_rg07_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg07 <= 9'h000 ;
	else if ( rl_rg07_en )
		rl_rg07 <= rl_rg07_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg08_t_c1 = ( rl_we01 & rl_d01 [119] ) ;	// line#=../rle.cpp:69,85
	rl_rg08_t_c2 = ( rl_we02 & rl_d02 [119] ) ;
	rl_rg08_t_c3 = ( U_187 & rl_d03 [119] ) ;	// line#=../rle.cpp:74
	rl_rg08_t = ( ( { 9{ rl_rg08_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg08_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg08_en = ( rl_rg08_t_c1 | rl_rg08_t_c2 | rl_rg08_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg08 <= 9'h000 ;
	else if ( rl_rg08_en )
		rl_rg08 <= rl_rg08_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg09_t_c1 = ( rl_we01 & rl_d01 [118] ) ;	// line#=../rle.cpp:69,85
	rl_rg09_t_c2 = ( rl_we02 & rl_d02 [118] ) ;
	rl_rg09_t_c3 = ( U_187 & rl_d03 [118] ) ;	// line#=../rle.cpp:74
	rl_rg09_t = ( ( { 9{ rl_rg09_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg09_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg09_en = ( rl_rg09_t_c1 | rl_rg09_t_c2 | rl_rg09_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg09 <= 9'h000 ;
	else if ( rl_rg09_en )
		rl_rg09 <= rl_rg09_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg10_t_c1 = ( rl_we01 & rl_d01 [117] ) ;	// line#=../rle.cpp:69,85
	rl_rg10_t_c2 = ( rl_we02 & rl_d02 [117] ) ;
	rl_rg10_t_c3 = ( U_187 & rl_d03 [117] ) ;	// line#=../rle.cpp:74
	rl_rg10_t = ( ( { 9{ rl_rg10_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg10_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg10_en = ( rl_rg10_t_c1 | rl_rg10_t_c2 | rl_rg10_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg10 <= 9'h000 ;
	else if ( rl_rg10_en )
		rl_rg10 <= rl_rg10_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg11_t_c1 = ( rl_we01 & rl_d01 [116] ) ;	// line#=../rle.cpp:69,85
	rl_rg11_t_c2 = ( rl_we02 & rl_d02 [116] ) ;
	rl_rg11_t_c3 = ( U_187 & rl_d03 [116] ) ;	// line#=../rle.cpp:74
	rl_rg11_t = ( ( { 9{ rl_rg11_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg11_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg11_en = ( rl_rg11_t_c1 | rl_rg11_t_c2 | rl_rg11_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg11 <= 9'h000 ;
	else if ( rl_rg11_en )
		rl_rg11 <= rl_rg11_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg12_t_c1 = ( rl_we01 & rl_d01 [115] ) ;	// line#=../rle.cpp:69,85
	rl_rg12_t_c2 = ( rl_we02 & rl_d02 [115] ) ;
	rl_rg12_t_c3 = ( U_187 & rl_d03 [115] ) ;	// line#=../rle.cpp:74
	rl_rg12_t = ( ( { 9{ rl_rg12_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg12_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg12_en = ( rl_rg12_t_c1 | rl_rg12_t_c2 | rl_rg12_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg12 <= 9'h000 ;
	else if ( rl_rg12_en )
		rl_rg12 <= rl_rg12_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg13_t_c1 = ( rl_we01 & rl_d01 [114] ) ;	// line#=../rle.cpp:69,85
	rl_rg13_t_c2 = ( rl_we02 & rl_d02 [114] ) ;
	rl_rg13_t_c3 = ( U_187 & rl_d03 [114] ) ;	// line#=../rle.cpp:74
	rl_rg13_t = ( ( { 9{ rl_rg13_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg13_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg13_en = ( rl_rg13_t_c1 | rl_rg13_t_c2 | rl_rg13_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg13 <= 9'h000 ;
	else if ( rl_rg13_en )
		rl_rg13 <= rl_rg13_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg14_t_c1 = ( rl_we01 & rl_d01 [113] ) ;	// line#=../rle.cpp:69,85
	rl_rg14_t_c2 = ( rl_we02 & rl_d02 [113] ) ;
	rl_rg14_t_c3 = ( U_187 & rl_d03 [113] ) ;	// line#=../rle.cpp:74
	rl_rg14_t = ( ( { 9{ rl_rg14_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg14_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg14_en = ( rl_rg14_t_c1 | rl_rg14_t_c2 | rl_rg14_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg14 <= 9'h000 ;
	else if ( rl_rg14_en )
		rl_rg14 <= rl_rg14_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg15_t_c1 = ( rl_we01 & rl_d01 [112] ) ;	// line#=../rle.cpp:69,85
	rl_rg15_t_c2 = ( rl_we02 & rl_d02 [112] ) ;
	rl_rg15_t_c3 = ( U_187 & rl_d03 [112] ) ;	// line#=../rle.cpp:74
	rl_rg15_t = ( ( { 9{ rl_rg15_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg15_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg15_en = ( rl_rg15_t_c1 | rl_rg15_t_c2 | rl_rg15_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg15 <= 9'h000 ;
	else if ( rl_rg15_en )
		rl_rg15 <= rl_rg15_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg16_t_c1 = ( rl_we01 & rl_d01 [111] ) ;	// line#=../rle.cpp:69,85
	rl_rg16_t_c2 = ( rl_we02 & rl_d02 [111] ) ;
	rl_rg16_t_c3 = ( U_187 & rl_d03 [111] ) ;	// line#=../rle.cpp:74
	rl_rg16_t = ( ( { 9{ rl_rg16_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg16_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg16_en = ( rl_rg16_t_c1 | rl_rg16_t_c2 | rl_rg16_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg16 <= 9'h000 ;
	else if ( rl_rg16_en )
		rl_rg16 <= rl_rg16_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg17_t_c1 = ( rl_we01 & rl_d01 [110] ) ;	// line#=../rle.cpp:69,85
	rl_rg17_t_c2 = ( rl_we02 & rl_d02 [110] ) ;
	rl_rg17_t_c3 = ( U_187 & rl_d03 [110] ) ;	// line#=../rle.cpp:74
	rl_rg17_t = ( ( { 9{ rl_rg17_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg17_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg17_en = ( rl_rg17_t_c1 | rl_rg17_t_c2 | rl_rg17_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg17 <= 9'h000 ;
	else if ( rl_rg17_en )
		rl_rg17 <= rl_rg17_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg18_t_c1 = ( rl_we01 & rl_d01 [109] ) ;	// line#=../rle.cpp:69,85
	rl_rg18_t_c2 = ( rl_we02 & rl_d02 [109] ) ;
	rl_rg18_t_c3 = ( U_187 & rl_d03 [109] ) ;	// line#=../rle.cpp:74
	rl_rg18_t = ( ( { 9{ rl_rg18_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg18_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg18_en = ( rl_rg18_t_c1 | rl_rg18_t_c2 | rl_rg18_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg18 <= 9'h000 ;
	else if ( rl_rg18_en )
		rl_rg18 <= rl_rg18_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg19_t_c1 = ( rl_we01 & rl_d01 [108] ) ;	// line#=../rle.cpp:69,85
	rl_rg19_t_c2 = ( rl_we02 & rl_d02 [108] ) ;
	rl_rg19_t_c3 = ( U_187 & rl_d03 [108] ) ;	// line#=../rle.cpp:74
	rl_rg19_t = ( ( { 9{ rl_rg19_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg19_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg19_en = ( rl_rg19_t_c1 | rl_rg19_t_c2 | rl_rg19_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg19 <= 9'h000 ;
	else if ( rl_rg19_en )
		rl_rg19 <= rl_rg19_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg20_t_c1 = ( rl_we01 & rl_d01 [107] ) ;	// line#=../rle.cpp:69,85
	rl_rg20_t_c2 = ( rl_we02 & rl_d02 [107] ) ;
	rl_rg20_t_c3 = ( U_187 & rl_d03 [107] ) ;	// line#=../rle.cpp:74
	rl_rg20_t = ( ( { 9{ rl_rg20_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg20_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg20_en = ( rl_rg20_t_c1 | rl_rg20_t_c2 | rl_rg20_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg20 <= 9'h000 ;
	else if ( rl_rg20_en )
		rl_rg20 <= rl_rg20_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg21_t_c1 = ( rl_we01 & rl_d01 [106] ) ;	// line#=../rle.cpp:69,85
	rl_rg21_t_c2 = ( rl_we02 & rl_d02 [106] ) ;
	rl_rg21_t_c3 = ( U_187 & rl_d03 [106] ) ;	// line#=../rle.cpp:74
	rl_rg21_t = ( ( { 9{ rl_rg21_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg21_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg21_en = ( rl_rg21_t_c1 | rl_rg21_t_c2 | rl_rg21_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg21 <= 9'h000 ;
	else if ( rl_rg21_en )
		rl_rg21 <= rl_rg21_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg22_t_c1 = ( rl_we01 & rl_d01 [105] ) ;	// line#=../rle.cpp:69,85
	rl_rg22_t_c2 = ( rl_we02 & rl_d02 [105] ) ;
	rl_rg22_t_c3 = ( U_187 & rl_d03 [105] ) ;	// line#=../rle.cpp:74
	rl_rg22_t = ( ( { 9{ rl_rg22_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg22_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg22_en = ( rl_rg22_t_c1 | rl_rg22_t_c2 | rl_rg22_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg22 <= 9'h000 ;
	else if ( rl_rg22_en )
		rl_rg22 <= rl_rg22_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg23_t_c1 = ( rl_we01 & rl_d01 [104] ) ;	// line#=../rle.cpp:69,85
	rl_rg23_t_c2 = ( rl_we02 & rl_d02 [104] ) ;
	rl_rg23_t_c3 = ( U_187 & rl_d03 [104] ) ;	// line#=../rle.cpp:74
	rl_rg23_t = ( ( { 9{ rl_rg23_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg23_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg23_en = ( rl_rg23_t_c1 | rl_rg23_t_c2 | rl_rg23_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg23 <= 9'h000 ;
	else if ( rl_rg23_en )
		rl_rg23 <= rl_rg23_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg24_t_c1 = ( rl_we01 & rl_d01 [103] ) ;	// line#=../rle.cpp:69,85
	rl_rg24_t_c2 = ( rl_we02 & rl_d02 [103] ) ;
	rl_rg24_t_c3 = ( U_187 & rl_d03 [103] ) ;	// line#=../rle.cpp:74
	rl_rg24_t = ( ( { 9{ rl_rg24_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg24_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg24_en = ( rl_rg24_t_c1 | rl_rg24_t_c2 | rl_rg24_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg24 <= 9'h000 ;
	else if ( rl_rg24_en )
		rl_rg24 <= rl_rg24_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg25_t_c1 = ( rl_we01 & rl_d01 [102] ) ;	// line#=../rle.cpp:69,85
	rl_rg25_t_c2 = ( rl_we02 & rl_d02 [102] ) ;
	rl_rg25_t_c3 = ( U_187 & rl_d03 [102] ) ;	// line#=../rle.cpp:74
	rl_rg25_t = ( ( { 9{ rl_rg25_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg25_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg25_en = ( rl_rg25_t_c1 | rl_rg25_t_c2 | rl_rg25_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg25 <= 9'h000 ;
	else if ( rl_rg25_en )
		rl_rg25 <= rl_rg25_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg26_t_c1 = ( rl_we01 & rl_d01 [101] ) ;	// line#=../rle.cpp:69,85
	rl_rg26_t_c2 = ( rl_we02 & rl_d02 [101] ) ;
	rl_rg26_t_c3 = ( U_187 & rl_d03 [101] ) ;	// line#=../rle.cpp:74
	rl_rg26_t = ( ( { 9{ rl_rg26_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg26_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg26_en = ( rl_rg26_t_c1 | rl_rg26_t_c2 | rl_rg26_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg26 <= 9'h000 ;
	else if ( rl_rg26_en )
		rl_rg26 <= rl_rg26_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg27_t_c1 = ( rl_we01 & rl_d01 [100] ) ;	// line#=../rle.cpp:69,85
	rl_rg27_t_c2 = ( rl_we02 & rl_d02 [100] ) ;
	rl_rg27_t_c3 = ( U_187 & rl_d03 [100] ) ;	// line#=../rle.cpp:74
	rl_rg27_t = ( ( { 9{ rl_rg27_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg27_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg27_en = ( rl_rg27_t_c1 | rl_rg27_t_c2 | rl_rg27_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg27 <= 9'h000 ;
	else if ( rl_rg27_en )
		rl_rg27 <= rl_rg27_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg28_t_c1 = ( rl_we01 & rl_d01 [99] ) ;	// line#=../rle.cpp:69,85
	rl_rg28_t_c2 = ( rl_we02 & rl_d02 [99] ) ;
	rl_rg28_t_c3 = ( U_187 & rl_d03 [99] ) ;	// line#=../rle.cpp:74
	rl_rg28_t = ( ( { 9{ rl_rg28_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg28_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg28_en = ( rl_rg28_t_c1 | rl_rg28_t_c2 | rl_rg28_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg28 <= 9'h000 ;
	else if ( rl_rg28_en )
		rl_rg28 <= rl_rg28_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg29_t_c1 = ( rl_we01 & rl_d01 [98] ) ;	// line#=../rle.cpp:69,85
	rl_rg29_t_c2 = ( rl_we02 & rl_d02 [98] ) ;
	rl_rg29_t_c3 = ( U_187 & rl_d03 [98] ) ;	// line#=../rle.cpp:74
	rl_rg29_t = ( ( { 9{ rl_rg29_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg29_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg29_en = ( rl_rg29_t_c1 | rl_rg29_t_c2 | rl_rg29_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg29 <= 9'h000 ;
	else if ( rl_rg29_en )
		rl_rg29 <= rl_rg29_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg30_t_c1 = ( rl_we01 & rl_d01 [97] ) ;	// line#=../rle.cpp:69,85
	rl_rg30_t_c2 = ( rl_we02 & rl_d02 [97] ) ;
	rl_rg30_t_c3 = ( U_187 & rl_d03 [97] ) ;	// line#=../rle.cpp:74
	rl_rg30_t = ( ( { 9{ rl_rg30_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg30_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg30_en = ( rl_rg30_t_c1 | rl_rg30_t_c2 | rl_rg30_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg30 <= 9'h000 ;
	else if ( rl_rg30_en )
		rl_rg30 <= rl_rg30_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg31_t_c1 = ( rl_we01 & rl_d01 [96] ) ;	// line#=../rle.cpp:69,85
	rl_rg31_t_c2 = ( rl_we02 & rl_d02 [96] ) ;
	rl_rg31_t_c3 = ( U_187 & rl_d03 [96] ) ;	// line#=../rle.cpp:74
	rl_rg31_t = ( ( { 9{ rl_rg31_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg31_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg31_en = ( rl_rg31_t_c1 | rl_rg31_t_c2 | rl_rg31_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg31 <= 9'h000 ;
	else if ( rl_rg31_en )
		rl_rg31 <= rl_rg31_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg32_t_c1 = ( rl_we01 & rl_d01 [95] ) ;	// line#=../rle.cpp:69,85
	rl_rg32_t_c2 = ( rl_we02 & rl_d02 [95] ) ;
	rl_rg32_t_c3 = ( U_187 & rl_d03 [95] ) ;	// line#=../rle.cpp:74
	rl_rg32_t = ( ( { 9{ rl_rg32_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg32_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg32_en = ( rl_rg32_t_c1 | rl_rg32_t_c2 | rl_rg32_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg32 <= 9'h000 ;
	else if ( rl_rg32_en )
		rl_rg32 <= rl_rg32_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg33_t_c1 = ( rl_we01 & rl_d01 [94] ) ;	// line#=../rle.cpp:69,85
	rl_rg33_t_c2 = ( rl_we02 & rl_d02 [94] ) ;
	rl_rg33_t_c3 = ( U_187 & rl_d03 [94] ) ;	// line#=../rle.cpp:74
	rl_rg33_t = ( ( { 9{ rl_rg33_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg33_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg33_en = ( rl_rg33_t_c1 | rl_rg33_t_c2 | rl_rg33_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg33 <= 9'h000 ;
	else if ( rl_rg33_en )
		rl_rg33 <= rl_rg33_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg34_t_c1 = ( rl_we01 & rl_d01 [93] ) ;	// line#=../rle.cpp:69,85
	rl_rg34_t_c2 = ( rl_we02 & rl_d02 [93] ) ;
	rl_rg34_t_c3 = ( U_187 & rl_d03 [93] ) ;	// line#=../rle.cpp:74
	rl_rg34_t = ( ( { 9{ rl_rg34_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg34_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg34_en = ( rl_rg34_t_c1 | rl_rg34_t_c2 | rl_rg34_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg34 <= 9'h000 ;
	else if ( rl_rg34_en )
		rl_rg34 <= rl_rg34_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg35_t_c1 = ( rl_we01 & rl_d01 [92] ) ;	// line#=../rle.cpp:69,85
	rl_rg35_t_c2 = ( rl_we02 & rl_d02 [92] ) ;
	rl_rg35_t_c3 = ( U_187 & rl_d03 [92] ) ;	// line#=../rle.cpp:74
	rl_rg35_t = ( ( { 9{ rl_rg35_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg35_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg35_en = ( rl_rg35_t_c1 | rl_rg35_t_c2 | rl_rg35_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg35 <= 9'h000 ;
	else if ( rl_rg35_en )
		rl_rg35 <= rl_rg35_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg36_t_c1 = ( rl_we01 & rl_d01 [91] ) ;	// line#=../rle.cpp:69,85
	rl_rg36_t_c2 = ( rl_we02 & rl_d02 [91] ) ;
	rl_rg36_t_c3 = ( U_187 & rl_d03 [91] ) ;	// line#=../rle.cpp:74
	rl_rg36_t = ( ( { 9{ rl_rg36_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg36_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg36_en = ( rl_rg36_t_c1 | rl_rg36_t_c2 | rl_rg36_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg36 <= 9'h000 ;
	else if ( rl_rg36_en )
		rl_rg36 <= rl_rg36_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg37_t_c1 = ( rl_we01 & rl_d01 [90] ) ;	// line#=../rle.cpp:69,85
	rl_rg37_t_c2 = ( rl_we02 & rl_d02 [90] ) ;
	rl_rg37_t_c3 = ( U_187 & rl_d03 [90] ) ;	// line#=../rle.cpp:74
	rl_rg37_t = ( ( { 9{ rl_rg37_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg37_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg37_en = ( rl_rg37_t_c1 | rl_rg37_t_c2 | rl_rg37_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg37 <= 9'h000 ;
	else if ( rl_rg37_en )
		rl_rg37 <= rl_rg37_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg38_t_c1 = ( rl_we01 & rl_d01 [89] ) ;	// line#=../rle.cpp:69,85
	rl_rg38_t_c2 = ( rl_we02 & rl_d02 [89] ) ;
	rl_rg38_t_c3 = ( U_187 & rl_d03 [89] ) ;	// line#=../rle.cpp:74
	rl_rg38_t = ( ( { 9{ rl_rg38_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg38_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg38_en = ( rl_rg38_t_c1 | rl_rg38_t_c2 | rl_rg38_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg38 <= 9'h000 ;
	else if ( rl_rg38_en )
		rl_rg38 <= rl_rg38_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg39_t_c1 = ( rl_we01 & rl_d01 [88] ) ;	// line#=../rle.cpp:69,85
	rl_rg39_t_c2 = ( rl_we02 & rl_d02 [88] ) ;
	rl_rg39_t_c3 = ( U_187 & rl_d03 [88] ) ;	// line#=../rle.cpp:74
	rl_rg39_t = ( ( { 9{ rl_rg39_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg39_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg39_en = ( rl_rg39_t_c1 | rl_rg39_t_c2 | rl_rg39_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg39 <= 9'h000 ;
	else if ( rl_rg39_en )
		rl_rg39 <= rl_rg39_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg40_t_c1 = ( rl_we01 & rl_d01 [87] ) ;	// line#=../rle.cpp:69,85
	rl_rg40_t_c2 = ( rl_we02 & rl_d02 [87] ) ;
	rl_rg40_t_c3 = ( U_187 & rl_d03 [87] ) ;	// line#=../rle.cpp:74
	rl_rg40_t = ( ( { 9{ rl_rg40_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg40_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg40_en = ( rl_rg40_t_c1 | rl_rg40_t_c2 | rl_rg40_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg40 <= 9'h000 ;
	else if ( rl_rg40_en )
		rl_rg40 <= rl_rg40_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg41_t_c1 = ( rl_we01 & rl_d01 [86] ) ;	// line#=../rle.cpp:69,85
	rl_rg41_t_c2 = ( rl_we02 & rl_d02 [86] ) ;
	rl_rg41_t_c3 = ( U_187 & rl_d03 [86] ) ;	// line#=../rle.cpp:74
	rl_rg41_t = ( ( { 9{ rl_rg41_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg41_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg41_en = ( rl_rg41_t_c1 | rl_rg41_t_c2 | rl_rg41_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg41 <= 9'h000 ;
	else if ( rl_rg41_en )
		rl_rg41 <= rl_rg41_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg42_t_c1 = ( rl_we01 & rl_d01 [85] ) ;	// line#=../rle.cpp:69,85
	rl_rg42_t_c2 = ( rl_we02 & rl_d02 [85] ) ;
	rl_rg42_t_c3 = ( U_187 & rl_d03 [85] ) ;	// line#=../rle.cpp:74
	rl_rg42_t = ( ( { 9{ rl_rg42_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg42_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg42_en = ( rl_rg42_t_c1 | rl_rg42_t_c2 | rl_rg42_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg42 <= 9'h000 ;
	else if ( rl_rg42_en )
		rl_rg42 <= rl_rg42_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg43_t_c1 = ( rl_we01 & rl_d01 [84] ) ;	// line#=../rle.cpp:69,85
	rl_rg43_t_c2 = ( rl_we02 & rl_d02 [84] ) ;
	rl_rg43_t_c3 = ( U_187 & rl_d03 [84] ) ;	// line#=../rle.cpp:74
	rl_rg43_t = ( ( { 9{ rl_rg43_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg43_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg43_en = ( rl_rg43_t_c1 | rl_rg43_t_c2 | rl_rg43_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg43 <= 9'h000 ;
	else if ( rl_rg43_en )
		rl_rg43 <= rl_rg43_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg44_t_c1 = ( rl_we01 & rl_d01 [83] ) ;	// line#=../rle.cpp:69,85
	rl_rg44_t_c2 = ( rl_we02 & rl_d02 [83] ) ;
	rl_rg44_t_c3 = ( U_187 & rl_d03 [83] ) ;	// line#=../rle.cpp:74
	rl_rg44_t = ( ( { 9{ rl_rg44_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg44_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg44_en = ( rl_rg44_t_c1 | rl_rg44_t_c2 | rl_rg44_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg44 <= 9'h000 ;
	else if ( rl_rg44_en )
		rl_rg44 <= rl_rg44_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg45_t_c1 = ( rl_we01 & rl_d01 [82] ) ;	// line#=../rle.cpp:69,85
	rl_rg45_t_c2 = ( rl_we02 & rl_d02 [82] ) ;
	rl_rg45_t_c3 = ( U_187 & rl_d03 [82] ) ;	// line#=../rle.cpp:74
	rl_rg45_t = ( ( { 9{ rl_rg45_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg45_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg45_en = ( rl_rg45_t_c1 | rl_rg45_t_c2 | rl_rg45_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg45 <= 9'h000 ;
	else if ( rl_rg45_en )
		rl_rg45 <= rl_rg45_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg46_t_c1 = ( rl_we01 & rl_d01 [81] ) ;	// line#=../rle.cpp:69,85
	rl_rg46_t_c2 = ( rl_we02 & rl_d02 [81] ) ;
	rl_rg46_t_c3 = ( U_187 & rl_d03 [81] ) ;	// line#=../rle.cpp:74
	rl_rg46_t = ( ( { 9{ rl_rg46_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg46_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg46_en = ( rl_rg46_t_c1 | rl_rg46_t_c2 | rl_rg46_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg46 <= 9'h000 ;
	else if ( rl_rg46_en )
		rl_rg46 <= rl_rg46_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg47_t_c1 = ( rl_we01 & rl_d01 [80] ) ;	// line#=../rle.cpp:69,85
	rl_rg47_t_c2 = ( rl_we02 & rl_d02 [80] ) ;
	rl_rg47_t_c3 = ( U_187 & rl_d03 [80] ) ;	// line#=../rle.cpp:74
	rl_rg47_t = ( ( { 9{ rl_rg47_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg47_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg47_en = ( rl_rg47_t_c1 | rl_rg47_t_c2 | rl_rg47_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg47 <= 9'h000 ;
	else if ( rl_rg47_en )
		rl_rg47 <= rl_rg47_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg48_t_c1 = ( rl_we01 & rl_d01 [79] ) ;	// line#=../rle.cpp:69,85
	rl_rg48_t_c2 = ( rl_we02 & rl_d02 [79] ) ;
	rl_rg48_t_c3 = ( U_187 & rl_d03 [79] ) ;	// line#=../rle.cpp:74
	rl_rg48_t = ( ( { 9{ rl_rg48_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg48_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg48_en = ( rl_rg48_t_c1 | rl_rg48_t_c2 | rl_rg48_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg48 <= 9'h000 ;
	else if ( rl_rg48_en )
		rl_rg48 <= rl_rg48_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg49_t_c1 = ( rl_we01 & rl_d01 [78] ) ;	// line#=../rle.cpp:69,85
	rl_rg49_t_c2 = ( rl_we02 & rl_d02 [78] ) ;
	rl_rg49_t_c3 = ( U_187 & rl_d03 [78] ) ;	// line#=../rle.cpp:74
	rl_rg49_t = ( ( { 9{ rl_rg49_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg49_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg49_en = ( rl_rg49_t_c1 | rl_rg49_t_c2 | rl_rg49_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg49 <= 9'h000 ;
	else if ( rl_rg49_en )
		rl_rg49 <= rl_rg49_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg50_t_c1 = ( rl_we01 & rl_d01 [77] ) ;	// line#=../rle.cpp:69,85
	rl_rg50_t_c2 = ( rl_we02 & rl_d02 [77] ) ;
	rl_rg50_t_c3 = ( U_187 & rl_d03 [77] ) ;	// line#=../rle.cpp:74
	rl_rg50_t = ( ( { 9{ rl_rg50_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg50_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg50_en = ( rl_rg50_t_c1 | rl_rg50_t_c2 | rl_rg50_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg50 <= 9'h000 ;
	else if ( rl_rg50_en )
		rl_rg50 <= rl_rg50_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg51_t_c1 = ( rl_we01 & rl_d01 [76] ) ;	// line#=../rle.cpp:69,85
	rl_rg51_t_c2 = ( rl_we02 & rl_d02 [76] ) ;
	rl_rg51_t_c3 = ( U_187 & rl_d03 [76] ) ;	// line#=../rle.cpp:74
	rl_rg51_t = ( ( { 9{ rl_rg51_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg51_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg51_en = ( rl_rg51_t_c1 | rl_rg51_t_c2 | rl_rg51_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg51 <= 9'h000 ;
	else if ( rl_rg51_en )
		rl_rg51 <= rl_rg51_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg52_t_c1 = ( rl_we01 & rl_d01 [75] ) ;	// line#=../rle.cpp:69,85
	rl_rg52_t_c2 = ( rl_we02 & rl_d02 [75] ) ;
	rl_rg52_t_c3 = ( U_187 & rl_d03 [75] ) ;	// line#=../rle.cpp:74
	rl_rg52_t = ( ( { 9{ rl_rg52_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg52_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg52_en = ( rl_rg52_t_c1 | rl_rg52_t_c2 | rl_rg52_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg52 <= 9'h000 ;
	else if ( rl_rg52_en )
		rl_rg52 <= rl_rg52_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg53_t_c1 = ( rl_we01 & rl_d01 [74] ) ;	// line#=../rle.cpp:69,85
	rl_rg53_t_c2 = ( rl_we02 & rl_d02 [74] ) ;
	rl_rg53_t_c3 = ( U_187 & rl_d03 [74] ) ;	// line#=../rle.cpp:74
	rl_rg53_t = ( ( { 9{ rl_rg53_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg53_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg53_en = ( rl_rg53_t_c1 | rl_rg53_t_c2 | rl_rg53_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg53 <= 9'h000 ;
	else if ( rl_rg53_en )
		rl_rg53 <= rl_rg53_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg54_t_c1 = ( rl_we01 & rl_d01 [73] ) ;	// line#=../rle.cpp:69,85
	rl_rg54_t_c2 = ( rl_we02 & rl_d02 [73] ) ;
	rl_rg54_t_c3 = ( U_187 & rl_d03 [73] ) ;	// line#=../rle.cpp:74
	rl_rg54_t = ( ( { 9{ rl_rg54_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg54_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg54_en = ( rl_rg54_t_c1 | rl_rg54_t_c2 | rl_rg54_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg54 <= 9'h000 ;
	else if ( rl_rg54_en )
		rl_rg54 <= rl_rg54_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg55_t_c1 = ( rl_we01 & rl_d01 [72] ) ;	// line#=../rle.cpp:69,85
	rl_rg55_t_c2 = ( rl_we02 & rl_d02 [72] ) ;
	rl_rg55_t_c3 = ( U_187 & rl_d03 [72] ) ;	// line#=../rle.cpp:74
	rl_rg55_t = ( ( { 9{ rl_rg55_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg55_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg55_en = ( rl_rg55_t_c1 | rl_rg55_t_c2 | rl_rg55_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg55 <= 9'h000 ;
	else if ( rl_rg55_en )
		rl_rg55 <= rl_rg55_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg56_t_c1 = ( rl_we01 & rl_d01 [71] ) ;	// line#=../rle.cpp:69,85
	rl_rg56_t_c2 = ( rl_we02 & rl_d02 [71] ) ;
	rl_rg56_t_c3 = ( U_187 & rl_d03 [71] ) ;	// line#=../rle.cpp:74
	rl_rg56_t = ( ( { 9{ rl_rg56_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg56_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg56_en = ( rl_rg56_t_c1 | rl_rg56_t_c2 | rl_rg56_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg56 <= 9'h000 ;
	else if ( rl_rg56_en )
		rl_rg56 <= rl_rg56_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg57_t_c1 = ( rl_we01 & rl_d01 [70] ) ;	// line#=../rle.cpp:69,85
	rl_rg57_t_c2 = ( rl_we02 & rl_d02 [70] ) ;
	rl_rg57_t_c3 = ( U_187 & rl_d03 [70] ) ;	// line#=../rle.cpp:74
	rl_rg57_t = ( ( { 9{ rl_rg57_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg57_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg57_en = ( rl_rg57_t_c1 | rl_rg57_t_c2 | rl_rg57_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg57 <= 9'h000 ;
	else if ( rl_rg57_en )
		rl_rg57 <= rl_rg57_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg58_t_c1 = ( rl_we01 & rl_d01 [69] ) ;	// line#=../rle.cpp:69,85
	rl_rg58_t_c2 = ( rl_we02 & rl_d02 [69] ) ;
	rl_rg58_t_c3 = ( U_187 & rl_d03 [69] ) ;	// line#=../rle.cpp:74
	rl_rg58_t = ( ( { 9{ rl_rg58_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg58_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg58_en = ( rl_rg58_t_c1 | rl_rg58_t_c2 | rl_rg58_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg58 <= 9'h000 ;
	else if ( rl_rg58_en )
		rl_rg58 <= rl_rg58_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg59_t_c1 = ( rl_we01 & rl_d01 [68] ) ;	// line#=../rle.cpp:69,85
	rl_rg59_t_c2 = ( rl_we02 & rl_d02 [68] ) ;
	rl_rg59_t_c3 = ( U_187 & rl_d03 [68] ) ;	// line#=../rle.cpp:74
	rl_rg59_t = ( ( { 9{ rl_rg59_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg59_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg59_en = ( rl_rg59_t_c1 | rl_rg59_t_c2 | rl_rg59_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg59 <= 9'h000 ;
	else if ( rl_rg59_en )
		rl_rg59 <= rl_rg59_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg60_t_c1 = ( rl_we01 & rl_d01 [67] ) ;	// line#=../rle.cpp:69,85
	rl_rg60_t_c2 = ( rl_we02 & rl_d02 [67] ) ;
	rl_rg60_t_c3 = ( U_187 & rl_d03 [67] ) ;	// line#=../rle.cpp:74
	rl_rg60_t = ( ( { 9{ rl_rg60_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg60_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg60_en = ( rl_rg60_t_c1 | rl_rg60_t_c2 | rl_rg60_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg60 <= 9'h000 ;
	else if ( rl_rg60_en )
		rl_rg60 <= rl_rg60_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg61_t_c1 = ( rl_we01 & rl_d01 [66] ) ;	// line#=../rle.cpp:69,85
	rl_rg61_t_c2 = ( rl_we02 & rl_d02 [66] ) ;
	rl_rg61_t_c3 = ( U_187 & rl_d03 [66] ) ;	// line#=../rle.cpp:74
	rl_rg61_t = ( ( { 9{ rl_rg61_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg61_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg61_en = ( rl_rg61_t_c1 | rl_rg61_t_c2 | rl_rg61_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg61 <= 9'h000 ;
	else if ( rl_rg61_en )
		rl_rg61 <= rl_rg61_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg62_t_c1 = ( rl_we01 & rl_d01 [65] ) ;	// line#=../rle.cpp:69,85
	rl_rg62_t_c2 = ( rl_we02 & rl_d02 [65] ) ;
	rl_rg62_t_c3 = ( U_187 & rl_d03 [65] ) ;	// line#=../rle.cpp:74
	rl_rg62_t = ( ( { 9{ rl_rg62_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg62_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg62_en = ( rl_rg62_t_c1 | rl_rg62_t_c2 | rl_rg62_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg62 <= 9'h000 ;
	else if ( rl_rg62_en )
		rl_rg62 <= rl_rg62_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg63_t_c1 = ( rl_we01 & rl_d01 [64] ) ;	// line#=../rle.cpp:69,85
	rl_rg63_t_c2 = ( rl_we02 & rl_d02 [64] ) ;
	rl_rg63_t_c3 = ( U_187 & rl_d03 [64] ) ;	// line#=../rle.cpp:74
	rl_rg63_t = ( ( { 9{ rl_rg63_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg63_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg63_en = ( rl_rg63_t_c1 | rl_rg63_t_c2 | rl_rg63_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg63 <= 9'h000 ;
	else if ( rl_rg63_en )
		rl_rg63 <= rl_rg63_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg64_t_c1 = ( rl_we01 & rl_d01 [63] ) ;	// line#=../rle.cpp:69,85
	rl_rg64_t_c2 = ( rl_we02 & rl_d02 [63] ) ;
	rl_rg64_t_c3 = ( U_187 & rl_d03 [63] ) ;	// line#=../rle.cpp:74
	rl_rg64_t = ( ( { 9{ rl_rg64_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg64_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg64_en = ( rl_rg64_t_c1 | rl_rg64_t_c2 | rl_rg64_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg64 <= 9'h000 ;
	else if ( rl_rg64_en )
		rl_rg64 <= rl_rg64_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg65_t_c1 = ( rl_we01 & rl_d01 [62] ) ;	// line#=../rle.cpp:69,85
	rl_rg65_t_c2 = ( rl_we02 & rl_d02 [62] ) ;
	rl_rg65_t_c3 = ( U_187 & rl_d03 [62] ) ;	// line#=../rle.cpp:74
	rl_rg65_t = ( ( { 9{ rl_rg65_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg65_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg65_en = ( rl_rg65_t_c1 | rl_rg65_t_c2 | rl_rg65_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg65 <= 9'h000 ;
	else if ( rl_rg65_en )
		rl_rg65 <= rl_rg65_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg66_t_c1 = ( rl_we01 & rl_d01 [61] ) ;	// line#=../rle.cpp:69,85
	rl_rg66_t_c2 = ( rl_we02 & rl_d02 [61] ) ;
	rl_rg66_t_c3 = ( U_187 & rl_d03 [61] ) ;	// line#=../rle.cpp:74
	rl_rg66_t = ( ( { 9{ rl_rg66_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg66_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg66_en = ( rl_rg66_t_c1 | rl_rg66_t_c2 | rl_rg66_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg66 <= 9'h000 ;
	else if ( rl_rg66_en )
		rl_rg66 <= rl_rg66_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg67_t_c1 = ( rl_we01 & rl_d01 [60] ) ;	// line#=../rle.cpp:69,85
	rl_rg67_t_c2 = ( rl_we02 & rl_d02 [60] ) ;
	rl_rg67_t_c3 = ( U_187 & rl_d03 [60] ) ;	// line#=../rle.cpp:74
	rl_rg67_t = ( ( { 9{ rl_rg67_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg67_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg67_en = ( rl_rg67_t_c1 | rl_rg67_t_c2 | rl_rg67_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg67 <= 9'h000 ;
	else if ( rl_rg67_en )
		rl_rg67 <= rl_rg67_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg68_t_c1 = ( rl_we01 & rl_d01 [59] ) ;	// line#=../rle.cpp:69,85
	rl_rg68_t_c2 = ( rl_we02 & rl_d02 [59] ) ;
	rl_rg68_t_c3 = ( U_187 & rl_d03 [59] ) ;	// line#=../rle.cpp:74
	rl_rg68_t = ( ( { 9{ rl_rg68_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg68_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg68_en = ( rl_rg68_t_c1 | rl_rg68_t_c2 | rl_rg68_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg68 <= 9'h000 ;
	else if ( rl_rg68_en )
		rl_rg68 <= rl_rg68_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg69_t_c1 = ( rl_we01 & rl_d01 [58] ) ;	// line#=../rle.cpp:69,85
	rl_rg69_t_c2 = ( rl_we02 & rl_d02 [58] ) ;
	rl_rg69_t_c3 = ( U_187 & rl_d03 [58] ) ;	// line#=../rle.cpp:74
	rl_rg69_t = ( ( { 9{ rl_rg69_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg69_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg69_en = ( rl_rg69_t_c1 | rl_rg69_t_c2 | rl_rg69_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg69 <= 9'h000 ;
	else if ( rl_rg69_en )
		rl_rg69 <= rl_rg69_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg70_t_c1 = ( rl_we01 & rl_d01 [57] ) ;	// line#=../rle.cpp:69,85
	rl_rg70_t_c2 = ( rl_we02 & rl_d02 [57] ) ;
	rl_rg70_t_c3 = ( U_187 & rl_d03 [57] ) ;	// line#=../rle.cpp:74
	rl_rg70_t = ( ( { 9{ rl_rg70_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg70_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg70_en = ( rl_rg70_t_c1 | rl_rg70_t_c2 | rl_rg70_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg70 <= 9'h000 ;
	else if ( rl_rg70_en )
		rl_rg70 <= rl_rg70_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg71_t_c1 = ( rl_we01 & rl_d01 [56] ) ;	// line#=../rle.cpp:69,85
	rl_rg71_t_c2 = ( rl_we02 & rl_d02 [56] ) ;
	rl_rg71_t_c3 = ( U_187 & rl_d03 [56] ) ;	// line#=../rle.cpp:74
	rl_rg71_t = ( ( { 9{ rl_rg71_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg71_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg71_en = ( rl_rg71_t_c1 | rl_rg71_t_c2 | rl_rg71_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg71 <= 9'h000 ;
	else if ( rl_rg71_en )
		rl_rg71 <= rl_rg71_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg72_t_c1 = ( rl_we01 & rl_d01 [55] ) ;	// line#=../rle.cpp:69,85
	rl_rg72_t_c2 = ( rl_we02 & rl_d02 [55] ) ;
	rl_rg72_t_c3 = ( U_187 & rl_d03 [55] ) ;	// line#=../rle.cpp:74
	rl_rg72_t = ( ( { 9{ rl_rg72_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg72_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg72_en = ( rl_rg72_t_c1 | rl_rg72_t_c2 | rl_rg72_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg72 <= 9'h000 ;
	else if ( rl_rg72_en )
		rl_rg72 <= rl_rg72_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg73_t_c1 = ( rl_we01 & rl_d01 [54] ) ;	// line#=../rle.cpp:69,85
	rl_rg73_t_c2 = ( rl_we02 & rl_d02 [54] ) ;
	rl_rg73_t_c3 = ( U_187 & rl_d03 [54] ) ;	// line#=../rle.cpp:74
	rl_rg73_t = ( ( { 9{ rl_rg73_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg73_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg73_en = ( rl_rg73_t_c1 | rl_rg73_t_c2 | rl_rg73_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg73 <= 9'h000 ;
	else if ( rl_rg73_en )
		rl_rg73 <= rl_rg73_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg74_t_c1 = ( rl_we01 & rl_d01 [53] ) ;	// line#=../rle.cpp:69,85
	rl_rg74_t_c2 = ( rl_we02 & rl_d02 [53] ) ;
	rl_rg74_t_c3 = ( U_187 & rl_d03 [53] ) ;	// line#=../rle.cpp:74
	rl_rg74_t = ( ( { 9{ rl_rg74_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg74_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg74_en = ( rl_rg74_t_c1 | rl_rg74_t_c2 | rl_rg74_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg74 <= 9'h000 ;
	else if ( rl_rg74_en )
		rl_rg74 <= rl_rg74_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg75_t_c1 = ( rl_we01 & rl_d01 [52] ) ;	// line#=../rle.cpp:69,85
	rl_rg75_t_c2 = ( rl_we02 & rl_d02 [52] ) ;
	rl_rg75_t_c3 = ( U_187 & rl_d03 [52] ) ;	// line#=../rle.cpp:74
	rl_rg75_t = ( ( { 9{ rl_rg75_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg75_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg75_en = ( rl_rg75_t_c1 | rl_rg75_t_c2 | rl_rg75_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg75 <= 9'h000 ;
	else if ( rl_rg75_en )
		rl_rg75 <= rl_rg75_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg76_t_c1 = ( rl_we01 & rl_d01 [51] ) ;	// line#=../rle.cpp:69,85
	rl_rg76_t_c2 = ( rl_we02 & rl_d02 [51] ) ;
	rl_rg76_t_c3 = ( U_187 & rl_d03 [51] ) ;	// line#=../rle.cpp:74
	rl_rg76_t = ( ( { 9{ rl_rg76_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg76_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg76_en = ( rl_rg76_t_c1 | rl_rg76_t_c2 | rl_rg76_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg76 <= 9'h000 ;
	else if ( rl_rg76_en )
		rl_rg76 <= rl_rg76_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg77_t_c1 = ( rl_we01 & rl_d01 [50] ) ;	// line#=../rle.cpp:69,85
	rl_rg77_t_c2 = ( rl_we02 & rl_d02 [50] ) ;
	rl_rg77_t_c3 = ( U_187 & rl_d03 [50] ) ;	// line#=../rle.cpp:74
	rl_rg77_t = ( ( { 9{ rl_rg77_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg77_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg77_en = ( rl_rg77_t_c1 | rl_rg77_t_c2 | rl_rg77_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg77 <= 9'h000 ;
	else if ( rl_rg77_en )
		rl_rg77 <= rl_rg77_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg78_t_c1 = ( rl_we01 & rl_d01 [49] ) ;	// line#=../rle.cpp:69,85
	rl_rg78_t_c2 = ( rl_we02 & rl_d02 [49] ) ;
	rl_rg78_t_c3 = ( U_187 & rl_d03 [49] ) ;	// line#=../rle.cpp:74
	rl_rg78_t = ( ( { 9{ rl_rg78_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg78_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg78_en = ( rl_rg78_t_c1 | rl_rg78_t_c2 | rl_rg78_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg78 <= 9'h000 ;
	else if ( rl_rg78_en )
		rl_rg78 <= rl_rg78_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg79_t_c1 = ( rl_we01 & rl_d01 [48] ) ;	// line#=../rle.cpp:69,85
	rl_rg79_t_c2 = ( rl_we02 & rl_d02 [48] ) ;
	rl_rg79_t_c3 = ( U_187 & rl_d03 [48] ) ;	// line#=../rle.cpp:74
	rl_rg79_t = ( ( { 9{ rl_rg79_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg79_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg79_en = ( rl_rg79_t_c1 | rl_rg79_t_c2 | rl_rg79_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg79 <= 9'h000 ;
	else if ( rl_rg79_en )
		rl_rg79 <= rl_rg79_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg80_t_c1 = ( rl_we01 & rl_d01 [47] ) ;	// line#=../rle.cpp:69,85
	rl_rg80_t_c2 = ( rl_we02 & rl_d02 [47] ) ;
	rl_rg80_t_c3 = ( U_187 & rl_d03 [47] ) ;	// line#=../rle.cpp:74
	rl_rg80_t = ( ( { 9{ rl_rg80_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg80_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg80_en = ( rl_rg80_t_c1 | rl_rg80_t_c2 | rl_rg80_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg80 <= 9'h000 ;
	else if ( rl_rg80_en )
		rl_rg80 <= rl_rg80_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg81_t_c1 = ( rl_we01 & rl_d01 [46] ) ;	// line#=../rle.cpp:69,85
	rl_rg81_t_c2 = ( rl_we02 & rl_d02 [46] ) ;
	rl_rg81_t_c3 = ( U_187 & rl_d03 [46] ) ;	// line#=../rle.cpp:74
	rl_rg81_t = ( ( { 9{ rl_rg81_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg81_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg81_en = ( rl_rg81_t_c1 | rl_rg81_t_c2 | rl_rg81_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg81 <= 9'h000 ;
	else if ( rl_rg81_en )
		rl_rg81 <= rl_rg81_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg82_t_c1 = ( rl_we01 & rl_d01 [45] ) ;	// line#=../rle.cpp:69,85
	rl_rg82_t_c2 = ( rl_we02 & rl_d02 [45] ) ;
	rl_rg82_t_c3 = ( U_187 & rl_d03 [45] ) ;	// line#=../rle.cpp:74
	rl_rg82_t = ( ( { 9{ rl_rg82_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg82_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg82_en = ( rl_rg82_t_c1 | rl_rg82_t_c2 | rl_rg82_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg82 <= 9'h000 ;
	else if ( rl_rg82_en )
		rl_rg82 <= rl_rg82_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg83_t_c1 = ( rl_we01 & rl_d01 [44] ) ;	// line#=../rle.cpp:69,85
	rl_rg83_t_c2 = ( rl_we02 & rl_d02 [44] ) ;
	rl_rg83_t_c3 = ( U_187 & rl_d03 [44] ) ;	// line#=../rle.cpp:74
	rl_rg83_t = ( ( { 9{ rl_rg83_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg83_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg83_en = ( rl_rg83_t_c1 | rl_rg83_t_c2 | rl_rg83_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg83 <= 9'h000 ;
	else if ( rl_rg83_en )
		rl_rg83 <= rl_rg83_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg84_t_c1 = ( rl_we01 & rl_d01 [43] ) ;	// line#=../rle.cpp:69,85
	rl_rg84_t_c2 = ( rl_we02 & rl_d02 [43] ) ;
	rl_rg84_t_c3 = ( U_187 & rl_d03 [43] ) ;	// line#=../rle.cpp:74
	rl_rg84_t = ( ( { 9{ rl_rg84_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg84_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg84_en = ( rl_rg84_t_c1 | rl_rg84_t_c2 | rl_rg84_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg84 <= 9'h000 ;
	else if ( rl_rg84_en )
		rl_rg84 <= rl_rg84_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg85_t_c1 = ( rl_we01 & rl_d01 [42] ) ;	// line#=../rle.cpp:69,85
	rl_rg85_t_c2 = ( rl_we02 & rl_d02 [42] ) ;
	rl_rg85_t_c3 = ( U_187 & rl_d03 [42] ) ;	// line#=../rle.cpp:74
	rl_rg85_t = ( ( { 9{ rl_rg85_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg85_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg85_en = ( rl_rg85_t_c1 | rl_rg85_t_c2 | rl_rg85_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg85 <= 9'h000 ;
	else if ( rl_rg85_en )
		rl_rg85 <= rl_rg85_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg86_t_c1 = ( rl_we01 & rl_d01 [41] ) ;	// line#=../rle.cpp:69,85
	rl_rg86_t_c2 = ( rl_we02 & rl_d02 [41] ) ;
	rl_rg86_t_c3 = ( U_187 & rl_d03 [41] ) ;	// line#=../rle.cpp:74
	rl_rg86_t = ( ( { 9{ rl_rg86_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg86_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg86_en = ( rl_rg86_t_c1 | rl_rg86_t_c2 | rl_rg86_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg86 <= 9'h000 ;
	else if ( rl_rg86_en )
		rl_rg86 <= rl_rg86_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg87_t_c1 = ( rl_we01 & rl_d01 [40] ) ;	// line#=../rle.cpp:69,85
	rl_rg87_t_c2 = ( rl_we02 & rl_d02 [40] ) ;
	rl_rg87_t_c3 = ( U_187 & rl_d03 [40] ) ;	// line#=../rle.cpp:74
	rl_rg87_t = ( ( { 9{ rl_rg87_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg87_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg87_en = ( rl_rg87_t_c1 | rl_rg87_t_c2 | rl_rg87_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg87 <= 9'h000 ;
	else if ( rl_rg87_en )
		rl_rg87 <= rl_rg87_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg88_t_c1 = ( rl_we01 & rl_d01 [39] ) ;	// line#=../rle.cpp:69,85
	rl_rg88_t_c2 = ( rl_we02 & rl_d02 [39] ) ;
	rl_rg88_t_c3 = ( U_187 & rl_d03 [39] ) ;	// line#=../rle.cpp:74
	rl_rg88_t = ( ( { 9{ rl_rg88_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg88_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg88_en = ( rl_rg88_t_c1 | rl_rg88_t_c2 | rl_rg88_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg88 <= 9'h000 ;
	else if ( rl_rg88_en )
		rl_rg88 <= rl_rg88_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg89_t_c1 = ( rl_we01 & rl_d01 [38] ) ;	// line#=../rle.cpp:69,85
	rl_rg89_t_c2 = ( rl_we02 & rl_d02 [38] ) ;
	rl_rg89_t_c3 = ( U_187 & rl_d03 [38] ) ;	// line#=../rle.cpp:74
	rl_rg89_t = ( ( { 9{ rl_rg89_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg89_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg89_en = ( rl_rg89_t_c1 | rl_rg89_t_c2 | rl_rg89_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg89 <= 9'h000 ;
	else if ( rl_rg89_en )
		rl_rg89 <= rl_rg89_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg90_t_c1 = ( rl_we01 & rl_d01 [37] ) ;	// line#=../rle.cpp:69,85
	rl_rg90_t_c2 = ( rl_we02 & rl_d02 [37] ) ;
	rl_rg90_t_c3 = ( U_187 & rl_d03 [37] ) ;	// line#=../rle.cpp:74
	rl_rg90_t = ( ( { 9{ rl_rg90_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg90_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg90_en = ( rl_rg90_t_c1 | rl_rg90_t_c2 | rl_rg90_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg90 <= 9'h000 ;
	else if ( rl_rg90_en )
		rl_rg90 <= rl_rg90_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg91_t_c1 = ( rl_we01 & rl_d01 [36] ) ;	// line#=../rle.cpp:69,85
	rl_rg91_t_c2 = ( rl_we02 & rl_d02 [36] ) ;
	rl_rg91_t_c3 = ( U_187 & rl_d03 [36] ) ;	// line#=../rle.cpp:74
	rl_rg91_t = ( ( { 9{ rl_rg91_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg91_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg91_en = ( rl_rg91_t_c1 | rl_rg91_t_c2 | rl_rg91_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg91 <= 9'h000 ;
	else if ( rl_rg91_en )
		rl_rg91 <= rl_rg91_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg92_t_c1 = ( rl_we01 & rl_d01 [35] ) ;	// line#=../rle.cpp:69,85
	rl_rg92_t_c2 = ( rl_we02 & rl_d02 [35] ) ;
	rl_rg92_t_c3 = ( U_187 & rl_d03 [35] ) ;	// line#=../rle.cpp:74
	rl_rg92_t = ( ( { 9{ rl_rg92_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg92_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg92_en = ( rl_rg92_t_c1 | rl_rg92_t_c2 | rl_rg92_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg92 <= 9'h000 ;
	else if ( rl_rg92_en )
		rl_rg92 <= rl_rg92_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg93_t_c1 = ( rl_we01 & rl_d01 [34] ) ;	// line#=../rle.cpp:69,85
	rl_rg93_t_c2 = ( rl_we02 & rl_d02 [34] ) ;
	rl_rg93_t_c3 = ( U_187 & rl_d03 [34] ) ;	// line#=../rle.cpp:74
	rl_rg93_t = ( ( { 9{ rl_rg93_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg93_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg93_en = ( rl_rg93_t_c1 | rl_rg93_t_c2 | rl_rg93_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg93 <= 9'h000 ;
	else if ( rl_rg93_en )
		rl_rg93 <= rl_rg93_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg94_t_c1 = ( rl_we01 & rl_d01 [33] ) ;	// line#=../rle.cpp:69,85
	rl_rg94_t_c2 = ( rl_we02 & rl_d02 [33] ) ;
	rl_rg94_t_c3 = ( U_187 & rl_d03 [33] ) ;	// line#=../rle.cpp:74
	rl_rg94_t = ( ( { 9{ rl_rg94_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg94_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg94_en = ( rl_rg94_t_c1 | rl_rg94_t_c2 | rl_rg94_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg94 <= 9'h000 ;
	else if ( rl_rg94_en )
		rl_rg94 <= rl_rg94_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg95_t_c1 = ( rl_we01 & rl_d01 [32] ) ;	// line#=../rle.cpp:69,85
	rl_rg95_t_c2 = ( rl_we02 & rl_d02 [32] ) ;
	rl_rg95_t_c3 = ( U_187 & rl_d03 [32] ) ;	// line#=../rle.cpp:74
	rl_rg95_t = ( ( { 9{ rl_rg95_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg95_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg95_en = ( rl_rg95_t_c1 | rl_rg95_t_c2 | rl_rg95_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg95 <= 9'h000 ;
	else if ( rl_rg95_en )
		rl_rg95 <= rl_rg95_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg96_t_c1 = ( rl_we01 & rl_d01 [31] ) ;	// line#=../rle.cpp:69,85
	rl_rg96_t_c2 = ( rl_we02 & rl_d02 [31] ) ;
	rl_rg96_t_c3 = ( U_187 & rl_d03 [31] ) ;	// line#=../rle.cpp:74
	rl_rg96_t = ( ( { 9{ rl_rg96_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg96_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg96_en = ( rl_rg96_t_c1 | rl_rg96_t_c2 | rl_rg96_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg96 <= 9'h000 ;
	else if ( rl_rg96_en )
		rl_rg96 <= rl_rg96_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg97_t_c1 = ( rl_we01 & rl_d01 [30] ) ;	// line#=../rle.cpp:69,85
	rl_rg97_t_c2 = ( rl_we02 & rl_d02 [30] ) ;
	rl_rg97_t_c3 = ( U_187 & rl_d03 [30] ) ;	// line#=../rle.cpp:74
	rl_rg97_t = ( ( { 9{ rl_rg97_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg97_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg97_en = ( rl_rg97_t_c1 | rl_rg97_t_c2 | rl_rg97_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg97 <= 9'h000 ;
	else if ( rl_rg97_en )
		rl_rg97 <= rl_rg97_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg98_t_c1 = ( rl_we01 & rl_d01 [29] ) ;	// line#=../rle.cpp:69,85
	rl_rg98_t_c2 = ( rl_we02 & rl_d02 [29] ) ;
	rl_rg98_t_c3 = ( U_187 & rl_d03 [29] ) ;	// line#=../rle.cpp:74
	rl_rg98_t = ( ( { 9{ rl_rg98_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg98_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg98_en = ( rl_rg98_t_c1 | rl_rg98_t_c2 | rl_rg98_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg98 <= 9'h000 ;
	else if ( rl_rg98_en )
		rl_rg98 <= rl_rg98_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg99_t_c1 = ( rl_we01 & rl_d01 [28] ) ;	// line#=../rle.cpp:69,85
	rl_rg99_t_c2 = ( rl_we02 & rl_d02 [28] ) ;
	rl_rg99_t_c3 = ( U_187 & rl_d03 [28] ) ;	// line#=../rle.cpp:74
	rl_rg99_t = ( ( { 9{ rl_rg99_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg99_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg99_en = ( rl_rg99_t_c1 | rl_rg99_t_c2 | rl_rg99_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg99 <= 9'h000 ;
	else if ( rl_rg99_en )
		rl_rg99 <= rl_rg99_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg100_t_c1 = ( rl_we01 & rl_d01 [27] ) ;	// line#=../rle.cpp:69,85
	rl_rg100_t_c2 = ( rl_we02 & rl_d02 [27] ) ;
	rl_rg100_t_c3 = ( U_187 & rl_d03 [27] ) ;	// line#=../rle.cpp:74
	rl_rg100_t = ( ( { 9{ rl_rg100_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg100_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg100_en = ( rl_rg100_t_c1 | rl_rg100_t_c2 | rl_rg100_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg100 <= 9'h000 ;
	else if ( rl_rg100_en )
		rl_rg100 <= rl_rg100_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg101_t_c1 = ( rl_we01 & rl_d01 [26] ) ;	// line#=../rle.cpp:69,85
	rl_rg101_t_c2 = ( rl_we02 & rl_d02 [26] ) ;
	rl_rg101_t_c3 = ( U_187 & rl_d03 [26] ) ;	// line#=../rle.cpp:74
	rl_rg101_t = ( ( { 9{ rl_rg101_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg101_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg101_en = ( rl_rg101_t_c1 | rl_rg101_t_c2 | rl_rg101_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg101 <= 9'h000 ;
	else if ( rl_rg101_en )
		rl_rg101 <= rl_rg101_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg102_t_c1 = ( rl_we01 & rl_d01 [25] ) ;	// line#=../rle.cpp:69,85
	rl_rg102_t_c2 = ( rl_we02 & rl_d02 [25] ) ;
	rl_rg102_t_c3 = ( U_187 & rl_d03 [25] ) ;	// line#=../rle.cpp:74
	rl_rg102_t = ( ( { 9{ rl_rg102_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg102_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg102_en = ( rl_rg102_t_c1 | rl_rg102_t_c2 | rl_rg102_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg102 <= 9'h000 ;
	else if ( rl_rg102_en )
		rl_rg102 <= rl_rg102_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg103_t_c1 = ( rl_we01 & rl_d01 [24] ) ;	// line#=../rle.cpp:69,85
	rl_rg103_t_c2 = ( rl_we02 & rl_d02 [24] ) ;
	rl_rg103_t_c3 = ( U_187 & rl_d03 [24] ) ;	// line#=../rle.cpp:74
	rl_rg103_t = ( ( { 9{ rl_rg103_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg103_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg103_en = ( rl_rg103_t_c1 | rl_rg103_t_c2 | rl_rg103_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg103 <= 9'h000 ;
	else if ( rl_rg103_en )
		rl_rg103 <= rl_rg103_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg104_t_c1 = ( rl_we01 & rl_d01 [23] ) ;	// line#=../rle.cpp:69,85
	rl_rg104_t_c2 = ( rl_we02 & rl_d02 [23] ) ;
	rl_rg104_t_c3 = ( U_187 & rl_d03 [23] ) ;	// line#=../rle.cpp:74
	rl_rg104_t = ( ( { 9{ rl_rg104_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg104_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg104_en = ( rl_rg104_t_c1 | rl_rg104_t_c2 | rl_rg104_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg104 <= 9'h000 ;
	else if ( rl_rg104_en )
		rl_rg104 <= rl_rg104_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg105_t_c1 = ( rl_we01 & rl_d01 [22] ) ;	// line#=../rle.cpp:69,85
	rl_rg105_t_c2 = ( rl_we02 & rl_d02 [22] ) ;
	rl_rg105_t_c3 = ( U_187 & rl_d03 [22] ) ;	// line#=../rle.cpp:74
	rl_rg105_t = ( ( { 9{ rl_rg105_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg105_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg105_en = ( rl_rg105_t_c1 | rl_rg105_t_c2 | rl_rg105_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg105 <= 9'h000 ;
	else if ( rl_rg105_en )
		rl_rg105 <= rl_rg105_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg106_t_c1 = ( rl_we01 & rl_d01 [21] ) ;	// line#=../rle.cpp:69,85
	rl_rg106_t_c2 = ( rl_we02 & rl_d02 [21] ) ;
	rl_rg106_t_c3 = ( U_187 & rl_d03 [21] ) ;	// line#=../rle.cpp:74
	rl_rg106_t = ( ( { 9{ rl_rg106_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg106_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg106_en = ( rl_rg106_t_c1 | rl_rg106_t_c2 | rl_rg106_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg106 <= 9'h000 ;
	else if ( rl_rg106_en )
		rl_rg106 <= rl_rg106_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg107_t_c1 = ( rl_we01 & rl_d01 [20] ) ;	// line#=../rle.cpp:69,85
	rl_rg107_t_c2 = ( rl_we02 & rl_d02 [20] ) ;
	rl_rg107_t_c3 = ( U_187 & rl_d03 [20] ) ;	// line#=../rle.cpp:74
	rl_rg107_t = ( ( { 9{ rl_rg107_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg107_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg107_en = ( rl_rg107_t_c1 | rl_rg107_t_c2 | rl_rg107_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg107 <= 9'h000 ;
	else if ( rl_rg107_en )
		rl_rg107 <= rl_rg107_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg108_t_c1 = ( rl_we01 & rl_d01 [19] ) ;	// line#=../rle.cpp:69,85
	rl_rg108_t_c2 = ( rl_we02 & rl_d02 [19] ) ;
	rl_rg108_t_c3 = ( U_187 & rl_d03 [19] ) ;	// line#=../rle.cpp:74
	rl_rg108_t = ( ( { 9{ rl_rg108_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg108_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg108_en = ( rl_rg108_t_c1 | rl_rg108_t_c2 | rl_rg108_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg108 <= 9'h000 ;
	else if ( rl_rg108_en )
		rl_rg108 <= rl_rg108_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg109_t_c1 = ( rl_we01 & rl_d01 [18] ) ;	// line#=../rle.cpp:69,85
	rl_rg109_t_c2 = ( rl_we02 & rl_d02 [18] ) ;
	rl_rg109_t_c3 = ( U_187 & rl_d03 [18] ) ;	// line#=../rle.cpp:74
	rl_rg109_t = ( ( { 9{ rl_rg109_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg109_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg109_en = ( rl_rg109_t_c1 | rl_rg109_t_c2 | rl_rg109_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg109 <= 9'h000 ;
	else if ( rl_rg109_en )
		rl_rg109 <= rl_rg109_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg110_t_c1 = ( rl_we01 & rl_d01 [17] ) ;	// line#=../rle.cpp:69,85
	rl_rg110_t_c2 = ( rl_we02 & rl_d02 [17] ) ;
	rl_rg110_t_c3 = ( U_187 & rl_d03 [17] ) ;	// line#=../rle.cpp:74
	rl_rg110_t = ( ( { 9{ rl_rg110_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg110_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg110_en = ( rl_rg110_t_c1 | rl_rg110_t_c2 | rl_rg110_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg110 <= 9'h000 ;
	else if ( rl_rg110_en )
		rl_rg110 <= rl_rg110_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg111_t_c1 = ( rl_we01 & rl_d01 [16] ) ;	// line#=../rle.cpp:69,85
	rl_rg111_t_c2 = ( rl_we02 & rl_d02 [16] ) ;
	rl_rg111_t_c3 = ( U_187 & rl_d03 [16] ) ;	// line#=../rle.cpp:74
	rl_rg111_t = ( ( { 9{ rl_rg111_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg111_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg111_en = ( rl_rg111_t_c1 | rl_rg111_t_c2 | rl_rg111_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg111 <= 9'h000 ;
	else if ( rl_rg111_en )
		rl_rg111 <= rl_rg111_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg112_t_c1 = ( rl_we01 & rl_d01 [15] ) ;	// line#=../rle.cpp:69,85
	rl_rg112_t_c2 = ( rl_we02 & rl_d02 [15] ) ;
	rl_rg112_t_c3 = ( U_187 & rl_d03 [15] ) ;	// line#=../rle.cpp:74
	rl_rg112_t = ( ( { 9{ rl_rg112_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg112_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg112_en = ( rl_rg112_t_c1 | rl_rg112_t_c2 | rl_rg112_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg112 <= 9'h000 ;
	else if ( rl_rg112_en )
		rl_rg112 <= rl_rg112_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg113_t_c1 = ( rl_we01 & rl_d01 [14] ) ;	// line#=../rle.cpp:69,85
	rl_rg113_t_c2 = ( rl_we02 & rl_d02 [14] ) ;
	rl_rg113_t_c3 = ( U_187 & rl_d03 [14] ) ;	// line#=../rle.cpp:74
	rl_rg113_t = ( ( { 9{ rl_rg113_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg113_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg113_en = ( rl_rg113_t_c1 | rl_rg113_t_c2 | rl_rg113_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg113 <= 9'h000 ;
	else if ( rl_rg113_en )
		rl_rg113 <= rl_rg113_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg114_t_c1 = ( rl_we01 & rl_d01 [13] ) ;	// line#=../rle.cpp:69,85
	rl_rg114_t_c2 = ( rl_we02 & rl_d02 [13] ) ;
	rl_rg114_t_c3 = ( U_187 & rl_d03 [13] ) ;	// line#=../rle.cpp:74
	rl_rg114_t = ( ( { 9{ rl_rg114_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg114_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg114_en = ( rl_rg114_t_c1 | rl_rg114_t_c2 | rl_rg114_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg114 <= 9'h000 ;
	else if ( rl_rg114_en )
		rl_rg114 <= rl_rg114_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg115_t_c1 = ( rl_we01 & rl_d01 [12] ) ;	// line#=../rle.cpp:69,85
	rl_rg115_t_c2 = ( rl_we02 & rl_d02 [12] ) ;
	rl_rg115_t_c3 = ( U_187 & rl_d03 [12] ) ;	// line#=../rle.cpp:74
	rl_rg115_t = ( ( { 9{ rl_rg115_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg115_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg115_en = ( rl_rg115_t_c1 | rl_rg115_t_c2 | rl_rg115_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg115 <= 9'h000 ;
	else if ( rl_rg115_en )
		rl_rg115 <= rl_rg115_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg116_t_c1 = ( rl_we01 & rl_d01 [11] ) ;	// line#=../rle.cpp:69,85
	rl_rg116_t_c2 = ( rl_we02 & rl_d02 [11] ) ;
	rl_rg116_t_c3 = ( U_187 & rl_d03 [11] ) ;	// line#=../rle.cpp:74
	rl_rg116_t = ( ( { 9{ rl_rg116_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg116_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg116_en = ( rl_rg116_t_c1 | rl_rg116_t_c2 | rl_rg116_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg116 <= 9'h000 ;
	else if ( rl_rg116_en )
		rl_rg116 <= rl_rg116_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg117_t_c1 = ( rl_we01 & rl_d01 [10] ) ;	// line#=../rle.cpp:69,85
	rl_rg117_t_c2 = ( rl_we02 & rl_d02 [10] ) ;
	rl_rg117_t_c3 = ( U_187 & rl_d03 [10] ) ;	// line#=../rle.cpp:74
	rl_rg117_t = ( ( { 9{ rl_rg117_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg117_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg117_en = ( rl_rg117_t_c1 | rl_rg117_t_c2 | rl_rg117_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg117 <= 9'h000 ;
	else if ( rl_rg117_en )
		rl_rg117 <= rl_rg117_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg118_t_c1 = ( rl_we01 & rl_d01 [9] ) ;	// line#=../rle.cpp:69,85
	rl_rg118_t_c2 = ( rl_we02 & rl_d02 [9] ) ;
	rl_rg118_t_c3 = ( U_187 & rl_d03 [9] ) ;	// line#=../rle.cpp:74
	rl_rg118_t = ( ( { 9{ rl_rg118_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg118_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg118_en = ( rl_rg118_t_c1 | rl_rg118_t_c2 | rl_rg118_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg118 <= 9'h000 ;
	else if ( rl_rg118_en )
		rl_rg118 <= rl_rg118_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg119_t_c1 = ( rl_we01 & rl_d01 [8] ) ;	// line#=../rle.cpp:69,85
	rl_rg119_t_c2 = ( rl_we02 & rl_d02 [8] ) ;
	rl_rg119_t_c3 = ( U_187 & rl_d03 [8] ) ;	// line#=../rle.cpp:74
	rl_rg119_t = ( ( { 9{ rl_rg119_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg119_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg119_en = ( rl_rg119_t_c1 | rl_rg119_t_c2 | rl_rg119_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg119 <= 9'h000 ;
	else if ( rl_rg119_en )
		rl_rg119 <= rl_rg119_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg120_t_c1 = ( rl_we01 & rl_d01 [7] ) ;	// line#=../rle.cpp:69,85
	rl_rg120_t_c2 = ( rl_we02 & rl_d02 [7] ) ;
	rl_rg120_t_c3 = ( U_187 & rl_d03 [7] ) ;	// line#=../rle.cpp:74
	rl_rg120_t = ( ( { 9{ rl_rg120_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg120_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg120_en = ( rl_rg120_t_c1 | rl_rg120_t_c2 | rl_rg120_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg120 <= 9'h000 ;
	else if ( rl_rg120_en )
		rl_rg120 <= rl_rg120_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg121_t_c1 = ( rl_we01 & rl_d01 [6] ) ;	// line#=../rle.cpp:69,85
	rl_rg121_t_c2 = ( rl_we02 & rl_d02 [6] ) ;
	rl_rg121_t_c3 = ( U_187 & rl_d03 [6] ) ;	// line#=../rle.cpp:74
	rl_rg121_t = ( ( { 9{ rl_rg121_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg121_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg121_en = ( rl_rg121_t_c1 | rl_rg121_t_c2 | rl_rg121_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg121 <= 9'h000 ;
	else if ( rl_rg121_en )
		rl_rg121 <= rl_rg121_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg122_t_c1 = ( rl_we01 & rl_d01 [5] ) ;	// line#=../rle.cpp:69,85
	rl_rg122_t_c2 = ( rl_we02 & rl_d02 [5] ) ;
	rl_rg122_t_c3 = ( U_187 & rl_d03 [5] ) ;	// line#=../rle.cpp:74
	rl_rg122_t = ( ( { 9{ rl_rg122_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg122_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg122_en = ( rl_rg122_t_c1 | rl_rg122_t_c2 | rl_rg122_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg122 <= 9'h000 ;
	else if ( rl_rg122_en )
		rl_rg122 <= rl_rg122_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg123_t_c1 = ( rl_we01 & rl_d01 [4] ) ;	// line#=../rle.cpp:69,85
	rl_rg123_t_c2 = ( rl_we02 & rl_d02 [4] ) ;
	rl_rg123_t_c3 = ( U_187 & rl_d03 [4] ) ;	// line#=../rle.cpp:74
	rl_rg123_t = ( ( { 9{ rl_rg123_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg123_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg123_en = ( rl_rg123_t_c1 | rl_rg123_t_c2 | rl_rg123_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg123 <= 9'h000 ;
	else if ( rl_rg123_en )
		rl_rg123 <= rl_rg123_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg124_t_c1 = ( rl_we01 & rl_d01 [3] ) ;	// line#=../rle.cpp:69,85
	rl_rg124_t_c2 = ( rl_we02 & rl_d02 [3] ) ;
	rl_rg124_t_c3 = ( U_187 & rl_d03 [3] ) ;	// line#=../rle.cpp:74
	rl_rg124_t = ( ( { 9{ rl_rg124_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg124_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg124_en = ( rl_rg124_t_c1 | rl_rg124_t_c2 | rl_rg124_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg124 <= 9'h000 ;
	else if ( rl_rg124_en )
		rl_rg124 <= rl_rg124_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg125_t_c1 = ( rl_we01 & rl_d01 [2] ) ;	// line#=../rle.cpp:69,85
	rl_rg125_t_c2 = ( rl_we02 & rl_d02 [2] ) ;
	rl_rg125_t_c3 = ( U_187 & rl_d03 [2] ) ;	// line#=../rle.cpp:74
	rl_rg125_t = ( ( { 9{ rl_rg125_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg125_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg125_en = ( rl_rg125_t_c1 | rl_rg125_t_c2 | rl_rg125_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg125 <= 9'h000 ;
	else if ( rl_rg125_en )
		rl_rg125 <= rl_rg125_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg126_t_c1 = ( rl_we01 & rl_d01 [1] ) ;	// line#=../rle.cpp:69,85
	rl_rg126_t_c2 = ( rl_we02 & rl_d02 [1] ) ;
	rl_rg126_t_c3 = ( U_187 & rl_d03 [1] ) ;	// line#=../rle.cpp:74
	rl_rg126_t = ( ( { 9{ rl_rg126_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg126_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg126_en = ( rl_rg126_t_c1 | rl_rg126_t_c2 | rl_rg126_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg126 <= 9'h000 ;
	else if ( rl_rg126_en )
		rl_rg126 <= rl_rg126_t ;	// line#=../rle.cpp:23,69,74,85
always @ ( zz_RD1 or rl_d03 or U_187 or rl_wd02 or rl_d02 or rl_we02 or rl_d01 or 
	rl_we01 )	// line#=../rle.cpp:23,74
	begin
	rl_rg127_t_c1 = ( rl_we01 & rl_d01 [0] ) ;	// line#=../rle.cpp:69,85
	rl_rg127_t_c2 = ( rl_we02 & rl_d02 [0] ) ;
	rl_rg127_t_c3 = ( U_187 & rl_d03 [0] ) ;	// line#=../rle.cpp:74
	rl_rg127_t = ( ( { 9{ rl_rg127_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg127_t_c3 } } & zz_RD1 )	// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:69,85
	end
assign	rl_rg127_en = ( rl_rg127_t_c1 | rl_rg127_t_c2 | rl_rg127_t_c3 ) ;	// line#=../rle.cpp:23,74
always @ ( posedge clk )	// line#=../rle.cpp:23,74
	if ( !rst )
		rl_rg127 <= 9'h000 ;
	else if ( rl_rg127_en )
		rl_rg127 <= rl_rg127_t ;	// line#=../rle.cpp:23,69,74,85
assign	CT_12 = ( ( ~|RG_j_k ) & M_102 ) ;	// line#=../rle.cpp:117,118
assign	M_102 = ~|{ ( RG_i [31] & RG_i [0] ) , ~RG_i [0] } ;	// line#=../rle.cpp:117,118,148,149
assign	CT_26 = ( ( ~|{ RG_j_k [31:3] , ~RG_j_k [2:0] } ) & M_102 ) ;	// line#=../rle.cpp:148,149
always @ ( RG_zz_02 or FF_d_02 )	// line#=../rle.cpp:61,62
	case ( FF_d_02 )
	1'h1 :
		M_01_t1 = ~|RG_zz_02 ;	// line#=../rle.cpp:61,62
	1'h0 :
		M_01_t1 = 1'h0 ;	// line#=../rle.cpp:61,62
	default :
		M_01_t1 = 1'hx ;
	endcase
assign	CT_31 = ~|{ RG_i_04 [31:7] , ~RG_i_04 [6] , RG_i_04 [5:0] } ;	// line#=../rle.cpp:66,67
assign	CT_32 = ~|rl_rd00 ;	// line#=../rle.cpp:77,78,83,84
always @ ( CT_32 )	// line#=../rle.cpp:77,78
	case ( CT_32 )
	1'h1 :
		JF_06 = 1'h1 ;
	1'h0 :
		JF_06 = 1'h0 ;
	default :
		JF_06 = 1'hx ;
	endcase
always @ ( CT_32 or RG_76_05 )	// line#=../rle.cpp:83,84
	case ( RG_76_05 )
	1'h1 :
		CT_35 = CT_32 ;	// line#=../rle.cpp:83,84
	1'h0 :
		CT_35 = 1'h0 ;	// line#=../rle.cpp:83,84
	default :
		CT_35 = 1'hx ;
	endcase
assign	FL01_01_Leos_all = ( ( ( ( FL01_01_eos & FL01_02_Leos ) & FL01_04_eos ) & 
	FL01_05_eos ) & FL01_06_eos ) ;
assign	FL01_02_Leos_all = ( FL01_02_eos & FL01_03_eos ) ;
assign	FL01_02_rdy = 1'h1 ;
assign	sub12s_91i1 = zz_RD3 ;	// line#=../rle.cpp:52,53
assign	sub12s_91i2 = RG_previous_dc ;	// line#=../rle.cpp:52
assign	lop8u_11i1 = RG_k ;	// line#=../rle.cpp:109,110
assign	lop8u_11i2 = 6'h24 ;	// line#=../rle.cpp:109,110
assign	incr4s1i1 = RG_j ;	// line#=../rle.cpp:34
assign	incr32s3i1 = RG_i_05 ;	// line#=../rle.cpp:74
assign	decr8u_71i1 = RG_len_05 [6:0] ;	// line#=../rle.cpp:77,78
assign	incr8u_71i1 = RG_k_05 [5:0] ;	// line#=../rle.cpp:142
assign	incr8u_61i1 = RG_k ;	// line#=../rle.cpp:111
assign	rl_ad03 = RG_k_05 ;	// line#=../rle.cpp:74
assign	U_05 = ( ST1_03d & lop8u_11ot ) ;	// line#=../rle.cpp:109,110
assign	U_06 = ( ST1_03d & ( ~lop8u_11ot ) ) ;	// line#=../rle.cpp:109,110
assign	U_07 = ( U_05 & M_107 ) ;	// line#=../rle.cpp:111
assign	U_08 = ( U_05 & M_103 ) ;	// line#=../rle.cpp:111
assign	U_09 = ( U_05 & M_112 ) ;	// line#=../rle.cpp:111
assign	U_10 = ( U_05 & M_119 ) ;	// line#=../rle.cpp:111
assign	U_11 = ( U_05 & M_117 ) ;	// line#=../rle.cpp:111
assign	U_12 = ( U_05 & M_122 ) ;	// line#=../rle.cpp:111
assign	U_13 = ( U_05 & M_124 ) ;	// line#=../rle.cpp:111
assign	U_14 = ( U_05 & M_115 ) ;	// line#=../rle.cpp:111
assign	C_02 = ( ( ~|RG_i ) & M_126 ) ;	// line#=../rle.cpp:112,113
assign	U_79 = ( U_05 & C_02 ) ;	// line#=../rle.cpp:112,113
assign	U_80 = ( U_05 & ( ~C_02 ) ) ;	// line#=../rle.cpp:112,113
assign	U_81 = ( U_80 & CT_12 ) ;	// line#=../rle.cpp:117,118
assign	U_82 = ( U_80 & ( ~CT_12 ) ) ;	// line#=../rle.cpp:117,118
assign	U_83 = ( U_82 & ( ~FF_d_02 ) ) ;	// line#=../rle.cpp:122,123
assign	U_84 = ( U_82 & FF_d_02 ) ;	// line#=../rle.cpp:122,123
assign	U_87 = ( ST1_04d & ( ~RG_k_05 [6] ) ) ;	// line#=../rle.cpp:140,141
assign	U_88 = ( ST1_04d & RG_k_05 [6] ) ;	// line#=../rle.cpp:140,141
assign	M_107 = ~|RG_i [2:0] ;	// line#=../rle.cpp:111,142
assign	U_89 = ( U_87 & M_107 ) ;	// line#=../rle.cpp:142
assign	M_103 = ~|( RG_i [2:0] ^ 3'h1 ) ;	// line#=../rle.cpp:111,142
assign	U_90 = ( U_87 & M_103 ) ;	// line#=../rle.cpp:142
assign	M_112 = ~|( RG_i [2:0] ^ 3'h2 ) ;	// line#=../rle.cpp:111,142
assign	U_91 = ( U_87 & M_112 ) ;	// line#=../rle.cpp:142
assign	M_119 = ~|( RG_i [2:0] ^ 3'h3 ) ;	// line#=../rle.cpp:111,142
assign	U_92 = ( U_87 & M_119 ) ;	// line#=../rle.cpp:142
assign	M_117 = ~|( RG_i [2:0] ^ 3'h4 ) ;	// line#=../rle.cpp:111,142
assign	U_93 = ( U_87 & M_117 ) ;	// line#=../rle.cpp:142
assign	M_122 = ~|( RG_i [2:0] ^ 3'h5 ) ;	// line#=../rle.cpp:111,142
assign	U_94 = ( U_87 & M_122 ) ;	// line#=../rle.cpp:142
assign	M_124 = ~|( RG_i [2:0] ^ 3'h6 ) ;	// line#=../rle.cpp:111,142
assign	U_95 = ( U_87 & M_124 ) ;	// line#=../rle.cpp:142
assign	M_115 = ~|( RG_i [2:0] ^ 3'h7 ) ;	// line#=../rle.cpp:111,142
assign	U_96 = ( U_87 & M_115 ) ;	// line#=../rle.cpp:142
assign	M_126 = ~|{ ( RG_j_k [31] & RG_j_k [0] ) , RG_j_k [0] } ;	// line#=../rle.cpp:112,113,143,144
assign	C_05 = ( ( ~|{ RG_i [31:3] , ~RG_i [2:0] } ) & M_126 ) ;	// line#=../rle.cpp:143,144
assign	U_161 = ( U_87 & C_05 ) ;	// line#=../rle.cpp:143,144
assign	U_162 = ( U_87 & ( ~C_05 ) ) ;	// line#=../rle.cpp:143,144
assign	U_163 = ( U_162 & CT_26 ) ;	// line#=../rle.cpp:148,149
assign	U_164 = ( U_162 & ( ~CT_26 ) ) ;	// line#=../rle.cpp:148,149
assign	U_165 = ( U_164 & ( ~FF_d_02 ) ) ;	// line#=../rle.cpp:153,154
assign	U_166 = ( U_164 & FF_d_02 ) ;	// line#=../rle.cpp:153,154
assign	U_168 = ( ST1_04d & ( ~JF_03 ) ) ;
assign	U_169 = ( ST1_05d & FL01_01_01a ) ;
assign	C_07 = ( RG_i_06 [31] | ( ~|RG_i_06 [30:6] ) ) ;	// line#=../rle.cpp:57,58
assign	U_170 = ( U_169 & C_07 ) ;	// line#=../rle.cpp:57,58
assign	U_173 = ( ST1_05d & FL01_02_01a ) ;
assign	U_176 = ( ST1_05d & FL01_03_01a ) ;
assign	U_180 = ( ST1_05d & FL01_04_01a ) ;
assign	U_181 = ( ST1_05d & FL01_05_01a ) ;
assign	U_182 = ( U_181 & CT_31 ) ;	// line#=../rle.cpp:66,67
assign	U_183 = ( U_181 & ( ~CT_31 ) ) ;	// line#=../rle.cpp:66,67
assign	U_185 = ( ST1_05d & FL01_06_01a ) ;
assign	U_186 = ( U_185 & RG_76_05 ) ;	// line#=../rle.cpp:66,67
assign	U_187 = ( U_185 & ( ~RG_76_05 ) ) ;	// line#=../rle.cpp:66,67
assign	U_188 = ( ST1_05d & ( ~|( FL01_01_streg ^ 2'h2 ) ) ) ;
assign	U_190 = ( ST1_05d & M_105 ) ;
assign	U_192 = ( U_188 & ( ~FL01_02_Lrdy ) ) ;
assign	C_11 = ( flag_r1 & flag_r2 ) ;
assign	U_195 = ( U_190 & C_11 ) ;
assign	U_198 = ( U_195 & ( ~FJ_05_11 ) ) ;
assign	U_200 = ( U_198 & ( ~FL01_02_Lrdy ) ) ;
assign	U_204 = ( ST1_05d & ( ~|( FL01_02_streg ^ 2'h1 ) ) ) ;
assign	U_205 = ( ST1_05d & ( ~|( FL01_02_streg ^ 2'h2 ) ) ) ;
assign	U_206 = ( ST1_05d & ( ~|( FL01_02_streg ^ 2'h3 ) ) ) ;
assign	U_207 = ( ( ST1_05d & ( ~|FL01_02_streg ) ) & flag_r3 ) ;
assign	U_208 = ( U_207 & FL01_01_ndat ) ;
assign	U_209 = ( U_207 & ( ~FL01_01_ndat ) ) ;
assign	U_212 = ( U_205 & FL01_02_Leos_all ) ;
assign	U_215 = ( U_212 & ( ~FL01_04_rdy ) ) ;
assign	U_216 = ( ST1_05d & ( ~FL01_03_streg ) ) ;
assign	U_217 = ( ST1_05d & FL01_03_streg ) ;
assign	U_221 = ( U_217 & ( ~FJ_07_08 ) ) ;
assign	U_224 = ( ST1_05d & ( ~FL01_04_streg ) ) ;
assign	U_225 = ( ST1_05d & FL01_04_streg ) ;
assign	U_228 = ( U_225 & FL01_02_Lndat ) ;
assign	U_230 = ( ST1_05d & ( ~FL01_05_streg ) ) ;
assign	U_231 = ( ST1_05d & FL01_05_streg ) ;
assign	U_236 = ( ST1_05d & ( ~FL01_06_streg ) ) ;
assign	U_237 = ( ST1_05d & FL01_06_streg ) ;
assign	U_242 = ( ST1_05d & FL01_01_break ) ;
assign	U_246 = ( ST1_05d & FL01_03_break ) ;
assign	U_258 = ( ST1_08d & ( ~FF_d_02 ) ) ;	// line#=../rle.cpp:77,78
assign	U_263 = ( ST1_11d & ( ~CT_35 ) ) ;	// line#=../rle.cpp:83,84
assign	U_264 = ( ST1_11d & RG_76_05 ) ;	// line#=../rle.cpp:83,84
assign	RG_previous_dc_en = ST1_11d ;
always @ ( posedge clk )
	if ( !rst )
		RG_previous_dc <= 9'h000 ;
	else if ( RG_previous_dc_en )
		RG_previous_dc <= RG_previous_dc_quantized_block ;
always @ ( FF_j or ST1_11d or incr4s1ot or ST1_02d or ST1_01d )
	RG_j_t = ( ( { 4{ ST1_01d } } & 4'hf /*-4'h1*/ )	// line#=../rle.cpp:34
		| ( { 4{ ST1_02d } } & incr4s1ot )		// line#=../rle.cpp:34
		| ( { 4{ ST1_11d } } & { 3'h0 , FF_j } ) ) ;
always @ ( posedge clk )
	RG_j <= RG_j_t ;	// line#=../rle.cpp:34
always @ ( incr32s3ot or U_187 or RG_i_05 or U_186 or U_185 or ST1_02d )
	begin
	RG_i_06_t_c1 = ( U_185 & U_186 ) ;
	RG_i_06_t_c2 = ( U_185 & U_187 ) ;	// line#=../rle.cpp:74
	RG_i_06_t = ( ( { 32{ ST1_02d } } & 32'h00000001 )	// line#=../rle.cpp:37
		| ( { 32{ RG_i_06_t_c1 } } & RG_i_05 )
		| ( { 32{ RG_i_06_t_c2 } } & incr32s3ot )	// line#=../rle.cpp:74
		) ;
	end
assign	RG_i_06_en = ( ST1_02d | RG_i_06_t_c1 | RG_i_06_t_c2 ) ;
always @ ( posedge clk )
	if ( RG_i_06_en )
		RG_i_06 <= RG_i_06_t ;	// line#=../rle.cpp:37,74
always @ ( U_06 )
	TR_01 = ( { 3{ U_06 } } & 3'h7 )	// line#=../rle.cpp:134
		 ;	// line#=../rle.cpp:105
always @ ( RG_i_06 or U_170 or decr32s1ot or U_165 or U_83 or incr32s2ot or U_173 or 
	U_166 or U_163 or U_84 or U_81 or TR_01 or M_129 )
	begin
	RG_i_t_c1 = ( ( ( ( U_81 | U_84 ) | U_163 ) | U_166 ) | U_173 ) ;	// line#=../rle.cpp:61,62,63,119,129,150
										// ,160
	RG_i_t_c2 = ( U_83 | U_165 ) ;	// line#=../rle.cpp:124,155
	RG_i_t = ( ( { 32{ M_129 } } & { 29'h00000000 , TR_01 } )	// line#=../rle.cpp:105,134
		| ( { 32{ RG_i_t_c1 } } & incr32s2ot )			// line#=../rle.cpp:61,62,63,119,129,150
									// ,160
		| ( { 32{ RG_i_t_c2 } } & decr32s1ot )			// line#=../rle.cpp:124,155
		| ( { 32{ U_170 } } & RG_i_06 ) ) ;
	end
assign	RG_i_en = ( M_129 | RG_i_t_c1 | RG_i_t_c2 | U_170 ) ;
always @ ( posedge clk )
	if ( RG_i_en )
		RG_i <= RG_i_t ;	// line#=../rle.cpp:61,62,63,105,119,124
					// ,129,134,150,155,160
always @ ( decr32s2ot or U_166 or U_84 or incr32s1ot or U_173 or U_165 or U_161 or 
	U_83 or U_79 or U_06 or U_170 or ST1_02d )
	begin
	RG_j_k_t_c1 = ( ( ST1_02d | U_170 ) | U_06 ) ;	// line#=../rle.cpp:59,105,135
	RG_j_k_t_c2 = ( ( ( ( U_79 | U_83 ) | U_161 ) | U_165 ) | U_173 ) ;	// line#=../rle.cpp:64,114,125,145,156
	RG_j_k_t_c3 = ( U_84 | U_166 ) ;	// line#=../rle.cpp:130,161
	RG_j_k_t = ( ( { 32{ RG_j_k_t_c1 } } & { 31'h00000000 , U_06 } )	// line#=../rle.cpp:59,105,135
		| ( { 32{ RG_j_k_t_c2 } } & incr32s1ot )			// line#=../rle.cpp:64,114,125,145,156
		| ( { 32{ RG_j_k_t_c3 } } & decr32s2ot )			// line#=../rle.cpp:130,161
		) ;
	end
assign	RG_j_k_en = ( RG_j_k_t_c1 | RG_j_k_t_c2 | RG_j_k_t_c3 ) ;
always @ ( posedge clk )
	if ( RG_j_k_en )
		RG_j_k <= RG_j_k_t ;	// line#=../rle.cpp:59,64,105,114,125,130
					// ,135,145,156,161
assign	RG_quantized_block_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_en )
		RG_quantized_block <= jpeg_in_a00 ;
assign	RG_quantized_block_1_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_1_en )
		RG_quantized_block_1 <= jpeg_in_a01 ;
assign	RG_quantized_block_2_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_2_en )
		RG_quantized_block_2 <= jpeg_in_a02 ;
assign	RG_quantized_block_3_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_3_en )
		RG_quantized_block_3 <= jpeg_in_a03 ;
assign	RG_quantized_block_4_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_4_en )
		RG_quantized_block_4 <= jpeg_in_a04 ;
assign	RG_quantized_block_5_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_5_en )
		RG_quantized_block_5 <= jpeg_in_a05 ;
assign	RG_quantized_block_6_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_6_en )
		RG_quantized_block_6 <= jpeg_in_a06 ;
assign	RG_quantized_block_7_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_7_en )
		RG_quantized_block_7 <= jpeg_in_a07 ;
assign	RG_quantized_block_8_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_8_en )
		RG_quantized_block_8 <= jpeg_in_a08 ;
assign	RG_quantized_block_9_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_9_en )
		RG_quantized_block_9 <= jpeg_in_a09 ;
assign	RG_quantized_block_10_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_10_en )
		RG_quantized_block_10 <= jpeg_in_a10 ;
assign	RG_quantized_block_11_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_11_en )
		RG_quantized_block_11 <= jpeg_in_a11 ;
assign	RG_quantized_block_12_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_12_en )
		RG_quantized_block_12 <= jpeg_in_a12 ;
assign	RG_quantized_block_13_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_13_en )
		RG_quantized_block_13 <= jpeg_in_a13 ;
assign	RG_quantized_block_14_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_14_en )
		RG_quantized_block_14 <= jpeg_in_a14 ;
assign	RG_quantized_block_15_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_15_en )
		RG_quantized_block_15 <= jpeg_in_a15 ;
assign	RG_quantized_block_16_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_16_en )
		RG_quantized_block_16 <= jpeg_in_a16 ;
assign	RG_quantized_block_17_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_17_en )
		RG_quantized_block_17 <= jpeg_in_a17 ;
assign	RG_quantized_block_18_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_18_en )
		RG_quantized_block_18 <= jpeg_in_a18 ;
assign	RG_quantized_block_19_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_19_en )
		RG_quantized_block_19 <= jpeg_in_a19 ;
assign	RG_quantized_block_20_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_20_en )
		RG_quantized_block_20 <= jpeg_in_a20 ;
assign	RG_quantized_block_21_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_21_en )
		RG_quantized_block_21 <= jpeg_in_a21 ;
assign	RG_quantized_block_22_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_22_en )
		RG_quantized_block_22 <= jpeg_in_a22 ;
assign	RG_quantized_block_23_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_23_en )
		RG_quantized_block_23 <= jpeg_in_a23 ;
assign	RG_quantized_block_24_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_24_en )
		RG_quantized_block_24 <= jpeg_in_a24 ;
assign	RG_quantized_block_25_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_25_en )
		RG_quantized_block_25 <= jpeg_in_a25 ;
assign	RG_quantized_block_26_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_26_en )
		RG_quantized_block_26 <= jpeg_in_a26 ;
assign	RG_quantized_block_27_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_27_en )
		RG_quantized_block_27 <= jpeg_in_a27 ;
assign	RG_quantized_block_28_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_28_en )
		RG_quantized_block_28 <= jpeg_in_a28 ;
assign	RG_quantized_block_29_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_29_en )
		RG_quantized_block_29 <= jpeg_in_a29 ;
assign	RG_quantized_block_30_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_30_en )
		RG_quantized_block_30 <= jpeg_in_a30 ;
assign	RG_quantized_block_31_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_31_en )
		RG_quantized_block_31 <= jpeg_in_a31 ;
assign	RG_quantized_block_32_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_32_en )
		RG_quantized_block_32 <= jpeg_in_a32 ;
assign	RG_quantized_block_33_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_33_en )
		RG_quantized_block_33 <= jpeg_in_a33 ;
assign	RG_quantized_block_34_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_34_en )
		RG_quantized_block_34 <= jpeg_in_a34 ;
assign	RG_quantized_block_35_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_35_en )
		RG_quantized_block_35 <= jpeg_in_a35 ;
assign	RG_quantized_block_36_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_36_en )
		RG_quantized_block_36 <= jpeg_in_a36 ;
assign	RG_quantized_block_37_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_37_en )
		RG_quantized_block_37 <= jpeg_in_a37 ;
assign	RG_quantized_block_38_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_38_en )
		RG_quantized_block_38 <= jpeg_in_a38 ;
assign	RG_quantized_block_39_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_39_en )
		RG_quantized_block_39 <= jpeg_in_a39 ;
assign	RG_quantized_block_40_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_40_en )
		RG_quantized_block_40 <= jpeg_in_a40 ;
assign	RG_quantized_block_41_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_41_en )
		RG_quantized_block_41 <= jpeg_in_a41 ;
assign	RG_quantized_block_42_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_42_en )
		RG_quantized_block_42 <= jpeg_in_a42 ;
assign	RG_quantized_block_43_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_43_en )
		RG_quantized_block_43 <= jpeg_in_a43 ;
assign	RG_quantized_block_44_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_44_en )
		RG_quantized_block_44 <= jpeg_in_a44 ;
assign	RG_quantized_block_45_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_45_en )
		RG_quantized_block_45 <= jpeg_in_a45 ;
assign	RG_quantized_block_46_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_46_en )
		RG_quantized_block_46 <= jpeg_in_a46 ;
assign	RG_quantized_block_47_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_47_en )
		RG_quantized_block_47 <= jpeg_in_a47 ;
assign	RG_quantized_block_48_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_48_en )
		RG_quantized_block_48 <= jpeg_in_a48 ;
assign	RG_quantized_block_49_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_49_en )
		RG_quantized_block_49 <= jpeg_in_a49 ;
assign	RG_quantized_block_50_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_50_en )
		RG_quantized_block_50 <= jpeg_in_a50 ;
assign	RG_quantized_block_51_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_51_en )
		RG_quantized_block_51 <= jpeg_in_a51 ;
assign	RG_quantized_block_52_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_52_en )
		RG_quantized_block_52 <= jpeg_in_a52 ;
assign	RG_quantized_block_53_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_53_en )
		RG_quantized_block_53 <= jpeg_in_a53 ;
assign	RG_quantized_block_54_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_54_en )
		RG_quantized_block_54 <= jpeg_in_a54 ;
assign	RG_quantized_block_55_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_55_en )
		RG_quantized_block_55 <= jpeg_in_a55 ;
assign	RG_quantized_block_56_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_56_en )
		RG_quantized_block_56 <= jpeg_in_a56 ;
assign	RG_quantized_block_57_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_57_en )
		RG_quantized_block_57 <= jpeg_in_a57 ;
assign	RG_quantized_block_58_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_58_en )
		RG_quantized_block_58 <= jpeg_in_a58 ;
assign	RG_quantized_block_59_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_59_en )
		RG_quantized_block_59 <= jpeg_in_a59 ;
always @ ( RG_k_quantized_block_03 or U_180 or jpeg_in_a60 or ST1_02d )
	RG_k_quantized_block_04_t = ( ( { 9{ ST1_02d } } & jpeg_in_a60 )	// line#=../rle.cpp:45
		| ( { 9{ U_180 } } & RG_k_quantized_block_03 ) ) ;
assign	RG_k_quantized_block_04_en = ( ST1_02d | U_180 ) ;
always @ ( posedge clk )
	if ( RG_k_quantized_block_04_en )
		RG_k_quantized_block_04 <= RG_k_quantized_block_04_t ;	// line#=../rle.cpp:45
always @ ( RG_k_02 or U_176 or jpeg_in_a61 or ST1_02d )
	RG_k_quantized_block_03_t = ( ( { 9{ ST1_02d } } & jpeg_in_a61 )	// line#=../rle.cpp:45
		| ( { 9{ U_176 } } & RG_k_02 [8:0] ) ) ;
assign	RG_k_quantized_block_03_en = ( ST1_02d | U_176 ) ;
always @ ( posedge clk )
	if ( RG_k_quantized_block_03_en )
		RG_k_quantized_block_03 <= RG_k_quantized_block_03_t ;	// line#=../rle.cpp:45
assign	RG_zz_02_en = U_173 ;
always @ ( posedge clk )
	if ( RG_zz_02_en )
		RG_zz_02 <= zz_RD2 ;
always @ ( zz_RD3 or U_88 or jpeg_in_a63 or ST1_02d )
	RG_previous_dc_quantized_block_t = ( ( { 9{ ST1_02d } } & jpeg_in_a63 )	// line#=../rle.cpp:45
		| ( { 9{ U_88 } } & zz_RD3 )					// line#=../rle.cpp:52,53
		) ;
assign	RG_previous_dc_quantized_block_en = ( ST1_02d | U_88 ) ;
always @ ( posedge clk )
	if ( RG_previous_dc_quantized_block_en )
		RG_previous_dc_quantized_block <= RG_previous_dc_quantized_block_t ;	// line#=../rle.cpp:45,52,53
always @ ( sub8u1ot or ST1_12d or incr8u1ot or ST1_09d or U_258 or incr8u2ot or 
	U_181 or ST1_02d )
	begin
	RG_len_05_t_c1 = ( U_258 | ST1_09d ) ;	// line#=../rle.cpp:79,80
	RG_len_05_t = ( ( { 8{ ST1_02d } } & 8'h01 )		// line#=../rle.cpp:39
		| ( { 8{ U_181 } } & incr8u2ot )		// line#=../rle.cpp:66,67,69,74
		| ( { 8{ RG_len_05_t_c1 } } & incr8u1ot )	// line#=../rle.cpp:79,80
		| ( { 8{ ST1_12d } } & sub8u1ot )		// line#=../rle.cpp:86
		) ;
	end
assign	RG_len_05_en = ( ST1_02d | U_181 | RG_len_05_t_c1 | ST1_12d ) ;
always @ ( posedge clk )
	if ( RG_len_05_en )
		RG_len_05 <= RG_len_05_t ;	// line#=../rle.cpp:39,66,67,69,74,79,80
						// ,86
always @ ( incr8u_61ot or ST1_03d )
	RG_k_t = ( { 6{ ST1_03d } } & incr8u_61ot )	// line#=../rle.cpp:111
		 ;	// line#=../rle.cpp:105
always @ ( posedge clk )
	RG_k <= RG_k_t ;	// line#=../rle.cpp:105,111
assign	M_129 = ( ST1_02d | U_06 ) ;
always @ ( CT_32 or ST1_07d or RG_i or U_173 or U_163 or U_79 or ST1_06d or U_161 or 
	U_81 or M_129 )
	begin
	FF_d_02_t_c1 = ( ( ( M_129 | U_81 ) | U_161 ) | ST1_06d ) ;	// line#=../rle.cpp:77,78,105,120,136,146
	FF_d_02_t_c2 = ( U_79 | U_163 ) ;	// line#=../rle.cpp:115,151
	FF_d_02_t = ( ( { 1{ FF_d_02_t_c2 } } & 1'h1 )				// line#=../rle.cpp:115,151
		| ( { 1{ U_173 } } & ( RG_i [31] | ( ~|RG_i [30:6] ) ) )	// line#=../rle.cpp:61,62
		| ( { 1{ ST1_07d } } & CT_32 )					// line#=../rle.cpp:77,78
		) ;	// line#=../rle.cpp:77,78,105,120,136,146
	end
assign	FF_d_02_en = ( FF_d_02_t_c1 | FF_d_02_t_c2 | U_173 | ST1_07d ) ;
always @ ( posedge clk )
	if ( FF_d_02_en )
		FF_d_02 <= FF_d_02_t ;	// line#=../rle.cpp:61,62,77,78,105,115
					// ,120,136,146,151
assign	FF_j_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:36
	if ( FF_j_en )
		FF_j <= 1'h0 ;
assign	RG_quantized_block_60_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_60_en )
		RG_quantized_block_60 <= jpeg_in_a62 ;
assign	RG_i_05_en = U_181 ;
always @ ( posedge clk )
	if ( RG_i_05_en )
		RG_i_05 <= RG_i_04 ;
assign	RG_i_04_en = U_180 ;
always @ ( posedge clk )
	if ( RG_i_04_en )
		RG_i_04 <= RG_i_03 ;
always @ ( CT_35 or ST1_11d or rl_rd00 or ST1_10d or FF_d_02 or ST1_08d or CT_32 or 
	ST1_06d or CT_31 or U_181 )
	RG_76_05_t = ( ( { 1{ U_181 } } & CT_31 )					// line#=../rle.cpp:66,67
		| ( { 1{ ST1_06d } } & CT_32 )						// line#=../rle.cpp:77,78
		| ( { 1{ ST1_08d } } & ( ~FF_d_02 ) )					// line#=../rle.cpp:77,78
		| ( { 1{ ST1_10d } } & ( ~|{ rl_rd00 [8:4] , ~rl_rd00 [3:0] } ) )	// line#=../rle.cpp:83,84
		| ( { 1{ ST1_11d } } & CT_35 )						// line#=../rle.cpp:83,84
		) ;
assign	RG_76_05_en = ( U_181 | ST1_06d | ST1_08d | ST1_10d | ST1_11d ) ;
always @ ( posedge clk )
	if ( RG_76_05_en )
		RG_76_05 <= RG_76_05_t ;	// line#=../rle.cpp:66,67,77,78,83,84
assign	RG_i_03_en = U_176 ;
always @ ( posedge clk )
	if ( RG_i_03_en )
		RG_i_03 <= RG_i_02 ;
assign	RG_i_02_en = U_173 ;
always @ ( posedge clk )
	if ( RG_i_02_en )
		RG_i_02 <= RG_i ;
assign	RG_k_02_en = U_173 ;
always @ ( posedge clk )	// line#=../rle.cpp:61,62
	if ( RG_k_02_en )
		RG_k_02 <= RG_j_k ;
always @ ( sub8u1ot or ST1_10d or incr8u1ot or M_134 or incr8u_71ot or ST1_04d or 
	RG_k or ST1_03d )
	RG_k_05_t = ( ( { 7{ ST1_03d } } & { 1'h0 , RG_k } )
		| ( { 7{ ST1_04d } } & incr8u_71ot )	// line#=../rle.cpp:142
		| ( { 7{ M_134 } } & incr8u1ot [6:0] )	// line#=../rle.cpp:68,69,73,74
		| ( { 7{ ST1_10d } } & sub8u1ot [6:0] )	// line#=../rle.cpp:83,84
		) ;
assign	RG_k_05_en = ( ST1_03d | ST1_04d | M_134 | ST1_10d ) ;
always @ ( posedge clk )
	if ( RG_k_05_en )
		RG_k_05 <= RG_k_05_t ;	// line#=../rle.cpp:68,69,73,74,83,84,142
assign	JF_01 = ~( ~|{ ~incr4s1ot [3] , incr4s1ot [2:0] } ) ;	// line#=../rle.cpp:34,35
assign	JF_03 = ~RG_k_05 [6] ;
assign	JF_03_port = JF_03 ;
assign	JF_07 = ~FF_d_02 ;	// line#=../rle.cpp:77,78
assign	JF_08 = ~CT_35 ;	// line#=../rle.cpp:83,84
assign	M_105 = ~|( FL01_01_streg ^ 2'h1 ) ;
assign	FL01_01_break = ( M_105 & FJ_05_11 ) ;
assign	FL01_02_break = ( ( U_206 | U_205 ) & FJ_07_08 ) ;
assign	FL01_03_break = ( FL01_03_streg & FJ_07_08 ) ;
always @ ( U_168 or U_237 )
	begin
	flag_r1_t_c1 = ( U_237 | U_168 ) ;
	flag_r1_t = ( { 1{ flag_r1_t_c1 } } & 1'h1 )
		 ;
	end
assign	flag_r1_en = ( flag_r1_t_c1 | U_198 ) ;
always @ ( posedge clk )
	if ( flag_r1_en )
		flag_r1 <= flag_r1_t ;
always @ ( U_168 or U_212 )
	begin
	flag_r2_t_c1 = ( U_212 | U_168 ) ;
	flag_r2_t = ( { 1{ flag_r2_t_c1 } } & 1'h1 )
		 ;
	end
assign	flag_r2_en = ( U_198 | flag_r2_t_c1 ) ;
always @ ( posedge clk )
	if ( flag_r2_en )
		flag_r2 <= flag_r2_t ;
always @ ( U_168 or U_225 )
	begin
	flag_r3_t_c1 = ( U_225 | U_168 ) ;
	flag_r3_t = ( { 1{ flag_r3_t_c1 } } & 1'h1 )
		 ;
	end
assign	flag_r3_en = ( flag_r3_t_c1 | U_208 ) ;
always @ ( posedge clk )
	if ( flag_r3_en )
		flag_r3 <= flag_r3_t ;
assign	FL01_01_01a = U_195 ;
assign	FL01_02_01a = U_206 ;
assign	FL01_03_01a = U_217 ;
assign	FL01_04_01a = U_225 ;
assign	FL01_05_01a = U_231 ;
assign	FL01_06_01a = U_237 ;
assign	FJ_05_11 = ( U_169 & ( ~C_07 ) ) ;	// line#=../rle.cpp:57,58
assign	FJ_07_08 = ( U_176 & ( ~( M_01_t1 & ( RG_k_02 [31] | ( ( ~|RG_k_02 [30:4] ) & ( 
	~&RG_k_02 [3:0] ) ) ) ) ) ) ;	// line#=../rle.cpp:61,62
assign	FL01_02_Leos = U_209 ;
assign	FL01_01_eos = ( M_135 | U_242 ) ;
assign	FL01_02_eos = ( U_209 | U_205 ) ;
assign	FL01_03_eos = ( M_136 | U_246 ) ;
assign	FL01_04_eos = M_137 ;
assign	FL01_05_eos = M_138 ;
assign	FL01_06_eos = M_139 ;
assign	M_128 = ( ( M_131 & ( ( ( U_190 & ( ~C_11 ) ) | ( U_198 & FL01_02_Lrdy ) ) | 
	( U_188 & FL01_02_Lrdy ) ) ) | U_168 ) ;
assign	M_131 = ( ST1_05d & ( ~FL01_01_break ) ) ;
assign	M_135 = ( ( ( ( U_195 & FJ_05_11 ) | ( U_200 & FL01_02_Lrdy ) ) | ( U_192 & 
	FL01_02_Lrdy ) ) | ( ST1_05d & ( ~|FL01_01_streg ) ) ) ;
always @ ( U_192 or FL01_02_Lrdy or U_200 or M_128 or M_135 or M_131 or U_242 )
	begin
	FL01_01_streg_t_c1 = ( ( U_242 | ( M_131 & M_135 ) ) | M_128 ) ;
	FL01_01_streg_t_c2 = ( M_131 & ( ( U_200 & ( ~FL01_02_Lrdy ) ) | ( U_192 & ( 
		~FL01_02_Lrdy ) ) ) ) ;
	FL01_01_streg_t = ( ( { 2{ FL01_01_streg_t_c1 } } & { 1'h0 , M_128 } )
		| ( { 2{ FL01_01_streg_t_c2 } } & 2'h2 ) ) ;
	end
assign	FL01_01_streg_en = ( FL01_01_streg_t_c1 | FL01_01_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_01_streg_en )
		FL01_01_streg <= FL01_01_streg_t ;
assign	M_127 = ( ST1_05d & FL01_02_break ) ;
always @ ( FL01_02_Leos_all or U_205 or U_215 or FL01_04_rdy or U_204 or U_208 or 
	U_206 )
	begin
	FL01_02_streg_t1_c1 = ( U_206 | U_208 ) ;
	FL01_02_streg_t1_c2 = ( ( U_204 & ( ~FL01_04_rdy ) ) | U_215 ) ;
	FL01_02_streg_t1_c3 = ( U_205 & ( ~FL01_02_Leos_all ) ) ;
	FL01_02_streg_t1 = ( ( { 2{ FL01_02_streg_t1_c1 } } & 2'h3 )
		| ( { 2{ FL01_02_streg_t1_c2 } } & 2'h1 )
		| ( { 2{ FL01_02_streg_t1_c3 } } & 2'h2 ) ) ;
	end
always @ ( FL01_02_streg_t1 or FL01_02_break or ST1_05d or U_168 or M_127 )
	begin
	FL01_02_streg_t_c1 = ( M_127 | U_168 ) ;
	FL01_02_streg_t_c2 = ( ST1_05d & ( ~FL01_02_break ) ) ;
	FL01_02_streg_t = ( ( { 2{ FL01_02_streg_t_c1 } } & { M_127 , 1'h0 } )
		| ( { 2{ FL01_02_streg_t_c2 } } & FL01_02_streg_t1 ) ) ;
	end
assign	FL01_02_streg_en = ( FL01_02_streg_t_c1 | FL01_02_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_02_streg_en )
		FL01_02_streg <= FL01_02_streg_t ;
assign	M_132 = ( ST1_05d & ( ~FL01_03_break ) ) ;
assign	M_136 = ( ( ( U_217 & FJ_07_08 ) | ( U_221 & ( ~FL01_02_ndat ) ) ) | ( U_216 & ( 
	~FL01_02_ndat ) ) ) ;
always @ ( U_216 or FL01_02_ndat or U_221 or M_136 or M_132 or U_168 or U_246 )
	begin
	FL01_03_streg_t_c1 = ( ( U_246 | U_168 ) | ( M_132 & M_136 ) ) ;
	FL01_03_streg_t_c2 = ( M_132 & ( ( U_221 & FL01_02_ndat ) | ( U_216 & FL01_02_ndat ) ) ) ;
	FL01_03_streg_t = ( { 1{ FL01_03_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_03_streg_en = ( FL01_03_streg_t_c1 | FL01_03_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_03_streg_en )
		FL01_03_streg <= FL01_03_streg_t ;
assign	M_137 = ( ( U_225 & ( ~FL01_02_Lndat ) ) | ( U_224 & ( ~FL01_02_Lndat ) ) ) ;
always @ ( FL01_02_Lndat or U_224 or U_228 or M_137 or ST1_05d or U_168 )
	begin
	FL01_04_streg_t_c1 = ( U_168 | ( ST1_05d & M_137 ) ) ;
	FL01_04_streg_t_c2 = ( ST1_05d & ( U_228 | ( U_224 & FL01_02_Lndat ) ) ) ;
	FL01_04_streg_t = ( { 1{ FL01_04_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_04_streg_en = ( FL01_04_streg_t_c1 | FL01_04_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_04_streg_en )
		FL01_04_streg <= FL01_04_streg_t ;
assign	M_138 = ( ( U_231 & ( ~FL01_04_ndat ) ) | ( U_230 & ( ~FL01_04_ndat ) ) ) ;
always @ ( U_230 or FL01_04_ndat or U_231 or M_138 or ST1_05d or U_168 )
	begin
	FL01_05_streg_t_c1 = ( U_168 | ( ST1_05d & M_138 ) ) ;
	FL01_05_streg_t_c2 = ( ST1_05d & ( ( U_231 & FL01_04_ndat ) | ( U_230 & FL01_04_ndat ) ) ) ;
	FL01_05_streg_t = ( { 1{ FL01_05_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_05_streg_en = ( FL01_05_streg_t_c1 | FL01_05_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_05_streg_en )
		FL01_05_streg <= FL01_05_streg_t ;
assign	M_139 = ( ( U_237 & ( ~FL01_05_ndat ) ) | ( U_236 & ( ~FL01_05_ndat ) ) ) ;
always @ ( U_236 or FL01_05_ndat or U_237 or M_139 or ST1_05d or U_168 )
	begin
	FL01_06_streg_t_c1 = ( U_168 | ( ST1_05d & M_139 ) ) ;
	FL01_06_streg_t_c2 = ( ST1_05d & ( ( U_237 & FL01_05_ndat ) | ( U_236 & FL01_05_ndat ) ) ) ;
	FL01_06_streg_t = ( { 1{ FL01_06_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_06_streg_en = ( FL01_06_streg_t_c1 | FL01_06_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_06_streg_en )
		FL01_06_streg <= FL01_06_streg_t ;
assign	FL01_01_ndat = ( U_198 | U_188 ) ;
assign	FL01_02_ndat = U_206 ;
assign	FL01_02_Lrdy = U_207 ;
assign	FL01_02_Lndat = ( U_204 | U_212 ) ;
assign	FL01_04_rdy = ( U_228 | U_224 ) ;
assign	FL01_04_ndat = U_225 ;
assign	FL01_05_ndat = U_231 ;
assign	jpeg_out_a00_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a00_r_en )
		jpeg_out_a00_r <= rl_rg00 ;
assign	jpeg_out_a01_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a01_r_en )
		jpeg_out_a01_r <= rl_rg01 ;
assign	jpeg_out_a02_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a02_r_en )
		jpeg_out_a02_r <= rl_rg02 ;
assign	jpeg_out_a03_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a03_r_en )
		jpeg_out_a03_r <= rl_rg03 ;
assign	jpeg_out_a04_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a04_r_en )
		jpeg_out_a04_r <= rl_rg04 ;
assign	jpeg_out_a05_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a05_r_en )
		jpeg_out_a05_r <= rl_rg05 ;
assign	jpeg_out_a06_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a06_r_en )
		jpeg_out_a06_r <= rl_rg06 ;
assign	jpeg_out_a07_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a07_r_en )
		jpeg_out_a07_r <= rl_rg07 ;
assign	jpeg_out_a08_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a08_r_en )
		jpeg_out_a08_r <= rl_rg08 ;
assign	jpeg_out_a09_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a09_r_en )
		jpeg_out_a09_r <= rl_rg09 ;
assign	jpeg_out_a10_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a10_r_en )
		jpeg_out_a10_r <= rl_rg10 ;
assign	jpeg_out_a11_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a11_r_en )
		jpeg_out_a11_r <= rl_rg11 ;
assign	jpeg_out_a12_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a12_r_en )
		jpeg_out_a12_r <= rl_rg12 ;
assign	jpeg_out_a13_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a13_r_en )
		jpeg_out_a13_r <= rl_rg13 ;
assign	jpeg_out_a14_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a14_r_en )
		jpeg_out_a14_r <= rl_rg14 ;
assign	jpeg_out_a15_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a15_r_en )
		jpeg_out_a15_r <= rl_rg15 ;
assign	jpeg_out_a16_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a16_r_en )
		jpeg_out_a16_r <= rl_rg16 ;
assign	jpeg_out_a17_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a17_r_en )
		jpeg_out_a17_r <= rl_rg17 ;
assign	jpeg_out_a18_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a18_r_en )
		jpeg_out_a18_r <= rl_rg18 ;
assign	jpeg_out_a19_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a19_r_en )
		jpeg_out_a19_r <= rl_rg19 ;
assign	jpeg_out_a20_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a20_r_en )
		jpeg_out_a20_r <= rl_rg20 ;
assign	jpeg_out_a21_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a21_r_en )
		jpeg_out_a21_r <= rl_rg21 ;
assign	jpeg_out_a22_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a22_r_en )
		jpeg_out_a22_r <= rl_rg22 ;
assign	jpeg_out_a23_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a23_r_en )
		jpeg_out_a23_r <= rl_rg23 ;
assign	jpeg_out_a24_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a24_r_en )
		jpeg_out_a24_r <= rl_rg24 ;
assign	jpeg_out_a25_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a25_r_en )
		jpeg_out_a25_r <= rl_rg25 ;
assign	jpeg_out_a26_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a26_r_en )
		jpeg_out_a26_r <= rl_rg26 ;
assign	jpeg_out_a27_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a27_r_en )
		jpeg_out_a27_r <= rl_rg27 ;
assign	jpeg_out_a28_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a28_r_en )
		jpeg_out_a28_r <= rl_rg28 ;
assign	jpeg_out_a29_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a29_r_en )
		jpeg_out_a29_r <= rl_rg29 ;
assign	jpeg_out_a30_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a30_r_en )
		jpeg_out_a30_r <= rl_rg30 ;
assign	jpeg_out_a31_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a31_r_en )
		jpeg_out_a31_r <= rl_rg31 ;
assign	jpeg_out_a32_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a32_r_en )
		jpeg_out_a32_r <= rl_rg32 ;
assign	jpeg_out_a33_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a33_r_en )
		jpeg_out_a33_r <= rl_rg33 ;
assign	jpeg_out_a34_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a34_r_en )
		jpeg_out_a34_r <= rl_rg34 ;
assign	jpeg_out_a35_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a35_r_en )
		jpeg_out_a35_r <= rl_rg35 ;
assign	jpeg_out_a36_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a36_r_en )
		jpeg_out_a36_r <= rl_rg36 ;
assign	jpeg_out_a37_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a37_r_en )
		jpeg_out_a37_r <= rl_rg37 ;
assign	jpeg_out_a38_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a38_r_en )
		jpeg_out_a38_r <= rl_rg38 ;
assign	jpeg_out_a39_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a39_r_en )
		jpeg_out_a39_r <= rl_rg39 ;
assign	jpeg_out_a40_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a40_r_en )
		jpeg_out_a40_r <= rl_rg40 ;
assign	jpeg_out_a41_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a41_r_en )
		jpeg_out_a41_r <= rl_rg41 ;
assign	jpeg_out_a42_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a42_r_en )
		jpeg_out_a42_r <= rl_rg42 ;
assign	jpeg_out_a43_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a43_r_en )
		jpeg_out_a43_r <= rl_rg43 ;
assign	jpeg_out_a44_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a44_r_en )
		jpeg_out_a44_r <= rl_rg44 ;
assign	jpeg_out_a45_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a45_r_en )
		jpeg_out_a45_r <= rl_rg45 ;
assign	jpeg_out_a46_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a46_r_en )
		jpeg_out_a46_r <= rl_rg46 ;
assign	jpeg_out_a47_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a47_r_en )
		jpeg_out_a47_r <= rl_rg47 ;
assign	jpeg_out_a48_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a48_r_en )
		jpeg_out_a48_r <= rl_rg48 ;
assign	jpeg_out_a49_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a49_r_en )
		jpeg_out_a49_r <= rl_rg49 ;
assign	jpeg_out_a50_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a50_r_en )
		jpeg_out_a50_r <= rl_rg50 ;
assign	jpeg_out_a51_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a51_r_en )
		jpeg_out_a51_r <= rl_rg51 ;
assign	jpeg_out_a52_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a52_r_en )
		jpeg_out_a52_r <= rl_rg52 ;
assign	jpeg_out_a53_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a53_r_en )
		jpeg_out_a53_r <= rl_rg53 ;
assign	jpeg_out_a54_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a54_r_en )
		jpeg_out_a54_r <= rl_rg54 ;
assign	jpeg_out_a55_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a55_r_en )
		jpeg_out_a55_r <= rl_rg55 ;
assign	jpeg_out_a56_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a56_r_en )
		jpeg_out_a56_r <= rl_rg56 ;
assign	jpeg_out_a57_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a57_r_en )
		jpeg_out_a57_r <= rl_rg57 ;
assign	jpeg_out_a58_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a58_r_en )
		jpeg_out_a58_r <= rl_rg58 ;
assign	jpeg_out_a59_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a59_r_en )
		jpeg_out_a59_r <= rl_rg59 ;
assign	jpeg_out_a60_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a60_r_en )
		jpeg_out_a60_r <= rl_rg60 ;
assign	jpeg_out_a61_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a61_r_en )
		jpeg_out_a61_r <= rl_rg61 ;
assign	jpeg_out_a62_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a62_r_en )
		jpeg_out_a62_r <= rl_rg62 ;
assign	jpeg_out_a63_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a63_r_en )
		jpeg_out_a63_r <= rl_rg63 ;
assign	jpeg_out_a64_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a64_r_en )
		jpeg_out_a64_r <= rl_rg64 ;
assign	jpeg_out_a65_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a65_r_en )
		jpeg_out_a65_r <= rl_rg65 ;
assign	jpeg_out_a66_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a66_r_en )
		jpeg_out_a66_r <= rl_rg66 ;
assign	jpeg_out_a67_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a67_r_en )
		jpeg_out_a67_r <= rl_rg67 ;
assign	jpeg_out_a68_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a68_r_en )
		jpeg_out_a68_r <= rl_rg68 ;
assign	jpeg_out_a69_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a69_r_en )
		jpeg_out_a69_r <= rl_rg69 ;
assign	jpeg_out_a70_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a70_r_en )
		jpeg_out_a70_r <= rl_rg70 ;
assign	jpeg_out_a71_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a71_r_en )
		jpeg_out_a71_r <= rl_rg71 ;
assign	jpeg_out_a72_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a72_r_en )
		jpeg_out_a72_r <= rl_rg72 ;
assign	jpeg_out_a73_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a73_r_en )
		jpeg_out_a73_r <= rl_rg73 ;
assign	jpeg_out_a74_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a74_r_en )
		jpeg_out_a74_r <= rl_rg74 ;
assign	jpeg_out_a75_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a75_r_en )
		jpeg_out_a75_r <= rl_rg75 ;
assign	jpeg_out_a76_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a76_r_en )
		jpeg_out_a76_r <= rl_rg76 ;
assign	jpeg_out_a77_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a77_r_en )
		jpeg_out_a77_r <= rl_rg77 ;
assign	jpeg_out_a78_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a78_r_en )
		jpeg_out_a78_r <= rl_rg78 ;
assign	jpeg_out_a79_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a79_r_en )
		jpeg_out_a79_r <= rl_rg79 ;
assign	jpeg_out_a80_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a80_r_en )
		jpeg_out_a80_r <= rl_rg80 ;
assign	jpeg_out_a81_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a81_r_en )
		jpeg_out_a81_r <= rl_rg81 ;
assign	jpeg_out_a82_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a82_r_en )
		jpeg_out_a82_r <= rl_rg82 ;
assign	jpeg_out_a83_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a83_r_en )
		jpeg_out_a83_r <= rl_rg83 ;
assign	jpeg_out_a84_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a84_r_en )
		jpeg_out_a84_r <= rl_rg84 ;
assign	jpeg_out_a85_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a85_r_en )
		jpeg_out_a85_r <= rl_rg85 ;
assign	jpeg_out_a86_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a86_r_en )
		jpeg_out_a86_r <= rl_rg86 ;
assign	jpeg_out_a87_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a87_r_en )
		jpeg_out_a87_r <= rl_rg87 ;
assign	jpeg_out_a88_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a88_r_en )
		jpeg_out_a88_r <= rl_rg88 ;
assign	jpeg_out_a89_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a89_r_en )
		jpeg_out_a89_r <= rl_rg89 ;
assign	jpeg_out_a90_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a90_r_en )
		jpeg_out_a90_r <= rl_rg90 ;
assign	jpeg_out_a91_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a91_r_en )
		jpeg_out_a91_r <= rl_rg91 ;
assign	jpeg_out_a92_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a92_r_en )
		jpeg_out_a92_r <= rl_rg92 ;
assign	jpeg_out_a93_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a93_r_en )
		jpeg_out_a93_r <= rl_rg93 ;
assign	jpeg_out_a94_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a94_r_en )
		jpeg_out_a94_r <= rl_rg94 ;
assign	jpeg_out_a95_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a95_r_en )
		jpeg_out_a95_r <= rl_rg95 ;
assign	jpeg_out_a96_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a96_r_en )
		jpeg_out_a96_r <= rl_rg96 ;
assign	jpeg_out_a97_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a97_r_en )
		jpeg_out_a97_r <= rl_rg97 ;
assign	jpeg_out_a98_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a98_r_en )
		jpeg_out_a98_r <= rl_rg98 ;
assign	jpeg_out_a99_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a99_r_en )
		jpeg_out_a99_r <= rl_rg99 ;
assign	jpeg_out_a100_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a100_r_en )
		jpeg_out_a100_r <= rl_rg100 ;
assign	jpeg_out_a101_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a101_r_en )
		jpeg_out_a101_r <= rl_rg101 ;
assign	jpeg_out_a102_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a102_r_en )
		jpeg_out_a102_r <= rl_rg102 ;
assign	jpeg_out_a103_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a103_r_en )
		jpeg_out_a103_r <= rl_rg103 ;
assign	jpeg_out_a104_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a104_r_en )
		jpeg_out_a104_r <= rl_rg104 ;
assign	jpeg_out_a105_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a105_r_en )
		jpeg_out_a105_r <= rl_rg105 ;
assign	jpeg_out_a106_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a106_r_en )
		jpeg_out_a106_r <= rl_rg106 ;
assign	jpeg_out_a107_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a107_r_en )
		jpeg_out_a107_r <= rl_rg107 ;
assign	jpeg_out_a108_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a108_r_en )
		jpeg_out_a108_r <= rl_rg108 ;
assign	jpeg_out_a109_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a109_r_en )
		jpeg_out_a109_r <= rl_rg109 ;
assign	jpeg_out_a110_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a110_r_en )
		jpeg_out_a110_r <= rl_rg110 ;
assign	jpeg_out_a111_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a111_r_en )
		jpeg_out_a111_r <= rl_rg111 ;
assign	jpeg_out_a112_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a112_r_en )
		jpeg_out_a112_r <= rl_rg112 ;
assign	jpeg_out_a113_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a113_r_en )
		jpeg_out_a113_r <= rl_rg113 ;
assign	jpeg_out_a114_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a114_r_en )
		jpeg_out_a114_r <= rl_rg114 ;
assign	jpeg_out_a115_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a115_r_en )
		jpeg_out_a115_r <= rl_rg115 ;
assign	jpeg_out_a116_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a116_r_en )
		jpeg_out_a116_r <= rl_rg116 ;
assign	jpeg_out_a117_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a117_r_en )
		jpeg_out_a117_r <= rl_rg117 ;
assign	jpeg_out_a118_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a118_r_en )
		jpeg_out_a118_r <= rl_rg118 ;
assign	jpeg_out_a119_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a119_r_en )
		jpeg_out_a119_r <= rl_rg119 ;
assign	jpeg_out_a120_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a120_r_en )
		jpeg_out_a120_r <= rl_rg120 ;
assign	jpeg_out_a121_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a121_r_en )
		jpeg_out_a121_r <= rl_rg121 ;
assign	jpeg_out_a122_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a122_r_en )
		jpeg_out_a122_r <= rl_rg122 ;
assign	jpeg_out_a123_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a123_r_en )
		jpeg_out_a123_r <= rl_rg123 ;
assign	jpeg_out_a124_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a124_r_en )
		jpeg_out_a124_r <= rl_rg124 ;
assign	jpeg_out_a125_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a125_r_en )
		jpeg_out_a125_r <= rl_rg125 ;
assign	jpeg_out_a126_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a126_r_en )
		jpeg_out_a126_r <= rl_rg126 ;
assign	jpeg_out_a127_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a127_r_en )
		jpeg_out_a127_r <= rl_rg127 ;
assign	jpeg_len_out_r_en = U_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:93
	if ( jpeg_len_out_r_en )
		jpeg_len_out_r <= { 4'h0 , RG_len_05 } ;
always @ ( U_263 )
	valid_r_t = ( { 1{ U_263 } } & 1'h1 )	// line#=../rle.cpp:95
		 ;	// line#=../rle.cpp:30
assign	valid_r_en = ( ST1_01d | U_263 ) ;
always @ ( posedge clk )
	if ( valid_r_en )
		valid_r <= valid_r_t ;	// line#=../rle.cpp:30,95
assign	sub8u1i1 = { ( ST1_12d & RG_len_05 [7] ) , RG_len_05 [6:0] } ;	// line#=../rle.cpp:77,78,83,84,86
always @ ( U_264 or ST1_10d or ST1_12d or ST1_07d )
	begin
	sub8u1i2_c1 = ( ST1_07d | ST1_12d ) ;	// line#=../rle.cpp:77,78,86
	sub8u1i2 = ( ( { 3{ sub8u1i2_c1 } } & 3'h2 )	// line#=../rle.cpp:77,78,86
		| ( { 3{ ST1_10d } } & 3'h4 )		// line#=../rle.cpp:83,84
		| ( { 3{ U_264 } } & 3'h3 )		// line#=../rle.cpp:83,84
		) ;
	end
assign	incr8u1i1 = RG_len_05 ;	// line#=../rle.cpp:68,73,79,80
assign	incr8u2i1 = incr8u1ot ;	// line#=../rle.cpp:68,69,73,74
assign	incr32s1i1 = RG_j_k ;	// line#=../rle.cpp:61,62,64,114,125,145
				// ,156
assign	incr32s2i1 = RG_i ;	// line#=../rle.cpp:61,62,63,119,129,150
				// ,160
assign	decr32s1i1 = RG_i ;	// line#=../rle.cpp:124,155
assign	decr32s2i1 = RG_j_k ;	// line#=../rle.cpp:130,161
always @ ( RG_i_05 or U_187 or RG_k_05 or U_89 or U_90 or U_91 or U_92 or U_93 or 
	U_94 or U_95 or U_96 or RG_k or U_07 or U_08 or U_09 or U_10 or U_11 or 
	U_12 or U_13 or U_14 )
	begin
	zz_AD1_c1 = ( ( ( ( ( ( ( U_14 | U_13 ) | U_12 ) | U_11 ) | U_10 ) | U_09 ) | 
		U_08 ) | U_07 ) ;	// line#=../rle.cpp:111
	zz_AD1_c2 = ( ( ( ( ( ( ( U_96 | U_95 ) | U_94 ) | U_93 ) | U_92 ) | U_91 ) | 
		U_90 ) | U_89 ) ;	// line#=../rle.cpp:142
	zz_AD1 = ( ( { 6{ zz_AD1_c1 } } & RG_k )		// line#=../rle.cpp:111
		| ( { 6{ zz_AD1_c2 } } & RG_k_05 [5:0] )	// line#=../rle.cpp:142
		| ( { 6{ U_187 } } & RG_i_05 [5:0] )		// line#=../rle.cpp:74
		) ;
	end
always @ ( RG_quantized_block_7 or RG_quantized_block_6 or RG_quantized_block_5 or 
	RG_quantized_block_4 or RG_quantized_block_3 or RG_quantized_block_2 or 
	RG_quantized_block_1 or RG_quantized_block or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_06 = RG_quantized_block ;	// line#=../rle.cpp:111
	3'h1 :
		TR_06 = RG_quantized_block_1 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_06 = RG_quantized_block_2 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_06 = RG_quantized_block_3 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_06 = RG_quantized_block_4 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_06 = RG_quantized_block_5 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_06 = RG_quantized_block_6 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_06 = RG_quantized_block_7 ;	// line#=../rle.cpp:111
	default :
		TR_06 = 9'hx ;
	endcase
always @ ( RG_quantized_block_15 or RG_quantized_block_14 or RG_quantized_block_13 or 
	RG_quantized_block_12 or RG_quantized_block_11 or RG_quantized_block_10 or 
	RG_quantized_block_9 or RG_quantized_block_8 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_07 = RG_quantized_block_8 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_07 = RG_quantized_block_9 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_07 = RG_quantized_block_10 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_07 = RG_quantized_block_11 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_07 = RG_quantized_block_12 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_07 = RG_quantized_block_13 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_07 = RG_quantized_block_14 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_07 = RG_quantized_block_15 ;	// line#=../rle.cpp:111
	default :
		TR_07 = 9'hx ;
	endcase
always @ ( RG_quantized_block_23 or RG_quantized_block_22 or RG_quantized_block_21 or 
	RG_quantized_block_20 or RG_quantized_block_19 or RG_quantized_block_18 or 
	RG_quantized_block_17 or RG_quantized_block_16 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_08 = RG_quantized_block_16 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_08 = RG_quantized_block_17 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_08 = RG_quantized_block_18 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_08 = RG_quantized_block_19 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_08 = RG_quantized_block_20 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_08 = RG_quantized_block_21 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_08 = RG_quantized_block_22 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_08 = RG_quantized_block_23 ;	// line#=../rle.cpp:111
	default :
		TR_08 = 9'hx ;
	endcase
always @ ( RG_quantized_block_31 or RG_quantized_block_30 or RG_quantized_block_29 or 
	RG_quantized_block_28 or RG_quantized_block_27 or RG_quantized_block_26 or 
	RG_quantized_block_25 or RG_quantized_block_24 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_09 = RG_quantized_block_24 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_09 = RG_quantized_block_25 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_09 = RG_quantized_block_26 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_09 = RG_quantized_block_27 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_09 = RG_quantized_block_28 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_09 = RG_quantized_block_29 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_09 = RG_quantized_block_30 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_09 = RG_quantized_block_31 ;	// line#=../rle.cpp:111
	default :
		TR_09 = 9'hx ;
	endcase
always @ ( RG_quantized_block_39 or RG_quantized_block_38 or RG_quantized_block_37 or 
	RG_quantized_block_36 or RG_quantized_block_35 or RG_quantized_block_34 or 
	RG_quantized_block_33 or RG_quantized_block_32 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_10 = RG_quantized_block_32 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_10 = RG_quantized_block_33 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_10 = RG_quantized_block_34 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_10 = RG_quantized_block_35 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_10 = RG_quantized_block_36 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_10 = RG_quantized_block_37 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_10 = RG_quantized_block_38 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_10 = RG_quantized_block_39 ;	// line#=../rle.cpp:111
	default :
		TR_10 = 9'hx ;
	endcase
always @ ( RG_quantized_block_47 or RG_quantized_block_46 or RG_quantized_block_45 or 
	RG_quantized_block_44 or RG_quantized_block_43 or RG_quantized_block_42 or 
	RG_quantized_block_41 or RG_quantized_block_40 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_11 = RG_quantized_block_40 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_11 = RG_quantized_block_41 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_11 = RG_quantized_block_42 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_11 = RG_quantized_block_43 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_11 = RG_quantized_block_44 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_11 = RG_quantized_block_45 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_11 = RG_quantized_block_46 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_11 = RG_quantized_block_47 ;	// line#=../rle.cpp:111
	default :
		TR_11 = 9'hx ;
	endcase
always @ ( RG_quantized_block_55 or RG_quantized_block_54 or RG_quantized_block_53 or 
	RG_quantized_block_52 or RG_quantized_block_51 or RG_quantized_block_50 or 
	RG_quantized_block_49 or RG_quantized_block_48 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_12 = RG_quantized_block_48 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_12 = RG_quantized_block_49 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_12 = RG_quantized_block_50 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_12 = RG_quantized_block_51 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_12 = RG_quantized_block_52 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_12 = RG_quantized_block_53 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_12 = RG_quantized_block_54 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_12 = RG_quantized_block_55 ;	// line#=../rle.cpp:111
	default :
		TR_12 = 9'hx ;
	endcase
always @ ( RG_previous_dc_quantized_block or RG_quantized_block_60 or RG_k_quantized_block_03 or 
	RG_k_quantized_block_04 or RG_quantized_block_59 or RG_quantized_block_58 or 
	RG_quantized_block_57 or RG_quantized_block_56 or RG_j_k )	// line#=../rle.cpp:111
	case ( RG_j_k [2:0] )
	3'h0 :
		TR_13 = RG_quantized_block_56 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_13 = RG_quantized_block_57 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_13 = RG_quantized_block_58 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_13 = RG_quantized_block_59 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_13 = RG_k_quantized_block_04 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_13 = RG_k_quantized_block_03 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_13 = RG_quantized_block_60 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_13 = RG_previous_dc_quantized_block ;	// line#=../rle.cpp:111
	default :
		TR_13 = 9'hx ;
	endcase
always @ ( U_96 or U_95 or U_94 or U_93 or U_92 or U_91 or U_90 or U_89 or TR_13 or 
	U_14 or TR_12 or U_13 or TR_11 or U_12 or TR_10 or U_11 or TR_09 or U_10 or 
	TR_08 or U_09 or TR_07 or U_08 or TR_06 or U_07 )
	zz_WD1 = ( ( { 9{ U_07 } } & TR_06 )	// line#=../rle.cpp:111
		| ( { 9{ U_08 } } & TR_07 )	// line#=../rle.cpp:111
		| ( { 9{ U_09 } } & TR_08 )	// line#=../rle.cpp:111
		| ( { 9{ U_10 } } & TR_09 )	// line#=../rle.cpp:111
		| ( { 9{ U_11 } } & TR_10 )	// line#=../rle.cpp:111
		| ( { 9{ U_12 } } & TR_11 )	// line#=../rle.cpp:111
		| ( { 9{ U_13 } } & TR_12 )	// line#=../rle.cpp:111
		| ( { 9{ U_14 } } & TR_13 )	// line#=../rle.cpp:111
		| ( { 9{ U_89 } } & TR_06 )	// line#=../rle.cpp:142
		| ( { 9{ U_90 } } & TR_07 )	// line#=../rle.cpp:142
		| ( { 9{ U_91 } } & TR_08 )	// line#=../rle.cpp:142
		| ( { 9{ U_92 } } & TR_09 )	// line#=../rle.cpp:142
		| ( { 9{ U_93 } } & TR_10 )	// line#=../rle.cpp:142
		| ( { 9{ U_94 } } & TR_11 )	// line#=../rle.cpp:142
		| ( { 9{ U_95 } } & TR_12 )	// line#=../rle.cpp:142
		| ( { 9{ U_96 } } & TR_13 )	// line#=../rle.cpp:142
		) ;
assign	M_104 = ~|( RG_j_k [2:0] ^ 3'h1 ) ;	// line#=../rle.cpp:111,142
assign	M_108 = ~|RG_j_k [2:0] ;	// line#=../rle.cpp:111,142
assign	M_113 = ~|( RG_j_k [2:0] ^ 3'h2 ) ;	// line#=../rle.cpp:111,142
assign	M_116 = ~|( RG_j_k [2:0] ^ 3'h7 ) ;	// line#=../rle.cpp:111,142
assign	M_118 = ~|( RG_j_k [2:0] ^ 3'h4 ) ;	// line#=../rle.cpp:111,142
assign	M_120 = ~|( RG_j_k [2:0] ^ 3'h3 ) ;	// line#=../rle.cpp:111,142
assign	M_123 = ~|( RG_j_k [2:0] ^ 3'h5 ) ;	// line#=../rle.cpp:111,142
assign	M_125 = ~|( RG_j_k [2:0] ^ 3'h6 ) ;	// line#=../rle.cpp:111,142
assign	zz_WE1 = ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( U_14 & M_116 ) | ( U_14 & M_125 ) ) | 
	( U_14 & M_123 ) ) | ( U_14 & M_118 ) ) | ( U_14 & M_120 ) ) | ( U_14 & M_113 ) ) | 
	( U_14 & M_104 ) ) | ( U_14 & M_108 ) ) | ( U_13 & M_116 ) ) | ( U_13 & M_125 ) ) | 
	( U_13 & M_123 ) ) | ( U_13 & M_118 ) ) | ( U_13 & M_120 ) ) | ( U_13 & M_113 ) ) | 
	( U_13 & M_104 ) ) | ( U_13 & M_108 ) ) | ( U_12 & M_116 ) ) | ( U_12 & M_125 ) ) | 
	( U_12 & M_123 ) ) | ( U_12 & M_118 ) ) | ( U_12 & M_120 ) ) | ( U_12 & M_113 ) ) | 
	( U_12 & M_104 ) ) | ( U_12 & M_108 ) ) | ( U_11 & M_116 ) ) | ( U_11 & M_125 ) ) | 
	( U_11 & M_123 ) ) | ( U_11 & M_118 ) ) | ( U_11 & M_120 ) ) | ( U_11 & M_113 ) ) | 
	( U_11 & M_104 ) ) | ( U_11 & M_108 ) ) | ( U_10 & M_116 ) ) | ( U_10 & M_125 ) ) | 
	( U_10 & M_123 ) ) | ( U_10 & M_118 ) ) | ( U_10 & M_120 ) ) | ( U_10 & M_113 ) ) | 
	( U_10 & M_104 ) ) | ( U_10 & M_108 ) ) | ( U_09 & M_116 ) ) | ( U_09 & M_125 ) ) | 
	( U_09 & M_123 ) ) | ( U_09 & M_118 ) ) | ( U_09 & M_120 ) ) | ( U_09 & M_113 ) ) | 
	( U_09 & M_104 ) ) | ( U_09 & M_108 ) ) | ( U_08 & M_116 ) ) | ( U_08 & M_125 ) ) | 
	( U_08 & M_123 ) ) | ( U_08 & M_118 ) ) | ( U_08 & M_120 ) ) | ( U_08 & M_113 ) ) | 
	( U_08 & M_104 ) ) | ( U_08 & M_108 ) ) | ( U_07 & M_116 ) ) | ( U_07 & M_125 ) ) | 
	( U_07 & M_123 ) ) | ( U_07 & M_118 ) ) | ( U_07 & M_120 ) ) | ( U_07 & M_113 ) ) | 
	( U_07 & M_104 ) ) | ( U_07 & M_108 ) ) | ( U_96 & M_116 ) ) | ( U_96 & M_125 ) ) | 
	( U_96 & M_123 ) ) | ( U_96 & M_118 ) ) | ( U_96 & M_120 ) ) | ( U_96 & M_113 ) ) | 
	( U_96 & M_104 ) ) | ( U_96 & M_108 ) ) | ( U_95 & M_116 ) ) | ( U_95 & M_125 ) ) | 
	( U_95 & M_123 ) ) | ( U_95 & M_118 ) ) | ( U_95 & M_120 ) ) | ( U_95 & M_113 ) ) | 
	( U_95 & M_104 ) ) | ( U_95 & M_108 ) ) | ( U_94 & M_116 ) ) | ( U_94 & M_125 ) ) | 
	( U_94 & M_123 ) ) | ( U_94 & M_118 ) ) | ( U_94 & M_120 ) ) | ( U_94 & M_113 ) ) | 
	( U_94 & M_104 ) ) | ( U_94 & M_108 ) ) | ( U_93 & M_116 ) ) | ( U_93 & M_125 ) ) | 
	( U_93 & M_123 ) ) | ( U_93 & M_118 ) ) | ( U_93 & M_120 ) ) | ( U_93 & M_113 ) ) | 
	( U_93 & M_104 ) ) | ( U_93 & M_108 ) ) | ( U_92 & M_116 ) ) | ( U_92 & M_125 ) ) | 
	( U_92 & M_123 ) ) | ( U_92 & M_118 ) ) | ( U_92 & M_120 ) ) | ( U_92 & M_113 ) ) | 
	( U_92 & M_104 ) ) | ( U_92 & M_108 ) ) | ( U_91 & M_116 ) ) | ( U_91 & M_125 ) ) | 
	( U_91 & M_123 ) ) | ( U_91 & M_118 ) ) | ( U_91 & M_120 ) ) | ( U_91 & M_113 ) ) | 
	( U_91 & M_104 ) ) | ( U_91 & M_108 ) ) | ( U_90 & M_116 ) ) | ( U_90 & M_125 ) ) | 
	( U_90 & M_123 ) ) | ( U_90 & M_118 ) ) | ( U_90 & M_120 ) ) | ( U_90 & M_113 ) ) | 
	( U_90 & M_104 ) ) | ( U_90 & M_108 ) ) | ( U_89 & M_116 ) ) | ( U_89 & M_125 ) ) | 
	( U_89 & M_123 ) ) | ( U_89 & M_118 ) ) | ( U_89 & M_120 ) ) | ( U_89 & M_113 ) ) | 
	( U_89 & M_104 ) ) | ( U_89 & M_108 ) ) ;
always @ ( sub8u1ot or ST1_10d or U_264 or ST1_07d or decr8u_71ot or ST1_06d )
	begin
	rl_ad00_c1 = ( ( ST1_07d | U_264 ) | ST1_10d ) ;	// line#=../rle.cpp:77,78,83,84
	rl_ad00 = ( ( { 7{ ST1_06d } } & decr8u_71ot )		// line#=../rle.cpp:77,78
		| ( { 7{ rl_ad00_c1 } } & sub8u1ot [6:0] )	// line#=../rle.cpp:77,78,83,84
		) ;
	end
assign	rl_ad01 = RG_k_05 ;	// line#=../rle.cpp:69,85
assign	rl_ad02 = RG_len_05 [6:0] ;	// line#=../rle.cpp:68,73,79,80
always @ ( RG_k_quantized_block_04 or U_183 )
	rl_wd02 = ( { 9{ U_183 } } & RG_k_quantized_block_04 )	// line#=../rle.cpp:73
		 ;	// line#=../rle.cpp:68,79,80
assign	rl_we01 = ( U_186 | ST1_12d ) ;	// line#=../rle.cpp:69,85
assign	M_134 = U_181 ;
assign	rl_we02 = ( ( M_134 | U_258 ) | ST1_09d ) ;	// line#=../rle.cpp:68,73,79,80

endmodule

module jpeg_incr8u_6 ( i1 ,o1 );
input	[5:0]	i1 ;
output	[5:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr8u_7 ( i1 ,o1 );
input	[5:0]	i1 ;
output	[6:0]	o1 ;

assign	o1 = ( { 1'h0 , i1 } + 1'h1 ) ;

endmodule

module jpeg_decr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_decr8u_7 ( i1 ,o1 );
input	[6:0]	i1 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_incr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr8u ( i1 ,o1 );
input	[7:0]	i1 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr4s ( i1 ,o1 );
input	[3:0]	i1 ;
output	[3:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_lop8u_1 ( i1 ,i2 ,o1 );
input	[5:0]	i1 ;
input	[5:0]	i2 ;
output		o1 ;
wire		M_01 ;

assign	M_01 = ( i1 < i2 ) ;
assign	o1 = M_01 ;

endmodule

module jpeg_sub12s_9 ( i1 ,i2 ,o1 );
input	[8:0]	i1 ;
input	[8:0]	i2 ;
output	[8:0]	o1 ;

assign	o1 = ( i1 - i2 ) ;

endmodule

module jpeg_sub8u ( i1 ,i2 ,o1 );
input	[7:0]	i1 ;
input	[2:0]	i2 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 - { 5'h00 , i2 } ) ;

endmodule

module jpeg_decoder_7to128 ( DECODER_in ,DECODER_out );
input	[6:0]	DECODER_in ;
output	[127:0]	DECODER_out ;
reg	[127:0]	DECODER_out ;

always @ ( DECODER_in )
	begin
	DECODER_out = 128'h00000000000000000000000000000000 ;
	DECODER_out [127 - DECODER_in] = 1'h1 ;
	end

endmodule

module jpeg_MEM_zz ( AD1 ,RD1 ,WD1 ,WE1 ,CLK1 ,RA2 ,RD2 ,RA3 ,RD3 );
input	[5:0]	AD1 ;
output	[8:0]	RD1 ;
input	[8:0]	WD1 ;
input		WE1 ;
input		CLK1 ;
input	[5:0]	RA2 ;
output	[8:0]	RD2 ;
input	[5:0]	RA3 ;
output	[8:0]	RD3 ;

jpeg_MEM_zz_subD INST_MEM_zz_subD_1 ( .RD1(RD1) ,.AD1(AD1) ,.WE1(WE1) ,.WD1(WD1) ,
	.CLK1(CLK1) ,.RD2(RD2) ,.RA2(RA2) );
jpeg_MEM_zz_subD INST_MEM_zz_subD_2 ( .RD1() ,.AD1(AD1) ,.WE1(WE1) ,.WD1(WD1) ,.CLK1(CLK1) ,
	.RD2(RD3) ,.RA2(RA3) );

endmodule

(* ram_extract = "yes" *)
module jpeg_MEM_zz_subD ( RD1 ,AD1 ,WE1 ,WD1 ,CLK1 ,RD2 ,RA2 );
output	[8:0]	RD1 ;
input	[5:0]	AD1 ;
input		WE1 ;
input	[8:0]	WD1 ;
input		CLK1 ;
output	[8:0]	RD2 ;
input	[5:0]	RA2 ;
(* ram_style = "distributed" *)reg	[8:0]	zz_r	[0:63] ;

assign	RD1 = zz_r[AD1] ;
assign	RD2 = zz_r[RA2] ;

always @ ( posedge CLK1 )
	begin
	if ( WE1 )
		zz_r [AD1] = WD1 ;
	end

endmodule
