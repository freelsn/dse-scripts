// verilog_out version 6.79.2
// options:  veriloggen jpeg_E.IFF
// bdlpars options:  -DDSE ../rle.cpp
// bdltran options:  -c1000 -s -Zresource_fcnt=GENERATE -Zresource_mcnt=GENERATE -lb /home/shuangnan/share/packages/zynq-1.BLIB -lfl /home/shuangnan/share/packages/zynq-1.FLIB jpeg.IFF -OX -a8196 -Zfu_cnt_incr_rate=0 -tcio 
// timestamp_0: 20180213181726_16339_92815
// timestamp_5: 20180213181731_17757_19297
// timestamp_9: 20180213181737_17757_90759
// timestamp_C: 20180213181737_17757_86776
// timestamp_E: 20180213181738_17757_06042
// timestamp_V: 20180213181742_20243_23258

module jpeg ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,jpeg_in_a04 ,
	jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,jpeg_in_a10 ,
	jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,jpeg_in_a16 ,
	jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,jpeg_in_a22 ,
	jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,jpeg_in_a28 ,
	jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,jpeg_in_a34 ,
	jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,jpeg_in_a40 ,
	jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,jpeg_in_a46 ,
	jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,jpeg_in_a52 ,
	jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,jpeg_in_a58 ,
	jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,jpeg_in_a64 ,
	jpeg_in_a65 ,jpeg_in_a66 ,jpeg_in_a67 ,jpeg_in_a68 ,jpeg_in_a69 ,jpeg_in_a70 ,
	jpeg_in_a71 ,jpeg_in_a72 ,jpeg_in_a73 ,jpeg_in_a74 ,jpeg_in_a75 ,jpeg_in_a76 ,
	jpeg_in_a77 ,jpeg_in_a78 ,jpeg_in_a79 ,jpeg_in_a80 ,jpeg_in_a81 ,jpeg_in_a82 ,
	jpeg_in_a83 ,jpeg_in_a84 ,jpeg_in_a85 ,jpeg_in_a86 ,jpeg_in_a87 ,jpeg_in_a88 ,
	jpeg_in_a89 ,jpeg_in_a90 ,jpeg_in_a91 ,jpeg_in_a92 ,jpeg_in_a93 ,jpeg_in_a94 ,
	jpeg_in_a95 ,jpeg_in_a96 ,jpeg_in_a97 ,jpeg_in_a98 ,jpeg_in_a99 ,jpeg_in_a100 ,
	jpeg_in_a101 ,jpeg_in_a102 ,jpeg_in_a103 ,jpeg_in_a104 ,jpeg_in_a105 ,jpeg_in_a106 ,
	jpeg_in_a107 ,jpeg_in_a108 ,jpeg_in_a109 ,jpeg_in_a110 ,jpeg_in_a111 ,jpeg_in_a112 ,
	jpeg_in_a113 ,jpeg_in_a114 ,jpeg_in_a115 ,jpeg_in_a116 ,jpeg_in_a117 ,jpeg_in_a118 ,
	jpeg_in_a119 ,jpeg_in_a120 ,jpeg_in_a121 ,jpeg_in_a122 ,jpeg_in_a123 ,jpeg_in_a124 ,
	jpeg_in_a125 ,jpeg_in_a126 ,jpeg_in_a127 ,jpeg_len_in ,jpeg_out_a00 ,jpeg_out_a01 ,
	jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,jpeg_out_a06 ,jpeg_out_a07 ,
	jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,jpeg_out_a12 ,jpeg_out_a13 ,
	jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,jpeg_out_a18 ,jpeg_out_a19 ,
	jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,jpeg_out_a24 ,jpeg_out_a25 ,
	jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,jpeg_out_a30 ,jpeg_out_a31 ,
	jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,jpeg_out_a36 ,jpeg_out_a37 ,
	jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,jpeg_out_a42 ,jpeg_out_a43 ,
	jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,jpeg_out_a48 ,jpeg_out_a49 ,
	jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,jpeg_out_a54 ,jpeg_out_a55 ,
	jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,jpeg_out_a60 ,jpeg_out_a61 ,
	jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,jpeg_out_a66 ,jpeg_out_a67 ,
	jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,jpeg_out_a72 ,jpeg_out_a73 ,
	jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,jpeg_out_a78 ,jpeg_out_a79 ,
	jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,jpeg_out_a84 ,jpeg_out_a85 ,
	jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,jpeg_out_a90 ,jpeg_out_a91 ,
	jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,jpeg_out_a96 ,jpeg_out_a97 ,
	jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,jpeg_out_a102 ,
	jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,jpeg_out_a107 ,
	jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,jpeg_out_a112 ,
	jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,jpeg_out_a117 ,
	jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,jpeg_out_a122 ,
	jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,jpeg_out_a127 ,
	jpeg_len_out ,valid );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a64 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a65 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a66 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a67 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a68 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a69 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a70 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a71 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a72 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a73 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a74 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a75 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a76 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a77 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a78 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a79 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a80 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a81 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a82 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a83 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a84 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a85 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a86 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a87 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a88 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a89 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a90 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a91 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a92 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a93 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a94 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a95 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a96 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a97 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a98 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a99 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a100 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a101 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a102 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a103 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a104 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a105 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a106 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a107 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a108 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a109 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a110 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a111 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a112 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a113 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a114 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a115 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a116 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a117 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a118 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a119 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a120 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a121 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a122 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a123 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a124 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a125 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a126 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a127 ;	// line#=../rle.h:56
input	[11:0]	jpeg_len_in ;	// line#=../rle.h:57
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
wire		ST1_01d ;
wire		ST1_02d ;
wire		ST1_03d ;
wire		ST1_04d ;
wire		ST1_05d ;
wire		ST1_06d ;
wire		ST1_07d ;
wire		ST1_08d ;
wire		ST1_09d ;
wire		ST1_10d ;
wire		ST1_11d ;
wire		ST1_12d ;
wire		ST1_13d ;
wire		ST1_14d ;
wire		ST1_15d ;
wire		ST1_16d ;
wire		ST1_17d ;
wire		ST1_18d ;
wire		ST1_19d ;
wire		ST1_20d ;
wire		ST1_21d ;
wire		ST1_22d ;
wire		ST1_23d ;
wire		ST1_24d ;
wire		ST1_25d ;
wire		ST1_26d ;
wire		ST1_27d ;
wire		ST1_28d ;
wire		ST1_29d ;
wire		ST1_30d ;
wire		ST1_31d ;
wire		ST1_32d ;
wire		ST1_33d ;
wire		ST1_34d ;
wire		ST1_35d ;
wire		ST1_36d ;
wire		ST1_37d ;
wire		ST1_38d ;
wire		ST1_39d ;
wire		ST1_40d ;
wire		ST1_41d ;
wire		ST1_42d ;
wire		ST1_43d ;
wire		ST1_44d ;
wire		ST1_45d ;
wire		ST1_46d ;
wire		ST1_47d ;
wire		ST1_48d ;
wire		ST1_49d ;
wire		ST1_50d ;
wire		ST1_51d ;
wire		ST1_52d ;
wire		ST1_53d ;
wire		ST1_54d ;
wire		ST1_55d ;
wire		ST1_56d ;
wire		JF_01 ;
wire		lop8u_11ot ;
wire		JF_03 ;
wire		CT_31 ;
wire		JF_05 ;
wire		FL01_01_Leos_all ;
wire		FL02_01_Leos_all ;

jpeg_fsm INST_fsm ( .clk(clk) ,.rst(rst) ,.ST1_56d(ST1_56d) ,.ST1_55d(ST1_55d) ,
	.ST1_54d(ST1_54d) ,.ST1_53d(ST1_53d) ,.ST1_52d(ST1_52d) ,.ST1_51d(ST1_51d) ,
	.ST1_50d(ST1_50d) ,.ST1_49d(ST1_49d) ,.ST1_48d(ST1_48d) ,.ST1_47d(ST1_47d) ,
	.ST1_46d(ST1_46d) ,.ST1_45d(ST1_45d) ,.ST1_44d(ST1_44d) ,.ST1_43d(ST1_43d) ,
	.ST1_42d(ST1_42d) ,.ST1_41d(ST1_41d) ,.ST1_40d(ST1_40d) ,.ST1_39d(ST1_39d) ,
	.ST1_38d(ST1_38d) ,.ST1_37d(ST1_37d) ,.ST1_36d(ST1_36d) ,.ST1_35d(ST1_35d) ,
	.ST1_34d(ST1_34d) ,.ST1_33d(ST1_33d) ,.ST1_32d(ST1_32d) ,.ST1_31d(ST1_31d) ,
	.ST1_30d(ST1_30d) ,.ST1_29d(ST1_29d) ,.ST1_28d(ST1_28d) ,.ST1_27d(ST1_27d) ,
	.ST1_26d(ST1_26d) ,.ST1_25d(ST1_25d) ,.ST1_24d(ST1_24d) ,.ST1_23d(ST1_23d) ,
	.ST1_22d(ST1_22d) ,.ST1_21d(ST1_21d) ,.ST1_20d(ST1_20d) ,.ST1_19d(ST1_19d) ,
	.ST1_18d(ST1_18d) ,.ST1_17d(ST1_17d) ,.ST1_16d(ST1_16d) ,.ST1_15d(ST1_15d) ,
	.ST1_14d(ST1_14d) ,.ST1_13d(ST1_13d) ,.ST1_12d(ST1_12d) ,.ST1_11d(ST1_11d) ,
	.ST1_10d(ST1_10d) ,.ST1_09d(ST1_09d) ,.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,
	.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,
	.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,.JF_01(JF_01) ,.lop8u_11ot(lop8u_11ot) ,
	.JF_03(JF_03) ,.CT_31(CT_31) ,.JF_05(JF_05) ,.FL01_01_Leos_all(FL01_01_Leos_all) ,
	.FL02_01_Leos_all(FL02_01_Leos_all) );
jpeg_dat INST_dat ( .clk(clk) ,.rst(rst) ,.jpeg_in_a00(jpeg_in_a00) ,.jpeg_in_a01(jpeg_in_a01) ,
	.jpeg_in_a02(jpeg_in_a02) ,.jpeg_in_a03(jpeg_in_a03) ,.jpeg_in_a04(jpeg_in_a04) ,
	.jpeg_in_a05(jpeg_in_a05) ,.jpeg_in_a06(jpeg_in_a06) ,.jpeg_in_a07(jpeg_in_a07) ,
	.jpeg_in_a08(jpeg_in_a08) ,.jpeg_in_a09(jpeg_in_a09) ,.jpeg_in_a10(jpeg_in_a10) ,
	.jpeg_in_a11(jpeg_in_a11) ,.jpeg_in_a12(jpeg_in_a12) ,.jpeg_in_a13(jpeg_in_a13) ,
	.jpeg_in_a14(jpeg_in_a14) ,.jpeg_in_a15(jpeg_in_a15) ,.jpeg_in_a16(jpeg_in_a16) ,
	.jpeg_in_a17(jpeg_in_a17) ,.jpeg_in_a18(jpeg_in_a18) ,.jpeg_in_a19(jpeg_in_a19) ,
	.jpeg_in_a20(jpeg_in_a20) ,.jpeg_in_a21(jpeg_in_a21) ,.jpeg_in_a22(jpeg_in_a22) ,
	.jpeg_in_a23(jpeg_in_a23) ,.jpeg_in_a24(jpeg_in_a24) ,.jpeg_in_a25(jpeg_in_a25) ,
	.jpeg_in_a26(jpeg_in_a26) ,.jpeg_in_a27(jpeg_in_a27) ,.jpeg_in_a28(jpeg_in_a28) ,
	.jpeg_in_a29(jpeg_in_a29) ,.jpeg_in_a30(jpeg_in_a30) ,.jpeg_in_a31(jpeg_in_a31) ,
	.jpeg_in_a32(jpeg_in_a32) ,.jpeg_in_a33(jpeg_in_a33) ,.jpeg_in_a34(jpeg_in_a34) ,
	.jpeg_in_a35(jpeg_in_a35) ,.jpeg_in_a36(jpeg_in_a36) ,.jpeg_in_a37(jpeg_in_a37) ,
	.jpeg_in_a38(jpeg_in_a38) ,.jpeg_in_a39(jpeg_in_a39) ,.jpeg_in_a40(jpeg_in_a40) ,
	.jpeg_in_a41(jpeg_in_a41) ,.jpeg_in_a42(jpeg_in_a42) ,.jpeg_in_a43(jpeg_in_a43) ,
	.jpeg_in_a44(jpeg_in_a44) ,.jpeg_in_a45(jpeg_in_a45) ,.jpeg_in_a46(jpeg_in_a46) ,
	.jpeg_in_a47(jpeg_in_a47) ,.jpeg_in_a48(jpeg_in_a48) ,.jpeg_in_a49(jpeg_in_a49) ,
	.jpeg_in_a50(jpeg_in_a50) ,.jpeg_in_a51(jpeg_in_a51) ,.jpeg_in_a52(jpeg_in_a52) ,
	.jpeg_in_a53(jpeg_in_a53) ,.jpeg_in_a54(jpeg_in_a54) ,.jpeg_in_a55(jpeg_in_a55) ,
	.jpeg_in_a56(jpeg_in_a56) ,.jpeg_in_a57(jpeg_in_a57) ,.jpeg_in_a58(jpeg_in_a58) ,
	.jpeg_in_a59(jpeg_in_a59) ,.jpeg_in_a60(jpeg_in_a60) ,.jpeg_in_a61(jpeg_in_a61) ,
	.jpeg_in_a62(jpeg_in_a62) ,.jpeg_in_a63(jpeg_in_a63) ,.jpeg_out_a00(jpeg_out_a00) ,
	.jpeg_out_a01(jpeg_out_a01) ,.jpeg_out_a02(jpeg_out_a02) ,.jpeg_out_a03(jpeg_out_a03) ,
	.jpeg_out_a04(jpeg_out_a04) ,.jpeg_out_a05(jpeg_out_a05) ,.jpeg_out_a06(jpeg_out_a06) ,
	.jpeg_out_a07(jpeg_out_a07) ,.jpeg_out_a08(jpeg_out_a08) ,.jpeg_out_a09(jpeg_out_a09) ,
	.jpeg_out_a10(jpeg_out_a10) ,.jpeg_out_a11(jpeg_out_a11) ,.jpeg_out_a12(jpeg_out_a12) ,
	.jpeg_out_a13(jpeg_out_a13) ,.jpeg_out_a14(jpeg_out_a14) ,.jpeg_out_a15(jpeg_out_a15) ,
	.jpeg_out_a16(jpeg_out_a16) ,.jpeg_out_a17(jpeg_out_a17) ,.jpeg_out_a18(jpeg_out_a18) ,
	.jpeg_out_a19(jpeg_out_a19) ,.jpeg_out_a20(jpeg_out_a20) ,.jpeg_out_a21(jpeg_out_a21) ,
	.jpeg_out_a22(jpeg_out_a22) ,.jpeg_out_a23(jpeg_out_a23) ,.jpeg_out_a24(jpeg_out_a24) ,
	.jpeg_out_a25(jpeg_out_a25) ,.jpeg_out_a26(jpeg_out_a26) ,.jpeg_out_a27(jpeg_out_a27) ,
	.jpeg_out_a28(jpeg_out_a28) ,.jpeg_out_a29(jpeg_out_a29) ,.jpeg_out_a30(jpeg_out_a30) ,
	.jpeg_out_a31(jpeg_out_a31) ,.jpeg_out_a32(jpeg_out_a32) ,.jpeg_out_a33(jpeg_out_a33) ,
	.jpeg_out_a34(jpeg_out_a34) ,.jpeg_out_a35(jpeg_out_a35) ,.jpeg_out_a36(jpeg_out_a36) ,
	.jpeg_out_a37(jpeg_out_a37) ,.jpeg_out_a38(jpeg_out_a38) ,.jpeg_out_a39(jpeg_out_a39) ,
	.jpeg_out_a40(jpeg_out_a40) ,.jpeg_out_a41(jpeg_out_a41) ,.jpeg_out_a42(jpeg_out_a42) ,
	.jpeg_out_a43(jpeg_out_a43) ,.jpeg_out_a44(jpeg_out_a44) ,.jpeg_out_a45(jpeg_out_a45) ,
	.jpeg_out_a46(jpeg_out_a46) ,.jpeg_out_a47(jpeg_out_a47) ,.jpeg_out_a48(jpeg_out_a48) ,
	.jpeg_out_a49(jpeg_out_a49) ,.jpeg_out_a50(jpeg_out_a50) ,.jpeg_out_a51(jpeg_out_a51) ,
	.jpeg_out_a52(jpeg_out_a52) ,.jpeg_out_a53(jpeg_out_a53) ,.jpeg_out_a54(jpeg_out_a54) ,
	.jpeg_out_a55(jpeg_out_a55) ,.jpeg_out_a56(jpeg_out_a56) ,.jpeg_out_a57(jpeg_out_a57) ,
	.jpeg_out_a58(jpeg_out_a58) ,.jpeg_out_a59(jpeg_out_a59) ,.jpeg_out_a60(jpeg_out_a60) ,
	.jpeg_out_a61(jpeg_out_a61) ,.jpeg_out_a62(jpeg_out_a62) ,.jpeg_out_a63(jpeg_out_a63) ,
	.jpeg_out_a64(jpeg_out_a64) ,.jpeg_out_a65(jpeg_out_a65) ,.jpeg_out_a66(jpeg_out_a66) ,
	.jpeg_out_a67(jpeg_out_a67) ,.jpeg_out_a68(jpeg_out_a68) ,.jpeg_out_a69(jpeg_out_a69) ,
	.jpeg_out_a70(jpeg_out_a70) ,.jpeg_out_a71(jpeg_out_a71) ,.jpeg_out_a72(jpeg_out_a72) ,
	.jpeg_out_a73(jpeg_out_a73) ,.jpeg_out_a74(jpeg_out_a74) ,.jpeg_out_a75(jpeg_out_a75) ,
	.jpeg_out_a76(jpeg_out_a76) ,.jpeg_out_a77(jpeg_out_a77) ,.jpeg_out_a78(jpeg_out_a78) ,
	.jpeg_out_a79(jpeg_out_a79) ,.jpeg_out_a80(jpeg_out_a80) ,.jpeg_out_a81(jpeg_out_a81) ,
	.jpeg_out_a82(jpeg_out_a82) ,.jpeg_out_a83(jpeg_out_a83) ,.jpeg_out_a84(jpeg_out_a84) ,
	.jpeg_out_a85(jpeg_out_a85) ,.jpeg_out_a86(jpeg_out_a86) ,.jpeg_out_a87(jpeg_out_a87) ,
	.jpeg_out_a88(jpeg_out_a88) ,.jpeg_out_a89(jpeg_out_a89) ,.jpeg_out_a90(jpeg_out_a90) ,
	.jpeg_out_a91(jpeg_out_a91) ,.jpeg_out_a92(jpeg_out_a92) ,.jpeg_out_a93(jpeg_out_a93) ,
	.jpeg_out_a94(jpeg_out_a94) ,.jpeg_out_a95(jpeg_out_a95) ,.jpeg_out_a96(jpeg_out_a96) ,
	.jpeg_out_a97(jpeg_out_a97) ,.jpeg_out_a98(jpeg_out_a98) ,.jpeg_out_a99(jpeg_out_a99) ,
	.jpeg_out_a100(jpeg_out_a100) ,.jpeg_out_a101(jpeg_out_a101) ,.jpeg_out_a102(jpeg_out_a102) ,
	.jpeg_out_a103(jpeg_out_a103) ,.jpeg_out_a104(jpeg_out_a104) ,.jpeg_out_a105(jpeg_out_a105) ,
	.jpeg_out_a106(jpeg_out_a106) ,.jpeg_out_a107(jpeg_out_a107) ,.jpeg_out_a108(jpeg_out_a108) ,
	.jpeg_out_a109(jpeg_out_a109) ,.jpeg_out_a110(jpeg_out_a110) ,.jpeg_out_a111(jpeg_out_a111) ,
	.jpeg_out_a112(jpeg_out_a112) ,.jpeg_out_a113(jpeg_out_a113) ,.jpeg_out_a114(jpeg_out_a114) ,
	.jpeg_out_a115(jpeg_out_a115) ,.jpeg_out_a116(jpeg_out_a116) ,.jpeg_out_a117(jpeg_out_a117) ,
	.jpeg_out_a118(jpeg_out_a118) ,.jpeg_out_a119(jpeg_out_a119) ,.jpeg_out_a120(jpeg_out_a120) ,
	.jpeg_out_a121(jpeg_out_a121) ,.jpeg_out_a122(jpeg_out_a122) ,.jpeg_out_a123(jpeg_out_a123) ,
	.jpeg_out_a124(jpeg_out_a124) ,.jpeg_out_a125(jpeg_out_a125) ,.jpeg_out_a126(jpeg_out_a126) ,
	.jpeg_out_a127(jpeg_out_a127) ,.jpeg_len_out(jpeg_len_out) ,.valid(valid) ,
	.ST1_56d(ST1_56d) ,.ST1_55d(ST1_55d) ,.ST1_54d(ST1_54d) ,.ST1_53d(ST1_53d) ,
	.ST1_52d(ST1_52d) ,.ST1_51d(ST1_51d) ,.ST1_50d(ST1_50d) ,.ST1_49d(ST1_49d) ,
	.ST1_48d(ST1_48d) ,.ST1_47d(ST1_47d) ,.ST1_46d(ST1_46d) ,.ST1_45d(ST1_45d) ,
	.ST1_44d(ST1_44d) ,.ST1_43d(ST1_43d) ,.ST1_42d(ST1_42d) ,.ST1_41d(ST1_41d) ,
	.ST1_40d(ST1_40d) ,.ST1_39d(ST1_39d) ,.ST1_38d(ST1_38d) ,.ST1_37d(ST1_37d) ,
	.ST1_36d(ST1_36d) ,.ST1_35d(ST1_35d) ,.ST1_34d(ST1_34d) ,.ST1_33d(ST1_33d) ,
	.ST1_32d(ST1_32d) ,.ST1_31d(ST1_31d) ,.ST1_30d(ST1_30d) ,.ST1_29d(ST1_29d) ,
	.ST1_28d(ST1_28d) ,.ST1_27d(ST1_27d) ,.ST1_26d(ST1_26d) ,.ST1_25d(ST1_25d) ,
	.ST1_24d(ST1_24d) ,.ST1_23d(ST1_23d) ,.ST1_22d(ST1_22d) ,.ST1_21d(ST1_21d) ,
	.ST1_20d(ST1_20d) ,.ST1_19d(ST1_19d) ,.ST1_18d(ST1_18d) ,.ST1_17d(ST1_17d) ,
	.ST1_16d(ST1_16d) ,.ST1_15d(ST1_15d) ,.ST1_14d(ST1_14d) ,.ST1_13d(ST1_13d) ,
	.ST1_12d(ST1_12d) ,.ST1_11d(ST1_11d) ,.ST1_10d(ST1_10d) ,.ST1_09d(ST1_09d) ,
	.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,
	.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,
	.JF_01(JF_01) ,.lop8u_11ot_port(lop8u_11ot) ,.JF_03(JF_03) ,.CT_31_port(CT_31) ,
	.JF_05_port(JF_05) ,.FL01_01_Leos_all(FL01_01_Leos_all) ,.FL02_01_Leos_all(FL02_01_Leos_all) );

endmodule

module jpeg_fsm ( clk ,rst ,ST1_56d ,ST1_55d ,ST1_54d ,ST1_53d ,ST1_52d ,ST1_51d ,
	ST1_50d ,ST1_49d ,ST1_48d ,ST1_47d ,ST1_46d ,ST1_45d ,ST1_44d ,ST1_43d ,
	ST1_42d ,ST1_41d ,ST1_40d ,ST1_39d ,ST1_38d ,ST1_37d ,ST1_36d ,ST1_35d ,
	ST1_34d ,ST1_33d ,ST1_32d ,ST1_31d ,ST1_30d ,ST1_29d ,ST1_28d ,ST1_27d ,
	ST1_26d ,ST1_25d ,ST1_24d ,ST1_23d ,ST1_22d ,ST1_21d ,ST1_20d ,ST1_19d ,
	ST1_18d ,ST1_17d ,ST1_16d ,ST1_15d ,ST1_14d ,ST1_13d ,ST1_12d ,ST1_11d ,
	ST1_10d ,ST1_09d ,ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,
	ST1_02d ,ST1_01d ,JF_01 ,lop8u_11ot ,JF_03 ,CT_31 ,JF_05 ,FL01_01_Leos_all ,
	FL02_01_Leos_all );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
output		ST1_56d ;
output		ST1_55d ;
output		ST1_54d ;
output		ST1_53d ;
output		ST1_52d ;
output		ST1_51d ;
output		ST1_50d ;
output		ST1_49d ;
output		ST1_48d ;
output		ST1_47d ;
output		ST1_46d ;
output		ST1_45d ;
output		ST1_44d ;
output		ST1_43d ;
output		ST1_42d ;
output		ST1_41d ;
output		ST1_40d ;
output		ST1_39d ;
output		ST1_38d ;
output		ST1_37d ;
output		ST1_36d ;
output		ST1_35d ;
output		ST1_34d ;
output		ST1_33d ;
output		ST1_32d ;
output		ST1_31d ;
output		ST1_30d ;
output		ST1_29d ;
output		ST1_28d ;
output		ST1_27d ;
output		ST1_26d ;
output		ST1_25d ;
output		ST1_24d ;
output		ST1_23d ;
output		ST1_22d ;
output		ST1_21d ;
output		ST1_20d ;
output		ST1_19d ;
output		ST1_18d ;
output		ST1_17d ;
output		ST1_16d ;
output		ST1_15d ;
output		ST1_14d ;
output		ST1_13d ;
output		ST1_12d ;
output		ST1_11d ;
output		ST1_10d ;
output		ST1_09d ;
output		ST1_08d ;
output		ST1_07d ;
output		ST1_06d ;
output		ST1_05d ;
output		ST1_04d ;
output		ST1_03d ;
output		ST1_02d ;
output		ST1_01d ;
input		JF_01 ;
input		lop8u_11ot ;
input		JF_03 ;
input		CT_31 ;
input		JF_05 ;
input		FL01_01_Leos_all ;
input		FL02_01_Leos_all ;
reg	[5:0]	B01_streg ;

parameter	ST1_01 = 6'h00 ;
parameter	ST1_02 = 6'h01 ;
parameter	ST1_03 = 6'h02 ;
parameter	ST1_04 = 6'h03 ;
parameter	ST1_05 = 6'h04 ;
parameter	ST1_06 = 6'h05 ;
parameter	ST1_07 = 6'h06 ;
parameter	ST1_08 = 6'h07 ;
parameter	ST1_09 = 6'h08 ;
parameter	ST1_10 = 6'h09 ;
parameter	ST1_11 = 6'h0a ;
parameter	ST1_12 = 6'h0b ;
parameter	ST1_13 = 6'h0c ;
parameter	ST1_14 = 6'h0d ;
parameter	ST1_15 = 6'h0e ;
parameter	ST1_16 = 6'h0f ;
parameter	ST1_17 = 6'h10 ;
parameter	ST1_18 = 6'h11 ;
parameter	ST1_19 = 6'h12 ;
parameter	ST1_20 = 6'h13 ;
parameter	ST1_21 = 6'h14 ;
parameter	ST1_22 = 6'h15 ;
parameter	ST1_23 = 6'h16 ;
parameter	ST1_24 = 6'h17 ;
parameter	ST1_25 = 6'h18 ;
parameter	ST1_26 = 6'h19 ;
parameter	ST1_27 = 6'h1a ;
parameter	ST1_28 = 6'h1b ;
parameter	ST1_29 = 6'h1c ;
parameter	ST1_30 = 6'h1d ;
parameter	ST1_31 = 6'h1e ;
parameter	ST1_32 = 6'h1f ;
parameter	ST1_33 = 6'h20 ;
parameter	ST1_34 = 6'h21 ;
parameter	ST1_35 = 6'h22 ;
parameter	ST1_36 = 6'h23 ;
parameter	ST1_37 = 6'h24 ;
parameter	ST1_38 = 6'h25 ;
parameter	ST1_39 = 6'h26 ;
parameter	ST1_40 = 6'h27 ;
parameter	ST1_41 = 6'h28 ;
parameter	ST1_42 = 6'h29 ;
parameter	ST1_43 = 6'h2a ;
parameter	ST1_44 = 6'h2b ;
parameter	ST1_45 = 6'h2c ;
parameter	ST1_46 = 6'h2d ;
parameter	ST1_47 = 6'h2e ;
parameter	ST1_48 = 6'h2f ;
parameter	ST1_49 = 6'h30 ;
parameter	ST1_50 = 6'h31 ;
parameter	ST1_51 = 6'h32 ;
parameter	ST1_52 = 6'h33 ;
parameter	ST1_53 = 6'h34 ;
parameter	ST1_54 = 6'h35 ;
parameter	ST1_55 = 6'h36 ;
parameter	ST1_56 = 6'h37 ;

assign	ST1_01d = ( ( B01_streg == ST1_01 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_02d = ( ( B01_streg == ST1_02 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_03d = ( ( B01_streg == ST1_03 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_04d = ( ( B01_streg == ST1_04 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_05d = ( ( B01_streg == ST1_05 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_06d = ( ( B01_streg == ST1_06 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_07d = ( ( B01_streg == ST1_07 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_08d = ( ( B01_streg == ST1_08 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_09d = ( ( B01_streg == ST1_09 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_10d = ( ( B01_streg == ST1_10 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_11d = ( ( B01_streg == ST1_11 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_12d = ( ( B01_streg == ST1_12 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_13d = ( ( B01_streg == ST1_13 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_14d = ( ( B01_streg == ST1_14 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_15d = ( ( B01_streg == ST1_15 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_16d = ( ( B01_streg == ST1_16 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_17d = ( ( B01_streg == ST1_17 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_18d = ( ( B01_streg == ST1_18 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_19d = ( ( B01_streg == ST1_19 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_20d = ( ( B01_streg == ST1_20 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_21d = ( ( B01_streg == ST1_21 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_22d = ( ( B01_streg == ST1_22 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_23d = ( ( B01_streg == ST1_23 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_24d = ( ( B01_streg == ST1_24 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_25d = ( ( B01_streg == ST1_25 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_26d = ( ( B01_streg == ST1_26 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_27d = ( ( B01_streg == ST1_27 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_28d = ( ( B01_streg == ST1_28 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_29d = ( ( B01_streg == ST1_29 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_30d = ( ( B01_streg == ST1_30 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_31d = ( ( B01_streg == ST1_31 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_32d = ( ( B01_streg == ST1_32 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_33d = ( ( B01_streg == ST1_33 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_34d = ( ( B01_streg == ST1_34 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_35d = ( ( B01_streg == ST1_35 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_36d = ( ( B01_streg == ST1_36 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_37d = ( ( B01_streg == ST1_37 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_38d = ( ( B01_streg == ST1_38 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_39d = ( ( B01_streg == ST1_39 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_40d = ( ( B01_streg == ST1_40 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_41d = ( ( B01_streg == ST1_41 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_42d = ( ( B01_streg == ST1_42 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_43d = ( ( B01_streg == ST1_43 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_44d = ( ( B01_streg == ST1_44 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_45d = ( ( B01_streg == ST1_45 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_46d = ( ( B01_streg == ST1_46 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_47d = ( ( B01_streg == ST1_47 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_48d = ( ( B01_streg == ST1_48 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_49d = ( ( B01_streg == ST1_49 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_50d = ( ( B01_streg == ST1_50 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_51d = ( ( B01_streg == ST1_51 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_52d = ( ( B01_streg == ST1_52 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_53d = ( ( B01_streg == ST1_53 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_54d = ( ( B01_streg == ST1_54 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_55d = ( ( B01_streg == ST1_55 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_56d = ( ( B01_streg == ST1_56 ) ? 1'h1 : 1'h0 ) ;
always @ ( posedge clk )
	if ( !rst )
		B01_streg <= ST1_01 ;
	else
		case ( B01_streg )
		ST1_01 :
			B01_streg <= ST1_02 ;
		ST1_02 :
			if ( ( JF_01 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_03 ;
		ST1_03 :
			if ( ( lop8u_11ot != 1'h0 ) )
				B01_streg <= ST1_03 ;
			else
				B01_streg <= ST1_04 ;
		ST1_04 :
			if ( ( JF_03 != 1'h0 ) )
				B01_streg <= ST1_04 ;
			else
				B01_streg <= ST1_05 ;
		ST1_05 :
			B01_streg <= ST1_06 ;
		ST1_06 :
			if ( ( CT_31 != 1'h0 ) )
				B01_streg <= ST1_10 ;
			else
				B01_streg <= ST1_07 ;
		ST1_07 :
			B01_streg <= ST1_08 ;
		ST1_08 :
			if ( ( JF_05 != 1'h0 ) )
				B01_streg <= ST1_09 ;
			else
				B01_streg <= ST1_11 ;
		ST1_09 :
			B01_streg <= ST1_11 ;
		ST1_10 :
			if ( ( FL01_01_Leos_all != 1'h0 ) )
				B01_streg <= ST1_12 ;
			else
				B01_streg <= ST1_10 ;
		ST1_11 :
			if ( ( FL02_01_Leos_all != 1'h0 ) )
				B01_streg <= ST1_14 ;
			else
				B01_streg <= ST1_11 ;
		ST1_12 :
			B01_streg <= ST1_13 ;
		ST1_13 :
			B01_streg <= ST1_06 ;
		ST1_14 :
			B01_streg <= ST1_15 ;
		ST1_15 :
			B01_streg <= ST1_16 ;
		ST1_16 :
			B01_streg <= ST1_17 ;
		ST1_17 :
			B01_streg <= ST1_18 ;
		ST1_18 :
			B01_streg <= ST1_19 ;
		ST1_19 :
			B01_streg <= ST1_20 ;
		ST1_20 :
			B01_streg <= ST1_21 ;
		ST1_21 :
			B01_streg <= ST1_22 ;
		ST1_22 :
			B01_streg <= ST1_23 ;
		ST1_23 :
			B01_streg <= ST1_24 ;
		ST1_24 :
			B01_streg <= ST1_25 ;
		ST1_25 :
			B01_streg <= ST1_26 ;
		ST1_26 :
			B01_streg <= ST1_27 ;
		ST1_27 :
			B01_streg <= ST1_28 ;
		ST1_28 :
			B01_streg <= ST1_29 ;
		ST1_29 :
			B01_streg <= ST1_30 ;
		ST1_30 :
			B01_streg <= ST1_31 ;
		ST1_31 :
			B01_streg <= ST1_32 ;
		ST1_32 :
			B01_streg <= ST1_33 ;
		ST1_33 :
			B01_streg <= ST1_34 ;
		ST1_34 :
			B01_streg <= ST1_35 ;
		ST1_35 :
			B01_streg <= ST1_36 ;
		ST1_36 :
			B01_streg <= ST1_37 ;
		ST1_37 :
			B01_streg <= ST1_38 ;
		ST1_38 :
			B01_streg <= ST1_39 ;
		ST1_39 :
			B01_streg <= ST1_40 ;
		ST1_40 :
			B01_streg <= ST1_41 ;
		ST1_41 :
			B01_streg <= ST1_42 ;
		ST1_42 :
			B01_streg <= ST1_43 ;
		ST1_43 :
			B01_streg <= ST1_44 ;
		ST1_44 :
			B01_streg <= ST1_45 ;
		ST1_45 :
			B01_streg <= ST1_46 ;
		ST1_46 :
			B01_streg <= ST1_47 ;
		ST1_47 :
			B01_streg <= ST1_48 ;
		ST1_48 :
			B01_streg <= ST1_49 ;
		ST1_49 :
			B01_streg <= ST1_50 ;
		ST1_50 :
			B01_streg <= ST1_51 ;
		ST1_51 :
			B01_streg <= ST1_52 ;
		ST1_52 :
			B01_streg <= ST1_53 ;
		ST1_53 :
			B01_streg <= ST1_54 ;
		ST1_54 :
			B01_streg <= ST1_55 ;
		ST1_55 :
			B01_streg <= ST1_56 ;
		ST1_56 :
			B01_streg <= ST1_02 ;
		default :
			B01_streg <= ST1_01 ;
		endcase

endmodule

module jpeg_dat ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,
	jpeg_in_a04 ,jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,
	jpeg_in_a10 ,jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,
	jpeg_in_a16 ,jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,
	jpeg_in_a22 ,jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,
	jpeg_in_a28 ,jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,
	jpeg_in_a34 ,jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,
	jpeg_in_a40 ,jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,
	jpeg_in_a46 ,jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,
	jpeg_in_a52 ,jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,
	jpeg_in_a58 ,jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,
	jpeg_out_a00 ,jpeg_out_a01 ,jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,
	jpeg_out_a06 ,jpeg_out_a07 ,jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,
	jpeg_out_a12 ,jpeg_out_a13 ,jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,
	jpeg_out_a18 ,jpeg_out_a19 ,jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,
	jpeg_out_a24 ,jpeg_out_a25 ,jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,
	jpeg_out_a30 ,jpeg_out_a31 ,jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,
	jpeg_out_a36 ,jpeg_out_a37 ,jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,
	jpeg_out_a42 ,jpeg_out_a43 ,jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,
	jpeg_out_a48 ,jpeg_out_a49 ,jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,
	jpeg_out_a54 ,jpeg_out_a55 ,jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,
	jpeg_out_a60 ,jpeg_out_a61 ,jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,
	jpeg_out_a66 ,jpeg_out_a67 ,jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,
	jpeg_out_a72 ,jpeg_out_a73 ,jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,
	jpeg_out_a78 ,jpeg_out_a79 ,jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,
	jpeg_out_a84 ,jpeg_out_a85 ,jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,
	jpeg_out_a90 ,jpeg_out_a91 ,jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,
	jpeg_out_a96 ,jpeg_out_a97 ,jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,
	jpeg_out_a102 ,jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,
	jpeg_out_a107 ,jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,
	jpeg_out_a112 ,jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,
	jpeg_out_a117 ,jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,
	jpeg_out_a122 ,jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,
	jpeg_out_a127 ,jpeg_len_out ,valid ,ST1_56d ,ST1_55d ,ST1_54d ,ST1_53d ,
	ST1_52d ,ST1_51d ,ST1_50d ,ST1_49d ,ST1_48d ,ST1_47d ,ST1_46d ,ST1_45d ,
	ST1_44d ,ST1_43d ,ST1_42d ,ST1_41d ,ST1_40d ,ST1_39d ,ST1_38d ,ST1_37d ,
	ST1_36d ,ST1_35d ,ST1_34d ,ST1_33d ,ST1_32d ,ST1_31d ,ST1_30d ,ST1_29d ,
	ST1_28d ,ST1_27d ,ST1_26d ,ST1_25d ,ST1_24d ,ST1_23d ,ST1_22d ,ST1_21d ,
	ST1_20d ,ST1_19d ,ST1_18d ,ST1_17d ,ST1_16d ,ST1_15d ,ST1_14d ,ST1_13d ,
	ST1_12d ,ST1_11d ,ST1_10d ,ST1_09d ,ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,
	ST1_04d ,ST1_03d ,ST1_02d ,ST1_01d ,JF_01 ,lop8u_11ot_port ,JF_03 ,CT_31_port ,
	JF_05_port ,FL01_01_Leos_all ,FL02_01_Leos_all );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
input		ST1_56d ;
input		ST1_55d ;
input		ST1_54d ;
input		ST1_53d ;
input		ST1_52d ;
input		ST1_51d ;
input		ST1_50d ;
input		ST1_49d ;
input		ST1_48d ;
input		ST1_47d ;
input		ST1_46d ;
input		ST1_45d ;
input		ST1_44d ;
input		ST1_43d ;
input		ST1_42d ;
input		ST1_41d ;
input		ST1_40d ;
input		ST1_39d ;
input		ST1_38d ;
input		ST1_37d ;
input		ST1_36d ;
input		ST1_35d ;
input		ST1_34d ;
input		ST1_33d ;
input		ST1_32d ;
input		ST1_31d ;
input		ST1_30d ;
input		ST1_29d ;
input		ST1_28d ;
input		ST1_27d ;
input		ST1_26d ;
input		ST1_25d ;
input		ST1_24d ;
input		ST1_23d ;
input		ST1_22d ;
input		ST1_21d ;
input		ST1_20d ;
input		ST1_19d ;
input		ST1_18d ;
input		ST1_17d ;
input		ST1_16d ;
input		ST1_15d ;
input		ST1_14d ;
input		ST1_13d ;
input		ST1_12d ;
input		ST1_11d ;
input		ST1_10d ;
input		ST1_09d ;
input		ST1_08d ;
input		ST1_07d ;
input		ST1_06d ;
input		ST1_05d ;
input		ST1_04d ;
input		ST1_03d ;
input		ST1_02d ;
input		ST1_01d ;
output		JF_01 ;
output		lop8u_11ot_port ;
output		JF_03 ;
output		CT_31_port ;
output		JF_05_port ;
output		FL01_01_Leos_all ;
output		FL02_01_Leos_all ;
wire		M_171 ;
wire		M_170 ;
wire		M_168 ;
wire		M_167 ;
wire		M_165 ;
wire		M_163 ;
wire		M_162 ;
wire		M_161 ;
wire		M_160 ;
wire		M_159 ;
wire		M_158 ;
wire		M_157 ;
wire		M_156 ;
wire		M_155 ;
wire		M_154 ;
wire		M_153 ;
wire		M_152 ;
wire		M_151 ;
wire		M_150 ;
wire		M_149 ;
wire		M_148 ;
wire		M_147 ;
wire		M_146 ;
wire		M_145 ;
wire		M_144 ;
wire		M_143 ;
wire		M_142 ;
wire		M_141 ;
wire		M_140 ;
wire		M_139 ;
wire		M_138 ;
wire		M_137 ;
wire		M_136 ;
wire		M_135 ;
wire		M_134 ;
wire		M_133 ;
wire		M_132 ;
wire		M_131 ;
wire		M_130 ;
wire		M_129 ;
wire		M_128 ;
wire		M_127 ;
wire		M_126 ;
wire		M_125 ;
wire		M_124 ;
wire		M_123 ;
wire		M_122 ;
wire		M_120 ;
wire		M_117 ;
wire		M_116 ;
wire		M_113 ;
wire		M_112 ;
wire		M_110 ;
wire		U_237 ;
wire		U_236 ;
wire		U_235 ;
wire		U_234 ;
wire		U_230 ;
wire		U_228 ;
wire		U_223 ;
wire		U_219 ;
wire		U_218 ;
wire		U_213 ;
wire		U_212 ;
wire		U_207 ;
wire		U_204 ;
wire		U_202 ;
wire		U_198 ;
wire		U_196 ;
wire		U_193 ;
wire		U_189 ;
wire		U_188 ;
wire		U_180 ;
wire		U_177 ;
wire		U_176 ;
wire		U_173 ;
wire		U_171 ;
wire		U_166 ;
wire		U_165 ;
wire		U_164 ;
wire		U_163 ;
wire		U_162 ;
wire		C_04 ;
wire		U_161 ;
wire		U_96 ;
wire		U_95 ;
wire		U_94 ;
wire		U_93 ;
wire		U_92 ;
wire		U_91 ;
wire		U_90 ;
wire		U_89 ;
wire		U_87 ;
wire		U_84 ;
wire		U_83 ;
wire		U_82 ;
wire		U_81 ;
wire		U_80 ;
wire		C_02 ;
wire		U_79 ;
wire		U_14 ;
wire		U_13 ;
wire		U_12 ;
wire		U_11 ;
wire		U_10 ;
wire		U_09 ;
wire		U_08 ;
wire		U_07 ;
wire		U_06 ;
wire		U_05 ;
wire	[1:0]	sub8u_7_11i2 ;
wire	[6:0]	sub8u_7_11i1 ;
wire	[6:0]	sub8u_7_11ot ;
wire	[2:0]	sub8u_71i2 ;
wire	[6:0]	sub8u_71i1 ;
wire	[6:0]	sub8u_71ot ;
wire	[31:0]	decr32s2i1 ;
wire	[31:0]	decr32s2ot ;
wire	[31:0]	decr32s1i1 ;
wire	[31:0]	decr32s1ot ;
wire	[6:0]	decr8u_71i1 ;
wire	[6:0]	decr8u_71ot ;
wire	[31:0]	incr32s3i1 ;
wire	[31:0]	incr32s3ot ;
wire	[31:0]	incr32s2i1 ;
wire	[31:0]	incr32s2ot ;
wire	[31:0]	incr32s1i1 ;
wire	[31:0]	incr32s1ot ;
wire	[7:0]	incr8u2ot ;
wire	[7:0]	incr8u1i1 ;
wire	[7:0]	incr8u1ot ;
wire	[3:0]	incr4s1i1 ;
wire	[3:0]	incr4s1ot ;
wire	[5:0]	lop8u_11i2 ;
wire	[5:0]	lop8u_11i1 ;
wire		lop8u_11ot ;
wire	[8:0]	sub12s_91i2 ;
wire	[8:0]	sub12s_91i1 ;
wire	[8:0]	sub12s_91ot ;
wire	[1:0]	sub8u1i2 ;
wire	[7:0]	sub8u1i1 ;
wire	[7:0]	sub8u1ot ;
wire		FL02_02_ndat ;
wire		FL02_01_ndat ;
wire		FL02_03_eos ;
wire		FL02_02_eos ;
wire		FL02_01_eos ;
wire		FL02_01_Leos_all ;
wire		FJ_14_17 ;
wire		FL02_03_01a ;
wire		FL02_02_01a ;
wire		FL02_01_01a ;
wire		FL02_03_break ;
wire		FL01_01_ndat ;
wire		FL01_02_eos ;
wire		FL01_01_eos ;
wire		FL01_01_Leos_all ;
wire		FJ_11_15 ;
wire		FL01_02_01a ;
wire		FL01_01_01a ;
wire		FL01_02_break ;
wire		CT_35 ;
wire		CT_31 ;
wire		JF_05 ;
wire		CT_26 ;
wire		JF_03 ;
wire		CT_12 ;
wire		JF_01 ;
wire		zz_WE2 ;
wire		rl_WE1 ;
wire	[8:0]	rl_RD1 ;
wire	[8:0]	rl_RD2 ;
wire	[8:0]	rl_RD3 ;
wire	[8:0]	zz_RD1 ;
wire		RG_previous_dc_en ;
wire		RG_quantized_block_en ;
wire		RG_quantized_block_1_en ;
wire		RG_quantized_block_2_en ;
wire		RG_quantized_block_3_en ;
wire		RG_quantized_block_4_en ;
wire		RG_quantized_block_5_en ;
wire		RG_quantized_block_6_en ;
wire		RG_quantized_block_7_en ;
wire		RG_quantized_block_8_en ;
wire		RG_quantized_block_9_en ;
wire		RG_quantized_block_10_en ;
wire		RG_quantized_block_11_en ;
wire		RG_quantized_block_12_en ;
wire		RG_quantized_block_13_en ;
wire		RG_quantized_block_14_en ;
wire		RG_quantized_block_15_en ;
wire		RG_quantized_block_16_en ;
wire		RG_quantized_block_17_en ;
wire		RG_quantized_block_18_en ;
wire		RG_quantized_block_19_en ;
wire		RG_quantized_block_20_en ;
wire		RG_quantized_block_21_en ;
wire		RG_quantized_block_22_en ;
wire		RG_quantized_block_23_en ;
wire		RG_quantized_block_24_en ;
wire		RG_quantized_block_25_en ;
wire		RG_quantized_block_26_en ;
wire		RG_quantized_block_27_en ;
wire		RG_quantized_block_28_en ;
wire		RG_quantized_block_29_en ;
wire		RG_quantized_block_30_en ;
wire		RG_quantized_block_31_en ;
wire		RG_quantized_block_32_en ;
wire		RG_quantized_block_33_en ;
wire		RG_quantized_block_34_en ;
wire		RG_quantized_block_35_en ;
wire		RG_quantized_block_36_en ;
wire		RG_quantized_block_37_en ;
wire		RG_quantized_block_38_en ;
wire		RG_quantized_block_39_en ;
wire		RG_quantized_block_40_en ;
wire		RG_quantized_block_41_en ;
wire		RG_quantized_block_42_en ;
wire		RG_quantized_block_43_en ;
wire		RG_quantized_block_44_en ;
wire		RG_quantized_block_45_en ;
wire		RG_quantized_block_46_en ;
wire		RG_quantized_block_47_en ;
wire		RG_quantized_block_48_en ;
wire		RG_quantized_block_49_en ;
wire		RG_quantized_block_50_en ;
wire		RG_quantized_block_51_en ;
wire		RG_quantized_block_52_en ;
wire		RG_quantized_block_53_en ;
wire		RG_quantized_block_54_en ;
wire		RG_quantized_block_55_en ;
wire		RG_quantized_block_56_en ;
wire		RG_quantized_block_57_en ;
wire		RG_quantized_block_58_en ;
wire		RG_quantized_block_59_en ;
wire		FF_j_en ;
wire		FF_i_en ;
wire		RG_len_03_en ;
wire		RG_i_02_en ;
wire		jpeg_out_a00_r_en ;
wire		jpeg_out_a01_r_en ;
wire		jpeg_out_a02_r_en ;
wire		jpeg_out_a03_r_en ;
wire		jpeg_out_a04_r_en ;
wire		jpeg_out_a05_r_en ;
wire		jpeg_out_a06_r_en ;
wire		jpeg_out_a07_r_en ;
wire		jpeg_out_a08_r_en ;
wire		jpeg_out_a09_r_en ;
wire		jpeg_out_a10_r_en ;
wire		jpeg_out_a11_r_en ;
wire		jpeg_out_a12_r_en ;
wire		jpeg_out_a13_r_en ;
wire		jpeg_out_a14_r_en ;
wire		jpeg_out_a15_r_en ;
wire		jpeg_out_a16_r_en ;
wire		jpeg_out_a17_r_en ;
wire		jpeg_out_a18_r_en ;
wire		jpeg_out_a19_r_en ;
wire		jpeg_out_a20_r_en ;
wire		jpeg_out_a21_r_en ;
wire		jpeg_out_a22_r_en ;
wire		jpeg_out_a23_r_en ;
wire		jpeg_out_a24_r_en ;
wire		jpeg_out_a25_r_en ;
wire		jpeg_out_a26_r_en ;
wire		jpeg_out_a27_r_en ;
wire		jpeg_out_a28_r_en ;
wire		jpeg_out_a29_r_en ;
wire		jpeg_out_a30_r_en ;
wire		jpeg_out_a31_r_en ;
wire		jpeg_out_a32_r_en ;
wire		jpeg_out_a33_r_en ;
wire		jpeg_out_a34_r_en ;
wire		jpeg_out_a35_r_en ;
wire		jpeg_out_a36_r_en ;
wire		jpeg_out_a37_r_en ;
wire		jpeg_out_a38_r_en ;
wire		jpeg_out_a39_r_en ;
wire		jpeg_out_a40_r_en ;
wire		jpeg_out_a41_r_en ;
wire		jpeg_out_a42_r_en ;
wire		jpeg_out_a43_r_en ;
wire		jpeg_out_a44_r_en ;
wire		jpeg_out_a45_r_en ;
wire		jpeg_out_a46_r_en ;
wire		jpeg_out_a47_r_en ;
wire		jpeg_out_a48_r_en ;
wire		jpeg_out_a49_r_en ;
wire		jpeg_out_a50_r_en ;
wire		jpeg_out_a51_r_en ;
wire		jpeg_out_a52_r_en ;
wire		jpeg_out_a53_r_en ;
wire		jpeg_out_a54_r_en ;
wire		jpeg_out_a55_r_en ;
wire		jpeg_out_a56_r_en ;
wire		jpeg_out_a57_r_en ;
wire		jpeg_out_a58_r_en ;
wire		jpeg_out_a59_r_en ;
wire		jpeg_out_a60_r_en ;
wire		jpeg_out_a61_r_en ;
wire		jpeg_out_a62_r_en ;
wire		jpeg_out_a63_r_en ;
wire		jpeg_out_a64_r_en ;
wire		jpeg_out_a65_r_en ;
wire		jpeg_out_a66_r_en ;
wire		jpeg_out_a67_r_en ;
wire		jpeg_out_a68_r_en ;
wire		jpeg_out_a69_r_en ;
wire		jpeg_out_a70_r_en ;
wire		jpeg_out_a71_r_en ;
wire		jpeg_out_a72_r_en ;
wire		jpeg_out_a73_r_en ;
wire		jpeg_out_a74_r_en ;
wire		jpeg_out_a75_r_en ;
wire		jpeg_out_a76_r_en ;
wire		jpeg_out_a77_r_en ;
wire		jpeg_out_a78_r_en ;
wire		jpeg_out_a79_r_en ;
wire		jpeg_out_a80_r_en ;
wire		jpeg_out_a81_r_en ;
wire		jpeg_out_a82_r_en ;
wire		jpeg_out_a83_r_en ;
wire		jpeg_out_a84_r_en ;
wire		jpeg_out_a85_r_en ;
wire		jpeg_out_a86_r_en ;
wire		jpeg_out_a87_r_en ;
wire		jpeg_out_a88_r_en ;
wire		jpeg_out_a89_r_en ;
wire		jpeg_out_a90_r_en ;
wire		jpeg_out_a91_r_en ;
wire		jpeg_out_a92_r_en ;
wire		jpeg_out_a93_r_en ;
wire		jpeg_out_a94_r_en ;
wire		jpeg_out_a95_r_en ;
wire		jpeg_out_a96_r_en ;
wire		jpeg_out_a97_r_en ;
wire		jpeg_out_a98_r_en ;
wire		jpeg_out_a99_r_en ;
wire		jpeg_out_a100_r_en ;
wire		jpeg_out_a101_r_en ;
wire		jpeg_out_a102_r_en ;
wire		jpeg_out_a103_r_en ;
wire		jpeg_out_a104_r_en ;
wire		jpeg_out_a105_r_en ;
wire		jpeg_out_a106_r_en ;
wire		jpeg_out_a107_r_en ;
wire		jpeg_out_a108_r_en ;
wire		jpeg_out_a109_r_en ;
wire		jpeg_out_a110_r_en ;
wire		jpeg_out_a111_r_en ;
wire		jpeg_out_a112_r_en ;
wire		jpeg_out_a113_r_en ;
wire		jpeg_out_a114_r_en ;
wire		jpeg_out_a115_r_en ;
wire		jpeg_out_a116_r_en ;
wire		jpeg_out_a117_r_en ;
wire		jpeg_out_a118_r_en ;
wire		jpeg_out_a119_r_en ;
wire		jpeg_out_a120_r_en ;
wire		jpeg_out_a121_r_en ;
wire		jpeg_out_a122_r_en ;
wire		jpeg_out_a123_r_en ;
wire		jpeg_out_a124_r_en ;
wire		jpeg_out_a125_r_en ;
wire		jpeg_out_a126_r_en ;
wire		jpeg_out_a127_r_en ;
wire		jpeg_len_out_r_en ;
wire		RG_j_03_en ;
wire		RG_i_k_01_en ;
wire		RG_i_j_01_en ;
wire		RG_k_quantized_block_02_en ;
wire		RG_quantized_block_rl_02_en ;
wire		RG_quantized_block_rl_02_1_en ;
wire		RG_previous_dc_quantized_block_en ;
wire		FF_d_en ;
wire		FF_len_en ;
wire		RG_len_01_1_en ;
wire		RG_82_01_en ;
wire		FL01_01_streg_en ;
wire		FL01_02_streg_en ;
wire		FL02_01_streg_en ;
wire		FL02_02_streg_en ;
wire		FL02_03_streg_en ;
wire		valid_r_en ;
reg	FL02_03_streg ;
reg	FL02_02_streg ;
reg	FL02_01_streg ;
reg	FL01_02_streg ;
reg	FL01_01_streg ;
reg	[8:0]	RG_previous_dc ;	// line#=../rle.h:66
reg	[3:0]	RG_j_03 ;	// line#=../rle.cpp:27
reg	[31:0]	RG_i_k_01 ;	// line#=../rle.cpp:25,105
reg	[31:0]	RG_i_j_01 ;	// line#=../rle.cpp:25,105
reg	[8:0]	RG_quantized_block ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_1 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_2 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_3 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_4 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_5 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_6 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_7 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_8 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_9 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_10 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_11 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_12 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_13 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_14 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_15 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_16 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_17 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_18 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_19 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_20 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_21 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_22 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_23 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_24 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_25 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_26 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_27 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_28 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_29 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_30 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_31 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_32 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_33 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_34 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_35 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_36 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_37 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_38 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_39 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_40 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_41 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_42 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_43 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_44 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_45 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_46 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_47 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_48 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_49 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_50 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_51 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_52 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_53 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_54 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_55 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_56 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_57 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_58 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_quantized_block_59 ;	// line#=../rle.cpp:22
reg	[8:0]	RG_k_quantized_block_02 ;	// line#=../rle.cpp:22,25
reg	[8:0]	RG_quantized_block_rl_02 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_02_1 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_previous_dc_quantized_block ;	// line#=../rle.cpp:22 ../rle.h:66
reg	[5:0]	RG_k ;	// line#=../rle.cpp:105
reg	FF_d ;	// line#=../rle.cpp:105
reg	FF_j ;	// line#=../rle.cpp:27
reg	FF_i ;	// line#=../rle.cpp:25
reg	FF_len ;	// line#=../rle.cpp:24
reg	[7:0]	RG_len_03 ;	// line#=../rle.cpp:24
reg	[7:0]	RG_len_02 ;	// line#=../rle.cpp:24
reg	[6:0]	RG_75_02 ;
reg	[7:0]	RG_len_01 ;	// line#=../rle.cpp:24
reg	[31:0]	RG_i_02 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_i_01 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_k_01 ;	// line#=../rle.cpp:25
reg	[6:0]	RG_80_01 ;
reg	[7:0]	RG_len_01_1 ;	// line#=../rle.cpp:24
reg	RG_82_01 ;
reg	[6:0]	RG_k_01_1 ;	// line#=../rle.cpp:105
reg	[8:0]	jpeg_out_a00_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a01_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a02_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a03_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a04_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a05_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a06_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a07_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a08_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a09_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a10_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a11_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a12_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a13_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a14_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a15_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a16_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a17_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a18_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a19_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a20_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a21_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a22_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a23_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a24_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a25_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a26_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a27_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a28_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a29_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a30_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a31_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a32_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a33_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a34_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a35_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a36_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a37_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a38_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a39_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a40_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a41_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a42_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a43_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a44_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a45_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a46_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a47_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a48_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a49_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a50_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a51_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a52_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a53_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a54_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a55_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a56_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a57_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a58_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a59_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a60_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a61_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a62_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a63_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a64_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a65_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a66_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a67_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a68_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a69_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a70_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a71_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a72_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a73_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a74_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a75_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a76_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a77_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a78_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a79_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a80_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a81_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a82_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a83_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a84_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a85_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a86_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a87_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a88_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a89_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a90_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a91_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a92_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a93_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a94_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a95_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a96_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a97_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a98_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a99_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a100_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a101_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a102_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a103_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a104_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a105_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a106_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a107_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a108_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a109_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a110_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a111_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a112_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a113_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a114_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a115_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a116_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a117_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a118_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a119_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a120_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a121_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a122_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a123_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a124_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a125_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a126_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a127_r ;	// line#=../rle.h:60
reg	[11:0]	jpeg_len_out_r ;	// line#=../rle.h:61
reg	valid_r ;	// line#=../rle.h:62
reg	M_02_t1 ;
reg	M_01_t1 ;
reg	M_03_t1 ;
reg	FL01_01_next ;
reg	FL02_01_next ;
reg	[3:0]	RG_j_03_t ;
reg	[2:0]	TR_01 ;
reg	[31:0]	RG_i_k_01_t ;
reg	RG_i_k_01_t_c1 ;
reg	RG_i_k_01_t_c2 ;
reg	RG_i_k_01_t_c3 ;
reg	TR_02 ;
reg	[31:0]	RG_i_j_01_t ;
reg	RG_i_j_01_t_c1 ;
reg	RG_i_j_01_t_c2 ;
reg	RG_i_j_01_t_c3 ;
reg	[8:0]	RG_k_quantized_block_02_t ;
reg	[8:0]	RG_quantized_block_rl_02_t ;
reg	[8:0]	RG_quantized_block_rl_02_1_t ;
reg	[8:0]	RG_previous_dc_quantized_block_t ;
reg	[5:0]	RG_k_t ;
reg	FF_d_t ;
reg	FF_d_t_c1 ;
reg	FF_d_t_c2 ;
reg	FF_len_t ;
reg	[6:0]	RG_80_01_t ;
reg	[7:0]	RG_len_01_1_t ;
reg	RG_82_01_t ;
reg	[6:0]	RG_k_01_1_t ;
reg	FL01_01_streg_t ;
reg	FL01_01_streg_t_c1 ;
reg	FL01_02_streg_t ;
reg	FL01_02_streg_t_c1 ;
reg	FL01_02_streg_t_c2 ;
reg	FL02_01_streg_t ;
reg	FL02_01_streg_t_c1 ;
reg	FL02_02_streg_t ;
reg	FL02_02_streg_t_c1 ;
reg	FL02_02_streg_t_c2 ;
reg	FL02_03_streg_t ;
reg	FL02_03_streg_t_c1 ;
reg	FL02_03_streg_t_c2 ;
reg	valid_r_t ;
reg	[5:0]	TR_04 ;
reg	[7:0]	incr8u2i1 ;
reg	incr8u2i1_c1 ;
reg	incr8u2i1_c2 ;
reg	[5:0]	zz_RA1 ;
reg	zz_RA1_c1 ;
reg	[5:0]	zz_WA2 ;
reg	zz_WA2_c1 ;
reg	zz_WA2_c2 ;
reg	[8:0]	TR_44 ;
reg	[8:0]	TR_45 ;
reg	[8:0]	TR_46 ;
reg	[8:0]	TR_47 ;
reg	[8:0]	TR_48 ;
reg	[8:0]	TR_49 ;
reg	[8:0]	TR_50 ;
reg	[8:0]	TR_51 ;
reg	[8:0]	zz_WD2 ;
reg	[1:0]	M_172 ;
reg	[1:0]	TR_17 ;
reg	[2:0]	TR_18 ;
reg	[3:0]	TR_06 ;
reg	TR_06_c1 ;
reg	[2:0]	TR_19 ;
reg	[2:0]	TR_32 ;
reg	[3:0]	TR_20 ;
reg	TR_20_c1 ;
reg	[4:0]	TR_07 ;
reg	TR_07_c1 ;
reg	[1:0]	TR_21 ;
reg	[2:0]	TR_22 ;
reg	[2:0]	TR_33 ;
reg	[3:0]	TR_23 ;
reg	TR_23_c1 ;
reg	[2:0]	TR_34 ;
reg	[1:0]	TR_41 ;
reg	[2:0]	TR_42 ;
reg	[3:0]	TR_35 ;
reg	TR_35_c1 ;
reg	[4:0]	TR_24 ;
reg	TR_24_c1 ;
reg	[5:0]	TR_08 ;
reg	TR_08_c1 ;
reg	[2:0]	TR_09 ;
reg	[2:0]	TR_25 ;
reg	[3:0]	TR_10 ;
reg	TR_10_c1 ;
reg	[1:0]	TR_26 ;
reg	[2:0]	TR_27 ;
reg	[2:0]	TR_36 ;
reg	[3:0]	TR_28 ;
reg	TR_28_c1 ;
reg	[4:0]	TR_11 ;
reg	TR_11_c1 ;
reg	[2:0]	TR_29 ;
reg	[1:0]	TR_37 ;
reg	[2:0]	TR_38 ;
reg	[3:0]	TR_30 ;
reg	TR_30_c1 ;
reg	[2:0]	TR_39 ;
reg	[2:0]	TR_43 ;
reg	[3:0]	TR_40 ;
reg	TR_40_c1 ;
reg	[4:0]	TR_31 ;
reg	TR_31_c1 ;
reg	[5:0]	TR_12 ;
reg	TR_12_c1 ;
reg	[6:0]	rl_AD1 ;
reg	rl_AD1_c1 ;
reg	rl_AD1_c2 ;
reg	rl_AD1_c3 ;
reg	[8:0]	rl_WD1 ;
reg	[5:0]	TR_13 ;
reg	[5:0]	TR_14 ;
reg	[6:0]	rl_RA2 ;
reg	rl_RA2_c1 ;
reg	[5:0]	TR_15 ;
reg	[5:0]	TR_16 ;
reg	[6:0]	rl_RA3 ;

jpeg_sub8u_7_1 INST_sub8u_7_1_1 ( .i1(sub8u_7_11i1) ,.i2(sub8u_7_11i2) ,.o1(sub8u_7_11ot) );	// line#=../rle.cpp:83,84
jpeg_sub8u_7 INST_sub8u_7_1 ( .i1(sub8u_71i1) ,.i2(sub8u_71i2) ,.o1(sub8u_71ot) );	// line#=../rle.cpp:83,84
jpeg_decr32s INST_decr32s_1 ( .i1(decr32s1i1) ,.o1(decr32s1ot) );	// line#=../rle.cpp:124,155
jpeg_decr32s INST_decr32s_2 ( .i1(decr32s2i1) ,.o1(decr32s2ot) );	// line#=../rle.cpp:130,161
jpeg_decr8u_7 INST_decr8u_7_1 ( .i1(decr8u_71i1) ,.o1(decr8u_71ot) );	// line#=../rle.cpp:77,78
jpeg_incr32s INST_incr32s_1 ( .i1(incr32s1i1) ,.o1(incr32s1ot) );	// line#=../rle.cpp:61,62,63,114,125,145
									// ,156
jpeg_incr32s INST_incr32s_2 ( .i1(incr32s2i1) ,.o1(incr32s2ot) );	// line#=../rle.cpp:64,119,129,150,160
jpeg_incr32s INST_incr32s_3 ( .i1(incr32s3i1) ,.o1(incr32s3ot) );	// line#=../rle.cpp:74
jpeg_incr8u INST_incr8u_1 ( .i1(incr8u1i1) ,.o1(incr8u1ot) );	// line#=../rle.cpp:68,73,79
jpeg_incr8u INST_incr8u_2 ( .i1(incr8u2i1) ,.o1(incr8u2ot) );	// line#=../rle.cpp:69,74,80,111,142
jpeg_incr4s INST_incr4s_1 ( .i1(incr4s1i1) ,.o1(incr4s1ot) );	// line#=../rle.cpp:34
jpeg_lop8u_1 INST_lop8u_1_1 ( .i1(lop8u_11i1) ,.i2(lop8u_11i2) ,.o1(lop8u_11ot) );	// line#=../rle.cpp:109,110
assign	lop8u_11ot_port = lop8u_11ot ;
jpeg_sub12s_9 INST_sub12s_9_1 ( .i1(sub12s_91i1) ,.i2(sub12s_91i2) ,.o1(sub12s_91ot) );	// line#=../rle.cpp:52
jpeg_sub8u INST_sub8u_1 ( .i1(sub8u1i1) ,.i2(sub8u1i2) ,.o1(sub8u1ot) );	// line#=../rle.cpp:77,78,83,84,86
assign	jpeg_out_a00 = jpeg_out_a00_r ;	// line#=../rle.h:60
assign	jpeg_out_a01 = jpeg_out_a01_r ;	// line#=../rle.h:60
assign	jpeg_out_a02 = jpeg_out_a02_r ;	// line#=../rle.h:60
assign	jpeg_out_a03 = jpeg_out_a03_r ;	// line#=../rle.h:60
assign	jpeg_out_a04 = jpeg_out_a04_r ;	// line#=../rle.h:60
assign	jpeg_out_a05 = jpeg_out_a05_r ;	// line#=../rle.h:60
assign	jpeg_out_a06 = jpeg_out_a06_r ;	// line#=../rle.h:60
assign	jpeg_out_a07 = jpeg_out_a07_r ;	// line#=../rle.h:60
assign	jpeg_out_a08 = jpeg_out_a08_r ;	// line#=../rle.h:60
assign	jpeg_out_a09 = jpeg_out_a09_r ;	// line#=../rle.h:60
assign	jpeg_out_a10 = jpeg_out_a10_r ;	// line#=../rle.h:60
assign	jpeg_out_a11 = jpeg_out_a11_r ;	// line#=../rle.h:60
assign	jpeg_out_a12 = jpeg_out_a12_r ;	// line#=../rle.h:60
assign	jpeg_out_a13 = jpeg_out_a13_r ;	// line#=../rle.h:60
assign	jpeg_out_a14 = jpeg_out_a14_r ;	// line#=../rle.h:60
assign	jpeg_out_a15 = jpeg_out_a15_r ;	// line#=../rle.h:60
assign	jpeg_out_a16 = jpeg_out_a16_r ;	// line#=../rle.h:60
assign	jpeg_out_a17 = jpeg_out_a17_r ;	// line#=../rle.h:60
assign	jpeg_out_a18 = jpeg_out_a18_r ;	// line#=../rle.h:60
assign	jpeg_out_a19 = jpeg_out_a19_r ;	// line#=../rle.h:60
assign	jpeg_out_a20 = jpeg_out_a20_r ;	// line#=../rle.h:60
assign	jpeg_out_a21 = jpeg_out_a21_r ;	// line#=../rle.h:60
assign	jpeg_out_a22 = jpeg_out_a22_r ;	// line#=../rle.h:60
assign	jpeg_out_a23 = jpeg_out_a23_r ;	// line#=../rle.h:60
assign	jpeg_out_a24 = jpeg_out_a24_r ;	// line#=../rle.h:60
assign	jpeg_out_a25 = jpeg_out_a25_r ;	// line#=../rle.h:60
assign	jpeg_out_a26 = jpeg_out_a26_r ;	// line#=../rle.h:60
assign	jpeg_out_a27 = jpeg_out_a27_r ;	// line#=../rle.h:60
assign	jpeg_out_a28 = jpeg_out_a28_r ;	// line#=../rle.h:60
assign	jpeg_out_a29 = jpeg_out_a29_r ;	// line#=../rle.h:60
assign	jpeg_out_a30 = jpeg_out_a30_r ;	// line#=../rle.h:60
assign	jpeg_out_a31 = jpeg_out_a31_r ;	// line#=../rle.h:60
assign	jpeg_out_a32 = jpeg_out_a32_r ;	// line#=../rle.h:60
assign	jpeg_out_a33 = jpeg_out_a33_r ;	// line#=../rle.h:60
assign	jpeg_out_a34 = jpeg_out_a34_r ;	// line#=../rle.h:60
assign	jpeg_out_a35 = jpeg_out_a35_r ;	// line#=../rle.h:60
assign	jpeg_out_a36 = jpeg_out_a36_r ;	// line#=../rle.h:60
assign	jpeg_out_a37 = jpeg_out_a37_r ;	// line#=../rle.h:60
assign	jpeg_out_a38 = jpeg_out_a38_r ;	// line#=../rle.h:60
assign	jpeg_out_a39 = jpeg_out_a39_r ;	// line#=../rle.h:60
assign	jpeg_out_a40 = jpeg_out_a40_r ;	// line#=../rle.h:60
assign	jpeg_out_a41 = jpeg_out_a41_r ;	// line#=../rle.h:60
assign	jpeg_out_a42 = jpeg_out_a42_r ;	// line#=../rle.h:60
assign	jpeg_out_a43 = jpeg_out_a43_r ;	// line#=../rle.h:60
assign	jpeg_out_a44 = jpeg_out_a44_r ;	// line#=../rle.h:60
assign	jpeg_out_a45 = jpeg_out_a45_r ;	// line#=../rle.h:60
assign	jpeg_out_a46 = jpeg_out_a46_r ;	// line#=../rle.h:60
assign	jpeg_out_a47 = jpeg_out_a47_r ;	// line#=../rle.h:60
assign	jpeg_out_a48 = jpeg_out_a48_r ;	// line#=../rle.h:60
assign	jpeg_out_a49 = jpeg_out_a49_r ;	// line#=../rle.h:60
assign	jpeg_out_a50 = jpeg_out_a50_r ;	// line#=../rle.h:60
assign	jpeg_out_a51 = jpeg_out_a51_r ;	// line#=../rle.h:60
assign	jpeg_out_a52 = jpeg_out_a52_r ;	// line#=../rle.h:60
assign	jpeg_out_a53 = jpeg_out_a53_r ;	// line#=../rle.h:60
assign	jpeg_out_a54 = jpeg_out_a54_r ;	// line#=../rle.h:60
assign	jpeg_out_a55 = jpeg_out_a55_r ;	// line#=../rle.h:60
assign	jpeg_out_a56 = jpeg_out_a56_r ;	// line#=../rle.h:60
assign	jpeg_out_a57 = jpeg_out_a57_r ;	// line#=../rle.h:60
assign	jpeg_out_a58 = jpeg_out_a58_r ;	// line#=../rle.h:60
assign	jpeg_out_a59 = jpeg_out_a59_r ;	// line#=../rle.h:60
assign	jpeg_out_a60 = jpeg_out_a60_r ;	// line#=../rle.h:60
assign	jpeg_out_a61 = jpeg_out_a61_r ;	// line#=../rle.h:60
assign	jpeg_out_a62 = jpeg_out_a62_r ;	// line#=../rle.h:60
assign	jpeg_out_a63 = jpeg_out_a63_r ;	// line#=../rle.h:60
assign	jpeg_out_a64 = jpeg_out_a64_r ;	// line#=../rle.h:60
assign	jpeg_out_a65 = jpeg_out_a65_r ;	// line#=../rle.h:60
assign	jpeg_out_a66 = jpeg_out_a66_r ;	// line#=../rle.h:60
assign	jpeg_out_a67 = jpeg_out_a67_r ;	// line#=../rle.h:60
assign	jpeg_out_a68 = jpeg_out_a68_r ;	// line#=../rle.h:60
assign	jpeg_out_a69 = jpeg_out_a69_r ;	// line#=../rle.h:60
assign	jpeg_out_a70 = jpeg_out_a70_r ;	// line#=../rle.h:60
assign	jpeg_out_a71 = jpeg_out_a71_r ;	// line#=../rle.h:60
assign	jpeg_out_a72 = jpeg_out_a72_r ;	// line#=../rle.h:60
assign	jpeg_out_a73 = jpeg_out_a73_r ;	// line#=../rle.h:60
assign	jpeg_out_a74 = jpeg_out_a74_r ;	// line#=../rle.h:60
assign	jpeg_out_a75 = jpeg_out_a75_r ;	// line#=../rle.h:60
assign	jpeg_out_a76 = jpeg_out_a76_r ;	// line#=../rle.h:60
assign	jpeg_out_a77 = jpeg_out_a77_r ;	// line#=../rle.h:60
assign	jpeg_out_a78 = jpeg_out_a78_r ;	// line#=../rle.h:60
assign	jpeg_out_a79 = jpeg_out_a79_r ;	// line#=../rle.h:60
assign	jpeg_out_a80 = jpeg_out_a80_r ;	// line#=../rle.h:60
assign	jpeg_out_a81 = jpeg_out_a81_r ;	// line#=../rle.h:60
assign	jpeg_out_a82 = jpeg_out_a82_r ;	// line#=../rle.h:60
assign	jpeg_out_a83 = jpeg_out_a83_r ;	// line#=../rle.h:60
assign	jpeg_out_a84 = jpeg_out_a84_r ;	// line#=../rle.h:60
assign	jpeg_out_a85 = jpeg_out_a85_r ;	// line#=../rle.h:60
assign	jpeg_out_a86 = jpeg_out_a86_r ;	// line#=../rle.h:60
assign	jpeg_out_a87 = jpeg_out_a87_r ;	// line#=../rle.h:60
assign	jpeg_out_a88 = jpeg_out_a88_r ;	// line#=../rle.h:60
assign	jpeg_out_a89 = jpeg_out_a89_r ;	// line#=../rle.h:60
assign	jpeg_out_a90 = jpeg_out_a90_r ;	// line#=../rle.h:60
assign	jpeg_out_a91 = jpeg_out_a91_r ;	// line#=../rle.h:60
assign	jpeg_out_a92 = jpeg_out_a92_r ;	// line#=../rle.h:60
assign	jpeg_out_a93 = jpeg_out_a93_r ;	// line#=../rle.h:60
assign	jpeg_out_a94 = jpeg_out_a94_r ;	// line#=../rle.h:60
assign	jpeg_out_a95 = jpeg_out_a95_r ;	// line#=../rle.h:60
assign	jpeg_out_a96 = jpeg_out_a96_r ;	// line#=../rle.h:60
assign	jpeg_out_a97 = jpeg_out_a97_r ;	// line#=../rle.h:60
assign	jpeg_out_a98 = jpeg_out_a98_r ;	// line#=../rle.h:60
assign	jpeg_out_a99 = jpeg_out_a99_r ;	// line#=../rle.h:60
assign	jpeg_out_a100 = jpeg_out_a100_r ;	// line#=../rle.h:60
assign	jpeg_out_a101 = jpeg_out_a101_r ;	// line#=../rle.h:60
assign	jpeg_out_a102 = jpeg_out_a102_r ;	// line#=../rle.h:60
assign	jpeg_out_a103 = jpeg_out_a103_r ;	// line#=../rle.h:60
assign	jpeg_out_a104 = jpeg_out_a104_r ;	// line#=../rle.h:60
assign	jpeg_out_a105 = jpeg_out_a105_r ;	// line#=../rle.h:60
assign	jpeg_out_a106 = jpeg_out_a106_r ;	// line#=../rle.h:60
assign	jpeg_out_a107 = jpeg_out_a107_r ;	// line#=../rle.h:60
assign	jpeg_out_a108 = jpeg_out_a108_r ;	// line#=../rle.h:60
assign	jpeg_out_a109 = jpeg_out_a109_r ;	// line#=../rle.h:60
assign	jpeg_out_a110 = jpeg_out_a110_r ;	// line#=../rle.h:60
assign	jpeg_out_a111 = jpeg_out_a111_r ;	// line#=../rle.h:60
assign	jpeg_out_a112 = jpeg_out_a112_r ;	// line#=../rle.h:60
assign	jpeg_out_a113 = jpeg_out_a113_r ;	// line#=../rle.h:60
assign	jpeg_out_a114 = jpeg_out_a114_r ;	// line#=../rle.h:60
assign	jpeg_out_a115 = jpeg_out_a115_r ;	// line#=../rle.h:60
assign	jpeg_out_a116 = jpeg_out_a116_r ;	// line#=../rle.h:60
assign	jpeg_out_a117 = jpeg_out_a117_r ;	// line#=../rle.h:60
assign	jpeg_out_a118 = jpeg_out_a118_r ;	// line#=../rle.h:60
assign	jpeg_out_a119 = jpeg_out_a119_r ;	// line#=../rle.h:60
assign	jpeg_out_a120 = jpeg_out_a120_r ;	// line#=../rle.h:60
assign	jpeg_out_a121 = jpeg_out_a121_r ;	// line#=../rle.h:60
assign	jpeg_out_a122 = jpeg_out_a122_r ;	// line#=../rle.h:60
assign	jpeg_out_a123 = jpeg_out_a123_r ;	// line#=../rle.h:60
assign	jpeg_out_a124 = jpeg_out_a124_r ;	// line#=../rle.h:60
assign	jpeg_out_a125 = jpeg_out_a125_r ;	// line#=../rle.h:60
assign	jpeg_out_a126 = jpeg_out_a126_r ;	// line#=../rle.h:60
assign	jpeg_out_a127 = jpeg_out_a127_r ;	// line#=../rle.h:60
assign	jpeg_len_out = jpeg_len_out_r ;	// line#=../rle.h:61
assign	valid = valid_r ;	// line#=../rle.h:62
always @ ( posedge clk )
	RG_len_02 <= RG_len_01 ;
always @ ( posedge clk )	// line#=../rle.cpp:83,84
	RG_75_02 <= RG_80_01 ;
always @ ( posedge clk )
	RG_len_01 <= RG_len_01_1 ;
always @ ( posedge clk )
	RG_i_01 <= RG_i_j_01 ;
always @ ( posedge clk )	// line#=../rle.cpp:61,62
	RG_k_01 <= RG_i_k_01 ;
assign	CT_12 = ( ( ~|RG_i_j_01 ) & M_110 ) ;	// line#=../rle.cpp:117,118
assign	M_110 = ~|{ ( RG_i_k_01 [31] & RG_i_k_01 [0] ) , ~RG_i_k_01 [0] } ;	// line#=../rle.cpp:117,118,148,149
assign	CT_26 = ( ( ~|{ RG_i_j_01 [31:3] , ~RG_i_j_01 [2:0] } ) & M_110 ) ;	// line#=../rle.cpp:148,149
always @ ( M_134 or RG_quantized_block_rl_02 )	// line#=../rle.cpp:77,78
	case ( ~|RG_quantized_block_rl_02 )
	1'h1 :
		M_02_t1 = M_134 ;	// line#=../rle.cpp:77,78
	1'h0 :
		M_02_t1 = 1'h0 ;	// line#=../rle.cpp:77,78
	default :
		M_02_t1 = 1'hx ;
	endcase
assign	CT_31 = ( RG_i_j_01 [31] | ( ~|RG_i_j_01 [30:6] ) ) ;	// line#=../rle.cpp:57,58,61,62
assign	CT_31_port = CT_31 ;
always @ ( zz_RD1 or RG_82_01 )	// line#=../rle.cpp:61,62
	case ( RG_82_01 )
	1'h1 :
		M_01_t1 = ~|zz_RD1 ;	// line#=../rle.cpp:61,62
	1'h0 :
		M_01_t1 = 1'h0 ;	// line#=../rle.cpp:61,62
	default :
		M_01_t1 = 1'hx ;
	endcase
assign	M_134 = ~|RG_quantized_block_rl_02_1 ;	// line#=../rle.cpp:77,78,83,84
always @ ( M_134 or RG_quantized_block_rl_02 )	// line#=../rle.cpp:83,84
	case ( ~|{ RG_quantized_block_rl_02 [8:4] , ~RG_quantized_block_rl_02 [3:0] } )
	1'h1 :
		M_03_t1 = M_134 ;	// line#=../rle.cpp:83,84
	1'h0 :
		M_03_t1 = 1'h0 ;	// line#=../rle.cpp:83,84
	default :
		M_03_t1 = 1'hx ;
	endcase
assign	CT_35 = ~|{ RG_i_02 [31:7] , ~RG_i_02 [6] , RG_i_02 [5:0] } ;	// line#=../rle.cpp:66,67
assign	FL01_01_Leos_all = ( FL01_01_eos & FL01_02_eos ) ;
always @ ( FL01_01_streg )
	case ( FL01_01_streg )
	1'h0 :
		FL01_01_next = 1'h0 ;
	1'h1 :
		FL01_01_next = 1'h1 ;
	default :
		FL01_01_next = 1'hx ;
	endcase
assign	FL02_01_Leos_all = ( ( FL02_01_eos & FL02_02_eos ) & FL02_03_eos ) ;
always @ ( FL02_01_streg )
	case ( FL02_01_streg )
	1'h0 :
		FL02_01_next = 1'h0 ;
	1'h1 :
		FL02_01_next = 1'h1 ;
	default :
		FL02_01_next = 1'hx ;
	endcase
jpeg_MEMB9W64 zz ( .RA1(zz_RA1) ,.RD1(zz_RD1) ,.RCLK1(clk) ,.WA2(zz_WA2) ,.WD2(zz_WD2) ,
	.WE2(zz_WE2) ,.WCLK2(clk) );	// line#=../rle.h:65
assign	sub12s_91i1 = zz_RD1 ;	// line#=../rle.cpp:52,53
assign	sub12s_91i2 = RG_previous_dc ;	// line#=../rle.cpp:52
assign	lop8u_11i1 = RG_k ;	// line#=../rle.cpp:109,110
assign	lop8u_11i2 = 6'h24 ;	// line#=../rle.cpp:109,110
assign	incr4s1i1 = RG_j_03 ;	// line#=../rle.cpp:34
assign	incr32s3i1 = RG_i_02 ;	// line#=../rle.cpp:74
assign	decr8u_71i1 = RG_len_01_1 [6:0] ;	// line#=../rle.cpp:77,78
assign	sub8u_71i1 = RG_len_01_1 [6:0] ;	// line#=../rle.cpp:83,84
assign	sub8u_71i2 = 3'h4 ;	// line#=../rle.cpp:83,84
assign	sub8u_7_11i1 = RG_len_01_1 [6:0] ;	// line#=../rle.cpp:83,84
assign	sub8u_7_11i2 = 2'h3 ;	// line#=../rle.cpp:83,84
assign	U_05 = ( ST1_03d & lop8u_11ot ) ;	// line#=../rle.cpp:109,110
assign	U_06 = ( ST1_03d & ( ~lop8u_11ot ) ) ;	// line#=../rle.cpp:109,110
assign	U_07 = ( U_05 & M_116 ) ;	// line#=../rle.cpp:111
assign	U_08 = ( U_05 & M_112 ) ;	// line#=../rle.cpp:111
assign	U_09 = ( U_05 & M_120 ) ;	// line#=../rle.cpp:111
assign	U_10 = ( U_05 & M_127 ) ;	// line#=../rle.cpp:111
assign	U_11 = ( U_05 & M_125 ) ;	// line#=../rle.cpp:111
assign	U_12 = ( U_05 & M_129 ) ;	// line#=../rle.cpp:111
assign	U_13 = ( U_05 & M_131 ) ;	// line#=../rle.cpp:111
assign	U_14 = ( U_05 & M_123 ) ;	// line#=../rle.cpp:111
assign	C_02 = ( ( ~|RG_i_k_01 ) & M_133 ) ;	// line#=../rle.cpp:112,113
assign	U_79 = ( U_05 & C_02 ) ;	// line#=../rle.cpp:112,113
assign	U_80 = ( U_05 & ( ~C_02 ) ) ;	// line#=../rle.cpp:112,113
assign	U_81 = ( U_80 & CT_12 ) ;	// line#=../rle.cpp:117,118
assign	U_82 = ( U_80 & ( ~CT_12 ) ) ;	// line#=../rle.cpp:117,118
assign	U_83 = ( U_82 & ( ~FF_d ) ) ;	// line#=../rle.cpp:122,123
assign	U_84 = ( U_82 & FF_d ) ;	// line#=../rle.cpp:122,123
assign	U_87 = ( ST1_04d & ( ~RG_k_01_1 [6] ) ) ;	// line#=../rle.cpp:140,141
assign	M_116 = ~|RG_i_k_01 [2:0] ;	// line#=../rle.cpp:111,142
assign	U_89 = ( U_87 & M_116 ) ;	// line#=../rle.cpp:142
assign	M_112 = ~|( RG_i_k_01 [2:0] ^ 3'h1 ) ;	// line#=../rle.cpp:111,142
assign	U_90 = ( U_87 & M_112 ) ;	// line#=../rle.cpp:142
assign	M_120 = ~|( RG_i_k_01 [2:0] ^ 3'h2 ) ;	// line#=../rle.cpp:111,142
assign	U_91 = ( U_87 & M_120 ) ;	// line#=../rle.cpp:142
assign	M_127 = ~|( RG_i_k_01 [2:0] ^ 3'h3 ) ;	// line#=../rle.cpp:111,142
assign	U_92 = ( U_87 & M_127 ) ;	// line#=../rle.cpp:142
assign	M_125 = ~|( RG_i_k_01 [2:0] ^ 3'h4 ) ;	// line#=../rle.cpp:111,142
assign	U_93 = ( U_87 & M_125 ) ;	// line#=../rle.cpp:142
assign	M_129 = ~|( RG_i_k_01 [2:0] ^ 3'h5 ) ;	// line#=../rle.cpp:111,142
assign	U_94 = ( U_87 & M_129 ) ;	// line#=../rle.cpp:142
assign	M_131 = ~|( RG_i_k_01 [2:0] ^ 3'h6 ) ;	// line#=../rle.cpp:111,142
assign	U_95 = ( U_87 & M_131 ) ;	// line#=../rle.cpp:142
assign	M_123 = ~|( RG_i_k_01 [2:0] ^ 3'h7 ) ;	// line#=../rle.cpp:111,142
assign	U_96 = ( U_87 & M_123 ) ;	// line#=../rle.cpp:142
assign	M_133 = ~|{ ( RG_i_j_01 [31] & RG_i_j_01 [0] ) , RG_i_j_01 [0] } ;	// line#=../rle.cpp:112,113,143,144
assign	C_04 = ( ( ~|{ RG_i_k_01 [31:3] , ~RG_i_k_01 [2:0] } ) & M_133 ) ;	// line#=../rle.cpp:143,144
assign	U_161 = ( U_87 & C_04 ) ;	// line#=../rle.cpp:143,144
assign	U_162 = ( U_87 & ( ~C_04 ) ) ;	// line#=../rle.cpp:143,144
assign	U_163 = ( U_162 & CT_26 ) ;	// line#=../rle.cpp:148,149
assign	U_164 = ( U_162 & ( ~CT_26 ) ) ;	// line#=../rle.cpp:148,149
assign	U_165 = ( U_164 & ( ~FF_d ) ) ;	// line#=../rle.cpp:153,154
assign	U_166 = ( U_164 & FF_d ) ;	// line#=../rle.cpp:153,154
assign	U_171 = ( ST1_06d & CT_31 ) ;	// line#=../rle.cpp:57,58
assign	U_173 = ( ST1_08d & ( ~M_02_t1 ) ) ;	// line#=../rle.cpp:77,78
assign	U_176 = ( ST1_08d & ( ~JF_05 ) ) ;
assign	U_177 = ( ST1_10d & FL01_01_01a ) ;
assign	U_180 = ( ST1_10d & FL01_02_01a ) ;
assign	U_188 = ( ST1_10d & ( ~FL01_02_streg ) ) ;
assign	U_189 = ( ST1_10d & FL01_02_streg ) ;
assign	U_193 = ( U_189 & ( ~FJ_11_15 ) ) ;
assign	U_196 = ( ST1_10d & FJ_11_15 ) ;
assign	U_198 = ( ST1_10d & FL01_02_break ) ;
assign	U_202 = ( ST1_11d & FL02_01_01a ) ;
assign	U_204 = ( ST1_11d & FL02_03_01a ) ;
assign	U_207 = ( U_204 & M_03_t1 ) ;	// line#=../rle.cpp:83,84
assign	U_212 = ( ST1_11d & ( ~FL02_02_streg ) ) ;
assign	U_213 = ( ST1_11d & FL02_02_streg ) ;
assign	U_218 = ( ST1_11d & ( ~FL02_03_streg ) ) ;
assign	U_219 = ( ST1_11d & FL02_03_streg ) ;
assign	U_223 = ( U_219 & ( ~FJ_14_17 ) ) ;
assign	U_228 = ( ST1_11d & FJ_14_17 ) ;
assign	U_230 = ( ST1_11d & FL02_03_break ) ;
assign	U_234 = ( ST1_12d & CT_35 ) ;	// line#=../rle.cpp:66,67
assign	U_235 = ( ST1_12d & ( ~CT_35 ) ) ;	// line#=../rle.cpp:66,67
assign	U_236 = ( ST1_13d & RG_82_01 ) ;	// line#=../rle.cpp:66,67
assign	U_237 = ( ST1_13d & ( ~RG_82_01 ) ) ;	// line#=../rle.cpp:66,67
assign	RG_previous_dc_en = ST1_56d ;
always @ ( posedge clk )
	if ( !rst )
		RG_previous_dc <= 9'h000 ;
	else if ( RG_previous_dc_en )
		RG_previous_dc <= RG_previous_dc_quantized_block ;
always @ ( FF_j or U_204 or incr4s1ot or ST1_02d or ST1_01d )
	RG_j_03_t = ( ( { 4{ ST1_01d } } & 4'hf /*-4'h1*/ )	// line#=../rle.cpp:34
		| ( { 4{ ST1_02d } } & incr4s1ot )		// line#=../rle.cpp:34
		| ( { 4{ U_204 } } & { 3'h0 , FF_j } )		// line#=../rle.cpp:83,84
		) ;
assign	RG_j_03_en = ( ST1_01d | ST1_02d | U_204 ) ;
always @ ( posedge clk )
	if ( RG_j_03_en )
		RG_j_03 <= RG_j_03_t ;	// line#=../rle.cpp:34,83,84
assign	M_136 = ( ST1_02d | ST1_06d ) ;
always @ ( U_06 )
	TR_01 = ( { 3{ U_06 } } & 3'h7 )	// line#=../rle.cpp:134
		 ;	// line#=../rle.cpp:59,105
always @ ( decr32s1ot or U_165 or U_83 or incr32s2ot or U_177 or U_166 or U_163 or 
	U_84 or U_81 or TR_01 or U_06 or M_136 )
	begin
	RG_i_k_01_t_c1 = ( M_136 | U_06 ) ;	// line#=../rle.cpp:59,105,134
	RG_i_k_01_t_c2 = ( ( ( ( U_81 | U_84 ) | U_163 ) | U_166 ) | U_177 ) ;	// line#=../rle.cpp:64,119,129,150,160
	RG_i_k_01_t_c3 = ( U_83 | U_165 ) ;	// line#=../rle.cpp:124,155
	RG_i_k_01_t = ( ( { 32{ RG_i_k_01_t_c1 } } & { 29'h00000000 , TR_01 } )	// line#=../rle.cpp:59,105,134
		| ( { 32{ RG_i_k_01_t_c2 } } & incr32s2ot )			// line#=../rle.cpp:64,119,129,150,160
		| ( { 32{ RG_i_k_01_t_c3 } } & decr32s1ot )			// line#=../rle.cpp:124,155
		) ;
	end
assign	RG_i_k_01_en = ( RG_i_k_01_t_c1 | RG_i_k_01_t_c2 | RG_i_k_01_t_c3 ) ;
always @ ( posedge clk )
	if ( RG_i_k_01_en )
		RG_i_k_01 <= RG_i_k_01_t ;	// line#=../rle.cpp:59,64,105,119,124,129
						// ,134,150,155,160
always @ ( FF_i or ST1_05d or U_06 )
	TR_02 = ( ( { 1{ U_06 } } & 1'h1 )	// line#=../rle.cpp:135
		| ( { 1{ ST1_05d } } & FF_i ) ) ;	// line#=../rle.cpp:105
always @ ( RG_i_02 or U_236 or incr32s3ot or U_237 or decr32s2ot or U_166 or U_84 or 
	incr32s1ot or U_177 or U_165 or U_161 or U_83 or U_79 or TR_02 or ST1_05d or 
	M_135 )
	begin
	RG_i_j_01_t_c1 = ( M_135 | ST1_05d ) ;	// line#=../rle.cpp:105,135
	RG_i_j_01_t_c2 = ( ( ( ( U_79 | U_83 ) | U_161 ) | U_165 ) | U_177 ) ;	// line#=../rle.cpp:61,62,63,114,125,145
										// ,156
	RG_i_j_01_t_c3 = ( U_84 | U_166 ) ;	// line#=../rle.cpp:130,161
	RG_i_j_01_t = ( ( { 32{ RG_i_j_01_t_c1 } } & { 31'h00000000 , TR_02 } )	// line#=../rle.cpp:105,135
		| ( { 32{ RG_i_j_01_t_c2 } } & incr32s1ot )			// line#=../rle.cpp:61,62,63,114,125,145
										// ,156
		| ( { 32{ RG_i_j_01_t_c3 } } & decr32s2ot )			// line#=../rle.cpp:130,161
		| ( { 32{ U_237 } } & incr32s3ot )				// line#=../rle.cpp:74
		| ( { 32{ U_236 } } & RG_i_02 ) ) ;
	end
assign	RG_i_j_01_en = ( RG_i_j_01_t_c1 | RG_i_j_01_t_c2 | RG_i_j_01_t_c3 | U_237 | 
	U_236 ) ;
always @ ( posedge clk )
	if ( RG_i_j_01_en )
		RG_i_j_01 <= RG_i_j_01_t ;	// line#=../rle.cpp:61,62,63,74,105,114
						// ,125,130,135,145,156,161
assign	RG_quantized_block_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_en )
		RG_quantized_block <= jpeg_in_a00 ;
assign	RG_quantized_block_1_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_1_en )
		RG_quantized_block_1 <= jpeg_in_a01 ;
assign	RG_quantized_block_2_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_2_en )
		RG_quantized_block_2 <= jpeg_in_a02 ;
assign	RG_quantized_block_3_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_3_en )
		RG_quantized_block_3 <= jpeg_in_a03 ;
assign	RG_quantized_block_4_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_4_en )
		RG_quantized_block_4 <= jpeg_in_a04 ;
assign	RG_quantized_block_5_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_5_en )
		RG_quantized_block_5 <= jpeg_in_a05 ;
assign	RG_quantized_block_6_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_6_en )
		RG_quantized_block_6 <= jpeg_in_a06 ;
assign	RG_quantized_block_7_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_7_en )
		RG_quantized_block_7 <= jpeg_in_a07 ;
assign	RG_quantized_block_8_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_8_en )
		RG_quantized_block_8 <= jpeg_in_a08 ;
assign	RG_quantized_block_9_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_9_en )
		RG_quantized_block_9 <= jpeg_in_a09 ;
assign	RG_quantized_block_10_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_10_en )
		RG_quantized_block_10 <= jpeg_in_a10 ;
assign	RG_quantized_block_11_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_11_en )
		RG_quantized_block_11 <= jpeg_in_a11 ;
assign	RG_quantized_block_12_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_12_en )
		RG_quantized_block_12 <= jpeg_in_a12 ;
assign	RG_quantized_block_13_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_13_en )
		RG_quantized_block_13 <= jpeg_in_a13 ;
assign	RG_quantized_block_14_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_14_en )
		RG_quantized_block_14 <= jpeg_in_a14 ;
assign	RG_quantized_block_15_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_15_en )
		RG_quantized_block_15 <= jpeg_in_a15 ;
assign	RG_quantized_block_16_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_16_en )
		RG_quantized_block_16 <= jpeg_in_a16 ;
assign	RG_quantized_block_17_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_17_en )
		RG_quantized_block_17 <= jpeg_in_a17 ;
assign	RG_quantized_block_18_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_18_en )
		RG_quantized_block_18 <= jpeg_in_a18 ;
assign	RG_quantized_block_19_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_19_en )
		RG_quantized_block_19 <= jpeg_in_a19 ;
assign	RG_quantized_block_20_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_20_en )
		RG_quantized_block_20 <= jpeg_in_a20 ;
assign	RG_quantized_block_21_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_21_en )
		RG_quantized_block_21 <= jpeg_in_a21 ;
assign	RG_quantized_block_22_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_22_en )
		RG_quantized_block_22 <= jpeg_in_a22 ;
assign	RG_quantized_block_23_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_23_en )
		RG_quantized_block_23 <= jpeg_in_a23 ;
assign	RG_quantized_block_24_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_24_en )
		RG_quantized_block_24 <= jpeg_in_a24 ;
assign	RG_quantized_block_25_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_25_en )
		RG_quantized_block_25 <= jpeg_in_a25 ;
assign	RG_quantized_block_26_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_26_en )
		RG_quantized_block_26 <= jpeg_in_a26 ;
assign	RG_quantized_block_27_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_27_en )
		RG_quantized_block_27 <= jpeg_in_a27 ;
assign	RG_quantized_block_28_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_28_en )
		RG_quantized_block_28 <= jpeg_in_a28 ;
assign	RG_quantized_block_29_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_29_en )
		RG_quantized_block_29 <= jpeg_in_a29 ;
assign	RG_quantized_block_30_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_30_en )
		RG_quantized_block_30 <= jpeg_in_a30 ;
assign	RG_quantized_block_31_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_31_en )
		RG_quantized_block_31 <= jpeg_in_a31 ;
assign	RG_quantized_block_32_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_32_en )
		RG_quantized_block_32 <= jpeg_in_a32 ;
assign	RG_quantized_block_33_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_33_en )
		RG_quantized_block_33 <= jpeg_in_a33 ;
assign	RG_quantized_block_34_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_34_en )
		RG_quantized_block_34 <= jpeg_in_a34 ;
assign	RG_quantized_block_35_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_35_en )
		RG_quantized_block_35 <= jpeg_in_a35 ;
assign	RG_quantized_block_36_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_36_en )
		RG_quantized_block_36 <= jpeg_in_a36 ;
assign	RG_quantized_block_37_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_37_en )
		RG_quantized_block_37 <= jpeg_in_a37 ;
assign	RG_quantized_block_38_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_38_en )
		RG_quantized_block_38 <= jpeg_in_a38 ;
assign	RG_quantized_block_39_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_39_en )
		RG_quantized_block_39 <= jpeg_in_a39 ;
assign	RG_quantized_block_40_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_40_en )
		RG_quantized_block_40 <= jpeg_in_a40 ;
assign	RG_quantized_block_41_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_41_en )
		RG_quantized_block_41 <= jpeg_in_a41 ;
assign	RG_quantized_block_42_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_42_en )
		RG_quantized_block_42 <= jpeg_in_a42 ;
assign	RG_quantized_block_43_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_43_en )
		RG_quantized_block_43 <= jpeg_in_a43 ;
assign	RG_quantized_block_44_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_44_en )
		RG_quantized_block_44 <= jpeg_in_a44 ;
assign	RG_quantized_block_45_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_45_en )
		RG_quantized_block_45 <= jpeg_in_a45 ;
assign	RG_quantized_block_46_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_46_en )
		RG_quantized_block_46 <= jpeg_in_a46 ;
assign	RG_quantized_block_47_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_47_en )
		RG_quantized_block_47 <= jpeg_in_a47 ;
assign	RG_quantized_block_48_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_48_en )
		RG_quantized_block_48 <= jpeg_in_a48 ;
assign	RG_quantized_block_49_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_49_en )
		RG_quantized_block_49 <= jpeg_in_a49 ;
assign	RG_quantized_block_50_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_50_en )
		RG_quantized_block_50 <= jpeg_in_a50 ;
assign	RG_quantized_block_51_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_51_en )
		RG_quantized_block_51 <= jpeg_in_a51 ;
assign	RG_quantized_block_52_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_52_en )
		RG_quantized_block_52 <= jpeg_in_a52 ;
assign	RG_quantized_block_53_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_53_en )
		RG_quantized_block_53 <= jpeg_in_a53 ;
assign	RG_quantized_block_54_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_54_en )
		RG_quantized_block_54 <= jpeg_in_a54 ;
assign	RG_quantized_block_55_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_55_en )
		RG_quantized_block_55 <= jpeg_in_a55 ;
assign	RG_quantized_block_56_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_56_en )
		RG_quantized_block_56 <= jpeg_in_a56 ;
assign	RG_quantized_block_57_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_57_en )
		RG_quantized_block_57 <= jpeg_in_a57 ;
assign	RG_quantized_block_58_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_58_en )
		RG_quantized_block_58 <= jpeg_in_a58 ;
assign	RG_quantized_block_59_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:45
	if ( RG_quantized_block_59_en )
		RG_quantized_block_59 <= jpeg_in_a59 ;
always @ ( RG_k_01 or U_180 or jpeg_in_a60 or ST1_02d )
	RG_k_quantized_block_02_t = ( ( { 9{ ST1_02d } } & jpeg_in_a60 )	// line#=../rle.cpp:45
		| ( { 9{ U_180 } } & RG_k_01 [8:0] ) ) ;
assign	RG_k_quantized_block_02_en = ( ST1_02d | U_180 ) ;
always @ ( posedge clk )
	if ( RG_k_quantized_block_02_en )
		RG_k_quantized_block_02 <= RG_k_quantized_block_02_t ;	// line#=../rle.cpp:45
jpeg_MEM_rl rl ( .AD1(rl_AD1) ,.RD1(rl_RD1) ,.WD1(rl_WD1) ,.WE1(rl_WE1) ,.CLK1(clk) ,
	.RA2(rl_RA2) ,.RD2(rl_RD2) ,.RA3(rl_RA3) ,.RD3(rl_RD3) );	// line#=../rle.cpp:23
always @ ( rl_RD3 or M_138 or jpeg_in_a61 or ST1_02d )
	RG_quantized_block_rl_02_t = ( ( { 9{ ST1_02d } } & jpeg_in_a61 )	// line#=../rle.cpp:45
		| ( { 9{ M_138 } } & rl_RD3 ) ) ;
assign	RG_quantized_block_rl_02_en = ( ST1_02d | M_138 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_02_en )
		RG_quantized_block_rl_02 <= RG_quantized_block_rl_02_t ;	// line#=../rle.cpp:45
assign	M_138 = ( ST1_07d | ( ST1_11d & FL02_02_01a ) ) ;
always @ ( rl_RD2 or M_138 or jpeg_in_a62 or ST1_02d )
	RG_quantized_block_rl_02_1_t = ( ( { 9{ ST1_02d } } & jpeg_in_a62 )	// line#=../rle.cpp:45
		| ( { 9{ M_138 } } & rl_RD2 )					// line#=../rle.cpp:77,78,83,84
		) ;
assign	RG_quantized_block_rl_02_1_en = ( ST1_02d | M_138 ) ;
always @ ( posedge clk )
	if ( RG_quantized_block_rl_02_1_en )
		RG_quantized_block_rl_02_1 <= RG_quantized_block_rl_02_1_t ;	// line#=../rle.cpp:45,77,78,83,84
always @ ( zz_RD1 or ST1_05d or jpeg_in_a63 or ST1_02d )
	RG_previous_dc_quantized_block_t = ( ( { 9{ ST1_02d } } & jpeg_in_a63 )	// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & zz_RD1 )					// line#=../rle.cpp:52,53
		) ;
assign	RG_previous_dc_quantized_block_en = ( ST1_02d | ST1_05d ) ;
always @ ( posedge clk )
	if ( RG_previous_dc_quantized_block_en )
		RG_previous_dc_quantized_block <= RG_previous_dc_quantized_block_t ;	// line#=../rle.cpp:45,52,53
always @ ( incr8u2ot or ST1_03d )
	RG_k_t = ( { 6{ ST1_03d } } & incr8u2ot [5:0] )	// line#=../rle.cpp:111
		 ;	// line#=../rle.cpp:105
always @ ( posedge clk )
	RG_k <= RG_k_t ;	// line#=../rle.cpp:105,111
assign	M_135 = ( ST1_02d | U_06 ) ;
always @ ( U_163 or U_79 or U_161 or U_81 or M_135 )
	begin
	FF_d_t_c1 = ( ( M_135 | U_81 ) | U_161 ) ;	// line#=../rle.cpp:105,120,136,146
	FF_d_t_c2 = ( U_79 | U_163 ) ;	// line#=../rle.cpp:115,151
	FF_d_t = ( { 1{ FF_d_t_c2 } } & 1'h1 )	// line#=../rle.cpp:115,151
		 ;	// line#=../rle.cpp:105,120,136,146
	end
assign	FF_d_en = ( FF_d_t_c1 | FF_d_t_c2 ) ;
always @ ( posedge clk )
	if ( FF_d_en )
		FF_d <= FF_d_t ;	// line#=../rle.cpp:105,115,120,136,146
					// ,151
assign	FF_j_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:36
	if ( FF_j_en )
		FF_j <= 1'h0 ;
assign	FF_i_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:37
	if ( FF_i_en )
		FF_i <= 1'h1 ;
always @ ( M_02_t1 or ST1_08d or ST1_02d )
	FF_len_t = ( ( { 1{ ST1_02d } } & 1'h1 )	// line#=../rle.cpp:39
		| ( { 1{ ST1_08d } } & ( ~M_02_t1 ) )	// line#=../rle.cpp:77,78
		) ;
assign	FF_len_en = ( ST1_02d | ST1_08d ) ;
always @ ( posedge clk )
	if ( FF_len_en )
		FF_len <= FF_len_t ;	// line#=../rle.cpp:39,77,78
assign	RG_len_03_en = U_204 ;
always @ ( posedge clk )
	if ( RG_len_03_en )
		RG_len_03 <= RG_len_02 ;
assign	RG_i_02_en = U_180 ;
always @ ( posedge clk )
	if ( RG_i_02_en )
		RG_i_02 <= RG_i_01 ;
always @ ( sub8u_71ot or U_202 or decr8u_71ot or ST1_06d )
	RG_80_01_t = ( ( { 7{ ST1_06d } } & decr8u_71ot )	// line#=../rle.cpp:77,78
		| ( { 7{ U_202 } } & sub8u_71ot )		// line#=../rle.cpp:83,84
		) ;
always @ ( posedge clk )
	RG_80_01 <= RG_80_01_t ;	// line#=../rle.cpp:77,78,83,84
always @ ( sub8u1ot or U_202 or incr8u2ot or M_139 or FF_len or ST1_05d )
	RG_len_01_1_t = ( ( { 8{ ST1_05d } } & { 7'h00 , FF_len } )
		| ( { 8{ M_139 } } & incr8u2ot )	// line#=../rle.cpp:69,74,80
		| ( { 8{ U_202 } } & sub8u1ot )		// line#=../rle.cpp:83,84,86
		) ;
assign	RG_len_01_1_en = ( ST1_05d | M_139 | U_202 ) ;
always @ ( posedge clk )
	if ( RG_len_01_1_en )
		RG_len_01_1 <= RG_len_01_1_t ;	// line#=../rle.cpp:69,74,80,83,84,86
always @ ( CT_35 or ST1_12d or U_177 or CT_31 or ST1_06d or RG_k_01_1 or ST1_04d )
	RG_82_01_t = ( ( { 1{ ST1_04d } } & ( ~RG_k_01_1 [6] ) )	// line#=../rle.cpp:140,141
		| ( { 1{ ST1_06d } } & CT_31 )				// line#=../rle.cpp:57,58
		| ( { 1{ U_177 } } & CT_31 )				// line#=../rle.cpp:61,62
		| ( { 1{ ST1_12d } } & CT_35 )				// line#=../rle.cpp:66,67
		) ;
assign	RG_82_01_en = ( ST1_04d | ST1_06d | U_177 | ST1_12d ) ;
always @ ( posedge clk )
	if ( RG_82_01_en )
		RG_82_01 <= RG_82_01_t ;	// line#=../rle.cpp:57,58,61,62,66,67,140
						// ,141
always @ ( sub8u_7_11ot or U_202 or sub8u1ot or ST1_06d or incr8u2ot or ST1_04d or 
	RG_k or ST1_03d )
	RG_k_01_1_t = ( ( { 7{ ST1_03d } } & { 1'h0 , RG_k } )
		| ( { 7{ ST1_04d } } & incr8u2ot [6:0] )	// line#=../rle.cpp:142
		| ( { 7{ ST1_06d } } & sub8u1ot [6:0] )		// line#=../rle.cpp:77,78
		| ( { 7{ U_202 } } & sub8u_7_11ot )		// line#=../rle.cpp:83,84
		) ;
always @ ( posedge clk )
	RG_k_01_1 <= RG_k_01_1_t ;	// line#=../rle.cpp:77,78,83,84,142
assign	JF_01 = ~( ~|{ ~incr4s1ot [3] , incr4s1ot [2:0] } ) ;	// line#=../rle.cpp:34,35
assign	JF_03 = ~RG_k_01_1 [6] ;
assign	JF_05 = ~M_02_t1 ;	// line#=../rle.cpp:77,78
assign	JF_05_port = JF_05 ;
assign	FL01_02_break = ( FL01_02_streg & FJ_11_15 ) ;
assign	M_171 = ( ST1_10d & FL01_01_streg ) ;
assign	FL01_01_01a = M_171 ;
assign	FL01_02_01a = U_189 ;
assign	FJ_11_15 = ( U_180 & ( ~( M_01_t1 & ( RG_k_01 [31] | ( ( ~|RG_k_01 [30:4] ) & ( 
	~&RG_k_01 [3:0] ) ) ) ) ) ) ;	// line#=../rle.cpp:61,62
assign	FL01_01_eos = ( ( ST1_10d & ( ~FL01_01_streg ) ) | U_196 ) ;
assign	FL01_02_eos = ( M_165 | U_198 ) ;
always @ ( U_171 or FL01_01_next or FJ_11_15 or ST1_10d )
	begin
	FL01_01_streg_t_c1 = ( ST1_10d & ( ~FJ_11_15 ) ) ;
	FL01_01_streg_t = ( ( { 1{ FL01_01_streg_t_c1 } } & FL01_01_next )
		| ( { 1{ U_171 } } & 1'h1 ) ) ;
	end
assign	FL01_01_streg_en = ( U_196 | FL01_01_streg_t_c1 | U_171 ) ;
always @ ( posedge clk )
	if ( FL01_01_streg_en )
		FL01_01_streg <= FL01_01_streg_t ;
assign	M_140 = ( ST1_10d & ( ~FL01_02_break ) ) ;
assign	M_165 = ( ( ( U_189 & FJ_11_15 ) | ( U_193 & ( ~FL01_01_ndat ) ) ) | ( U_188 & ( 
	~FL01_01_ndat ) ) ) ;
always @ ( U_188 or FL01_01_ndat or U_193 or M_165 or M_140 or U_171 or U_198 )
	begin
	FL01_02_streg_t_c1 = ( ( U_198 | U_171 ) | ( M_140 & M_165 ) ) ;
	FL01_02_streg_t_c2 = ( M_140 & ( ( U_193 & FL01_01_ndat ) | ( U_188 & FL01_01_ndat ) ) ) ;
	FL01_02_streg_t = ( { 1{ FL01_02_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_02_streg_en = ( FL01_02_streg_t_c1 | FL01_02_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_02_streg_en )
		FL01_02_streg <= FL01_02_streg_t ;
assign	FL01_01_ndat = M_171 ;
assign	FL02_03_break = ( FL02_03_streg & FJ_14_17 ) ;
assign	M_170 = ( ST1_11d & FL02_01_streg ) ;
assign	FL02_01_01a = M_170 ;
assign	FL02_02_01a = U_213 ;
assign	FL02_03_01a = U_219 ;
assign	FJ_14_17 = ( U_204 & ( ~M_03_t1 ) ) ;	// line#=../rle.cpp:83,84
assign	FL02_01_eos = ( ( ST1_11d & ( ~FL02_01_streg ) ) | U_228 ) ;
assign	FL02_02_eos = ( M_167 | U_228 ) ;
assign	FL02_03_eos = ( M_168 | U_230 ) ;
always @ ( ST1_09d or U_176 or FL02_01_next or M_141 )
	begin
	FL02_01_streg_t_c1 = ( U_176 | ST1_09d ) ;
	FL02_01_streg_t = ( ( { 1{ M_141 } } & FL02_01_next )
		| ( { 1{ FL02_01_streg_t_c1 } } & 1'h1 ) ) ;
	end
assign	FL02_01_streg_en = ( U_228 | M_141 | FL02_01_streg_t_c1 ) ;
always @ ( posedge clk )
	if ( FL02_01_streg_en )
		FL02_01_streg <= FL02_01_streg_t ;
assign	M_141 = ( ST1_11d & ( ~FJ_14_17 ) ) ;
assign	M_167 = ( ( U_213 & ( ~FL02_01_ndat ) ) | ( U_212 & ( ~FL02_01_ndat ) ) ) ;
always @ ( U_212 or FL02_01_ndat or U_213 or M_167 or M_141 or ST1_09d or U_176 or 
	U_228 )
	begin
	FL02_02_streg_t_c1 = ( ( ( U_228 | U_176 ) | ST1_09d ) | ( M_141 & M_167 ) ) ;
	FL02_02_streg_t_c2 = ( M_141 & ( ( U_213 & FL02_01_ndat ) | ( U_212 & FL02_01_ndat ) ) ) ;
	FL02_02_streg_t = ( { 1{ FL02_02_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL02_02_streg_en = ( FL02_02_streg_t_c1 | FL02_02_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL02_02_streg_en )
		FL02_02_streg <= FL02_02_streg_t ;
assign	M_142 = ( ST1_11d & ( ~FL02_03_break ) ) ;
assign	M_168 = ( ( ( U_219 & FJ_14_17 ) | ( U_223 & ( ~FL02_02_ndat ) ) ) | ( U_218 & ( 
	~FL02_02_ndat ) ) ) ;
always @ ( U_218 or FL02_02_ndat or U_223 or M_168 or M_142 or ST1_09d or U_176 or 
	U_230 )
	begin
	FL02_03_streg_t_c1 = ( ( ( U_230 | U_176 ) | ST1_09d ) | ( M_142 & M_168 ) ) ;
	FL02_03_streg_t_c2 = ( M_142 & ( ( U_223 & FL02_02_ndat ) | ( U_218 & FL02_02_ndat ) ) ) ;
	FL02_03_streg_t = ( { 1{ FL02_03_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL02_03_streg_en = ( FL02_03_streg_t_c1 | FL02_03_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL02_03_streg_en )
		FL02_03_streg <= FL02_03_streg_t ;
assign	FL02_01_ndat = M_170 ;
assign	FL02_02_ndat = U_213 ;
assign	jpeg_out_a00_r_en = ST1_14d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a00_r_en )
		jpeg_out_a00_r <= rl_RD1 ;
assign	jpeg_out_a01_r_en = ST1_14d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a01_r_en )
		jpeg_out_a01_r <= rl_RD3 ;
assign	jpeg_out_a02_r_en = ST1_14d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a02_r_en )
		jpeg_out_a02_r <= rl_RD2 ;
assign	jpeg_out_a03_r_en = ST1_15d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a03_r_en )
		jpeg_out_a03_r <= rl_RD3 ;
assign	jpeg_out_a04_r_en = ST1_15d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a04_r_en )
		jpeg_out_a04_r <= rl_RD2 ;
assign	jpeg_out_a05_r_en = ST1_15d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a05_r_en )
		jpeg_out_a05_r <= rl_RD1 ;
assign	jpeg_out_a06_r_en = ST1_16d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a06_r_en )
		jpeg_out_a06_r <= rl_RD3 ;
assign	jpeg_out_a07_r_en = ST1_16d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a07_r_en )
		jpeg_out_a07_r <= rl_RD2 ;
assign	jpeg_out_a08_r_en = ST1_16d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a08_r_en )
		jpeg_out_a08_r <= rl_RD1 ;
assign	jpeg_out_a09_r_en = ST1_17d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a09_r_en )
		jpeg_out_a09_r <= rl_RD3 ;
assign	jpeg_out_a10_r_en = ST1_17d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a10_r_en )
		jpeg_out_a10_r <= rl_RD2 ;
assign	jpeg_out_a11_r_en = ST1_17d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a11_r_en )
		jpeg_out_a11_r <= rl_RD1 ;
assign	jpeg_out_a12_r_en = ST1_18d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a12_r_en )
		jpeg_out_a12_r <= rl_RD3 ;
assign	jpeg_out_a13_r_en = ST1_18d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a13_r_en )
		jpeg_out_a13_r <= rl_RD2 ;
assign	jpeg_out_a14_r_en = ST1_18d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a14_r_en )
		jpeg_out_a14_r <= rl_RD1 ;
assign	jpeg_out_a15_r_en = ST1_19d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a15_r_en )
		jpeg_out_a15_r <= rl_RD3 ;
assign	jpeg_out_a16_r_en = ST1_19d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a16_r_en )
		jpeg_out_a16_r <= rl_RD2 ;
assign	jpeg_out_a17_r_en = ST1_19d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a17_r_en )
		jpeg_out_a17_r <= rl_RD1 ;
assign	jpeg_out_a18_r_en = ST1_20d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a18_r_en )
		jpeg_out_a18_r <= rl_RD3 ;
assign	jpeg_out_a19_r_en = ST1_20d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a19_r_en )
		jpeg_out_a19_r <= rl_RD2 ;
assign	jpeg_out_a20_r_en = ST1_20d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a20_r_en )
		jpeg_out_a20_r <= rl_RD1 ;
assign	jpeg_out_a21_r_en = ST1_21d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a21_r_en )
		jpeg_out_a21_r <= rl_RD3 ;
assign	jpeg_out_a22_r_en = ST1_21d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a22_r_en )
		jpeg_out_a22_r <= rl_RD2 ;
assign	jpeg_out_a23_r_en = ST1_21d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a23_r_en )
		jpeg_out_a23_r <= rl_RD1 ;
assign	jpeg_out_a24_r_en = ST1_22d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a24_r_en )
		jpeg_out_a24_r <= rl_RD3 ;
assign	jpeg_out_a25_r_en = ST1_22d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a25_r_en )
		jpeg_out_a25_r <= rl_RD2 ;
assign	jpeg_out_a26_r_en = ST1_22d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a26_r_en )
		jpeg_out_a26_r <= rl_RD1 ;
assign	jpeg_out_a27_r_en = ST1_23d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a27_r_en )
		jpeg_out_a27_r <= rl_RD3 ;
assign	jpeg_out_a28_r_en = ST1_23d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a28_r_en )
		jpeg_out_a28_r <= rl_RD2 ;
assign	jpeg_out_a29_r_en = ST1_23d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a29_r_en )
		jpeg_out_a29_r <= rl_RD1 ;
assign	jpeg_out_a30_r_en = ST1_24d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a30_r_en )
		jpeg_out_a30_r <= rl_RD3 ;
assign	jpeg_out_a31_r_en = ST1_24d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a31_r_en )
		jpeg_out_a31_r <= rl_RD2 ;
assign	jpeg_out_a32_r_en = ST1_24d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a32_r_en )
		jpeg_out_a32_r <= rl_RD1 ;
assign	jpeg_out_a33_r_en = ST1_25d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a33_r_en )
		jpeg_out_a33_r <= rl_RD3 ;
assign	jpeg_out_a34_r_en = ST1_25d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a34_r_en )
		jpeg_out_a34_r <= rl_RD2 ;
assign	jpeg_out_a35_r_en = ST1_25d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a35_r_en )
		jpeg_out_a35_r <= rl_RD1 ;
assign	jpeg_out_a36_r_en = ST1_26d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a36_r_en )
		jpeg_out_a36_r <= rl_RD3 ;
assign	jpeg_out_a37_r_en = ST1_26d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a37_r_en )
		jpeg_out_a37_r <= rl_RD2 ;
assign	jpeg_out_a38_r_en = ST1_26d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a38_r_en )
		jpeg_out_a38_r <= rl_RD1 ;
assign	jpeg_out_a39_r_en = ST1_27d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a39_r_en )
		jpeg_out_a39_r <= rl_RD3 ;
assign	jpeg_out_a40_r_en = ST1_27d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a40_r_en )
		jpeg_out_a40_r <= rl_RD2 ;
assign	jpeg_out_a41_r_en = ST1_27d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a41_r_en )
		jpeg_out_a41_r <= rl_RD1 ;
assign	jpeg_out_a42_r_en = ST1_28d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a42_r_en )
		jpeg_out_a42_r <= rl_RD3 ;
assign	jpeg_out_a43_r_en = ST1_28d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a43_r_en )
		jpeg_out_a43_r <= rl_RD2 ;
assign	jpeg_out_a44_r_en = ST1_28d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a44_r_en )
		jpeg_out_a44_r <= rl_RD1 ;
assign	jpeg_out_a45_r_en = ST1_29d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a45_r_en )
		jpeg_out_a45_r <= rl_RD3 ;
assign	jpeg_out_a46_r_en = ST1_29d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a46_r_en )
		jpeg_out_a46_r <= rl_RD2 ;
assign	jpeg_out_a47_r_en = ST1_29d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a47_r_en )
		jpeg_out_a47_r <= rl_RD1 ;
assign	jpeg_out_a48_r_en = ST1_30d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a48_r_en )
		jpeg_out_a48_r <= rl_RD3 ;
assign	jpeg_out_a49_r_en = ST1_30d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a49_r_en )
		jpeg_out_a49_r <= rl_RD2 ;
assign	jpeg_out_a50_r_en = ST1_30d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a50_r_en )
		jpeg_out_a50_r <= rl_RD1 ;
assign	jpeg_out_a51_r_en = ST1_31d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a51_r_en )
		jpeg_out_a51_r <= rl_RD3 ;
assign	jpeg_out_a52_r_en = ST1_31d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a52_r_en )
		jpeg_out_a52_r <= rl_RD2 ;
assign	jpeg_out_a53_r_en = ST1_31d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a53_r_en )
		jpeg_out_a53_r <= rl_RD1 ;
assign	jpeg_out_a54_r_en = ST1_32d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a54_r_en )
		jpeg_out_a54_r <= rl_RD3 ;
assign	jpeg_out_a55_r_en = ST1_32d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a55_r_en )
		jpeg_out_a55_r <= rl_RD2 ;
assign	jpeg_out_a56_r_en = ST1_32d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a56_r_en )
		jpeg_out_a56_r <= rl_RD1 ;
assign	jpeg_out_a57_r_en = ST1_33d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a57_r_en )
		jpeg_out_a57_r <= rl_RD3 ;
assign	jpeg_out_a58_r_en = ST1_33d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a58_r_en )
		jpeg_out_a58_r <= rl_RD2 ;
assign	jpeg_out_a59_r_en = ST1_33d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a59_r_en )
		jpeg_out_a59_r <= rl_RD1 ;
assign	jpeg_out_a60_r_en = ST1_34d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a60_r_en )
		jpeg_out_a60_r <= rl_RD3 ;
assign	jpeg_out_a61_r_en = ST1_34d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a61_r_en )
		jpeg_out_a61_r <= rl_RD2 ;
assign	jpeg_out_a62_r_en = ST1_34d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a62_r_en )
		jpeg_out_a62_r <= rl_RD1 ;
assign	jpeg_out_a63_r_en = ST1_35d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a63_r_en )
		jpeg_out_a63_r <= rl_RD2 ;
assign	jpeg_out_a64_r_en = ST1_35d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a64_r_en )
		jpeg_out_a64_r <= rl_RD3 ;
assign	jpeg_out_a65_r_en = ST1_35d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a65_r_en )
		jpeg_out_a65_r <= rl_RD1 ;
assign	jpeg_out_a66_r_en = ST1_36d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a66_r_en )
		jpeg_out_a66_r <= rl_RD2 ;
assign	jpeg_out_a67_r_en = ST1_36d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a67_r_en )
		jpeg_out_a67_r <= rl_RD3 ;
assign	jpeg_out_a68_r_en = ST1_36d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a68_r_en )
		jpeg_out_a68_r <= rl_RD1 ;
assign	jpeg_out_a69_r_en = ST1_37d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a69_r_en )
		jpeg_out_a69_r <= rl_RD2 ;
assign	jpeg_out_a70_r_en = ST1_37d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a70_r_en )
		jpeg_out_a70_r <= rl_RD3 ;
assign	jpeg_out_a71_r_en = ST1_37d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a71_r_en )
		jpeg_out_a71_r <= rl_RD1 ;
assign	jpeg_out_a72_r_en = ST1_38d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a72_r_en )
		jpeg_out_a72_r <= rl_RD2 ;
assign	jpeg_out_a73_r_en = ST1_38d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a73_r_en )
		jpeg_out_a73_r <= rl_RD3 ;
assign	jpeg_out_a74_r_en = ST1_38d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a74_r_en )
		jpeg_out_a74_r <= rl_RD1 ;
assign	jpeg_out_a75_r_en = ST1_39d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a75_r_en )
		jpeg_out_a75_r <= rl_RD2 ;
assign	jpeg_out_a76_r_en = ST1_39d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a76_r_en )
		jpeg_out_a76_r <= rl_RD3 ;
assign	jpeg_out_a77_r_en = ST1_39d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a77_r_en )
		jpeg_out_a77_r <= rl_RD1 ;
assign	jpeg_out_a78_r_en = ST1_40d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a78_r_en )
		jpeg_out_a78_r <= rl_RD2 ;
assign	jpeg_out_a79_r_en = ST1_40d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a79_r_en )
		jpeg_out_a79_r <= rl_RD3 ;
assign	jpeg_out_a80_r_en = ST1_40d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a80_r_en )
		jpeg_out_a80_r <= rl_RD1 ;
assign	jpeg_out_a81_r_en = ST1_41d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a81_r_en )
		jpeg_out_a81_r <= rl_RD2 ;
assign	jpeg_out_a82_r_en = ST1_41d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a82_r_en )
		jpeg_out_a82_r <= rl_RD3 ;
assign	jpeg_out_a83_r_en = ST1_41d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a83_r_en )
		jpeg_out_a83_r <= rl_RD1 ;
assign	jpeg_out_a84_r_en = ST1_42d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a84_r_en )
		jpeg_out_a84_r <= rl_RD2 ;
assign	jpeg_out_a85_r_en = ST1_42d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a85_r_en )
		jpeg_out_a85_r <= rl_RD3 ;
assign	jpeg_out_a86_r_en = ST1_42d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a86_r_en )
		jpeg_out_a86_r <= rl_RD1 ;
assign	jpeg_out_a87_r_en = ST1_43d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a87_r_en )
		jpeg_out_a87_r <= rl_RD2 ;
assign	jpeg_out_a88_r_en = ST1_43d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a88_r_en )
		jpeg_out_a88_r <= rl_RD3 ;
assign	jpeg_out_a89_r_en = ST1_43d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a89_r_en )
		jpeg_out_a89_r <= rl_RD1 ;
assign	jpeg_out_a90_r_en = ST1_44d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a90_r_en )
		jpeg_out_a90_r <= rl_RD2 ;
assign	jpeg_out_a91_r_en = ST1_44d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a91_r_en )
		jpeg_out_a91_r <= rl_RD3 ;
assign	jpeg_out_a92_r_en = ST1_44d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a92_r_en )
		jpeg_out_a92_r <= rl_RD1 ;
assign	jpeg_out_a93_r_en = ST1_45d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a93_r_en )
		jpeg_out_a93_r <= rl_RD2 ;
assign	jpeg_out_a94_r_en = ST1_45d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a94_r_en )
		jpeg_out_a94_r <= rl_RD3 ;
assign	jpeg_out_a95_r_en = ST1_45d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a95_r_en )
		jpeg_out_a95_r <= rl_RD1 ;
assign	jpeg_out_a96_r_en = ST1_46d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a96_r_en )
		jpeg_out_a96_r <= rl_RD2 ;
assign	jpeg_out_a97_r_en = ST1_46d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a97_r_en )
		jpeg_out_a97_r <= rl_RD3 ;
assign	jpeg_out_a98_r_en = ST1_46d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a98_r_en )
		jpeg_out_a98_r <= rl_RD1 ;
assign	jpeg_out_a99_r_en = ST1_47d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a99_r_en )
		jpeg_out_a99_r <= rl_RD2 ;
assign	jpeg_out_a100_r_en = ST1_47d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a100_r_en )
		jpeg_out_a100_r <= rl_RD3 ;
assign	jpeg_out_a101_r_en = ST1_47d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a101_r_en )
		jpeg_out_a101_r <= rl_RD1 ;
assign	jpeg_out_a102_r_en = ST1_48d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a102_r_en )
		jpeg_out_a102_r <= rl_RD2 ;
assign	jpeg_out_a103_r_en = ST1_48d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a103_r_en )
		jpeg_out_a103_r <= rl_RD3 ;
assign	jpeg_out_a104_r_en = ST1_48d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a104_r_en )
		jpeg_out_a104_r <= rl_RD1 ;
assign	jpeg_out_a105_r_en = ST1_49d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a105_r_en )
		jpeg_out_a105_r <= rl_RD2 ;
assign	jpeg_out_a106_r_en = ST1_49d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a106_r_en )
		jpeg_out_a106_r <= rl_RD3 ;
assign	jpeg_out_a107_r_en = ST1_49d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a107_r_en )
		jpeg_out_a107_r <= rl_RD1 ;
assign	jpeg_out_a108_r_en = ST1_50d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a108_r_en )
		jpeg_out_a108_r <= rl_RD2 ;
assign	jpeg_out_a109_r_en = ST1_50d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a109_r_en )
		jpeg_out_a109_r <= rl_RD3 ;
assign	jpeg_out_a110_r_en = ST1_50d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a110_r_en )
		jpeg_out_a110_r <= rl_RD1 ;
assign	jpeg_out_a111_r_en = ST1_51d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a111_r_en )
		jpeg_out_a111_r <= rl_RD2 ;
assign	jpeg_out_a112_r_en = ST1_51d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a112_r_en )
		jpeg_out_a112_r <= rl_RD3 ;
assign	jpeg_out_a113_r_en = ST1_51d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a113_r_en )
		jpeg_out_a113_r <= rl_RD1 ;
assign	jpeg_out_a114_r_en = ST1_52d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a114_r_en )
		jpeg_out_a114_r <= rl_RD2 ;
assign	jpeg_out_a115_r_en = ST1_52d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a115_r_en )
		jpeg_out_a115_r <= rl_RD3 ;
assign	jpeg_out_a116_r_en = ST1_52d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a116_r_en )
		jpeg_out_a116_r <= rl_RD1 ;
assign	jpeg_out_a117_r_en = ST1_53d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a117_r_en )
		jpeg_out_a117_r <= rl_RD2 ;
assign	jpeg_out_a118_r_en = ST1_53d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a118_r_en )
		jpeg_out_a118_r <= rl_RD3 ;
assign	jpeg_out_a119_r_en = ST1_53d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a119_r_en )
		jpeg_out_a119_r <= rl_RD1 ;
assign	jpeg_out_a120_r_en = ST1_54d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a120_r_en )
		jpeg_out_a120_r <= rl_RD2 ;
assign	jpeg_out_a121_r_en = ST1_54d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a121_r_en )
		jpeg_out_a121_r <= rl_RD3 ;
assign	jpeg_out_a122_r_en = ST1_54d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a122_r_en )
		jpeg_out_a122_r <= rl_RD1 ;
assign	jpeg_out_a123_r_en = ST1_55d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a123_r_en )
		jpeg_out_a123_r <= rl_RD2 ;
assign	jpeg_out_a124_r_en = ST1_55d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a124_r_en )
		jpeg_out_a124_r <= rl_RD3 ;
assign	jpeg_out_a125_r_en = ST1_55d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a125_r_en )
		jpeg_out_a125_r <= rl_RD1 ;
assign	jpeg_out_a126_r_en = ST1_56d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a126_r_en )
		jpeg_out_a126_r <= rl_RD1 ;
assign	jpeg_out_a127_r_en = ST1_56d ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a127_r_en )
		jpeg_out_a127_r <= rl_RD2 ;
assign	jpeg_len_out_r_en = ST1_14d ;
always @ ( posedge clk )	// line#=../rle.cpp:93
	if ( jpeg_len_out_r_en )
		jpeg_len_out_r <= { 4'h0 , RG_len_03 } ;
always @ ( ST1_56d )
	valid_r_t = ( { 1{ ST1_56d } } & 1'h1 )	// line#=../rle.cpp:95
		 ;	// line#=../rle.cpp:30
assign	valid_r_en = ( ST1_01d | ST1_56d ) ;
always @ ( posedge clk )
	if ( valid_r_en )
		valid_r <= valid_r_t ;	// line#=../rle.cpp:30,95
assign	sub8u1i1 = { ( U_202 & RG_len_01_1 [7] ) , RG_len_01_1 [6:0] } ;	// line#=../rle.cpp:77,78,83,84,86
assign	sub8u1i2 = 2'h2 ;	// line#=../rle.cpp:77,78,83,84,86
assign	incr8u1i1 = RG_len_01_1 ;	// line#=../rle.cpp:68,73,79
always @ ( RG_k_01_1 or U_87 or RG_k or U_05 )
	TR_04 = ( ( { 6{ U_05 } } & RG_k )		// line#=../rle.cpp:111
		| ( { 6{ U_87 } } & RG_k_01_1 [5:0] )	// line#=../rle.cpp:142
		) ;
always @ ( TR_04 or U_87 or U_05 or incr8u1ot or ST1_13d or ST1_09d )
	begin
	incr8u2i1_c1 = ( ST1_09d | ST1_13d ) ;	// line#=../rle.cpp:68,69,73,74,79,80
	incr8u2i1_c2 = ( U_05 | U_87 ) ;	// line#=../rle.cpp:111,142
	incr8u2i1 = ( ( { 8{ incr8u2i1_c1 } } & incr8u1ot )	// line#=../rle.cpp:68,69,73,74,79,80
		| ( { 8{ incr8u2i1_c2 } } & { 2'h0 , TR_04 } )	// line#=../rle.cpp:111,142
		) ;
	end
assign	incr32s1i1 = RG_i_j_01 ;	// line#=../rle.cpp:61,62,63,114,125,145
					// ,156
assign	incr32s2i1 = RG_i_k_01 ;	// line#=../rle.cpp:61,62,64,119,129,150
					// ,160
assign	decr32s1i1 = RG_i_k_01 ;	// line#=../rle.cpp:124,155
assign	decr32s2i1 = RG_i_j_01 ;	// line#=../rle.cpp:130,161
always @ ( RG_i_j_01 or CT_31 or U_177 or RG_i_02 or U_235 )	// line#=../rle.cpp:61,62,140,141
	begin
	zz_RA1_c1 = ( U_177 & CT_31 ) ;	// line#=../rle.cpp:61,62
	zz_RA1 = ( ( { 6{ U_235 } } & RG_i_02 [5:0] )		// line#=../rle.cpp:74
		| ( { 6{ zz_RA1_c1 } } & RG_i_j_01 [5:0] )	// line#=../rle.cpp:61,62
		) ;	// line#=../rle.cpp:52,53
	end
always @ ( RG_k_01_1 or U_89 or U_90 or U_91 or U_92 or U_93 or U_94 or U_95 or 
	U_96 or RG_k or U_07 or U_08 or U_09 or U_10 or U_11 or U_12 or U_13 or 
	U_14 )
	begin
	zz_WA2_c1 = ( ( ( ( ( ( ( U_14 | U_13 ) | U_12 ) | U_11 ) | U_10 ) | U_09 ) | 
		U_08 ) | U_07 ) ;	// line#=../rle.cpp:111
	zz_WA2_c2 = ( ( ( ( ( ( ( U_96 | U_95 ) | U_94 ) | U_93 ) | U_92 ) | U_91 ) | 
		U_90 ) | U_89 ) ;	// line#=../rle.cpp:142
	zz_WA2 = ( ( { 6{ zz_WA2_c1 } } & RG_k )		// line#=../rle.cpp:111
		| ( { 6{ zz_WA2_c2 } } & RG_k_01_1 [5:0] )	// line#=../rle.cpp:142
		) ;
	end
always @ ( RG_quantized_block_7 or RG_quantized_block_6 or RG_quantized_block_5 or 
	RG_quantized_block_4 or RG_quantized_block_3 or RG_quantized_block_2 or 
	RG_quantized_block_1 or RG_quantized_block or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_44 = RG_quantized_block ;	// line#=../rle.cpp:111
	3'h1 :
		TR_44 = RG_quantized_block_1 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_44 = RG_quantized_block_2 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_44 = RG_quantized_block_3 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_44 = RG_quantized_block_4 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_44 = RG_quantized_block_5 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_44 = RG_quantized_block_6 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_44 = RG_quantized_block_7 ;	// line#=../rle.cpp:111
	default :
		TR_44 = 9'hx ;
	endcase
always @ ( RG_quantized_block_15 or RG_quantized_block_14 or RG_quantized_block_13 or 
	RG_quantized_block_12 or RG_quantized_block_11 or RG_quantized_block_10 or 
	RG_quantized_block_9 or RG_quantized_block_8 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_45 = RG_quantized_block_8 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_45 = RG_quantized_block_9 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_45 = RG_quantized_block_10 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_45 = RG_quantized_block_11 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_45 = RG_quantized_block_12 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_45 = RG_quantized_block_13 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_45 = RG_quantized_block_14 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_45 = RG_quantized_block_15 ;	// line#=../rle.cpp:111
	default :
		TR_45 = 9'hx ;
	endcase
always @ ( RG_quantized_block_23 or RG_quantized_block_22 or RG_quantized_block_21 or 
	RG_quantized_block_20 or RG_quantized_block_19 or RG_quantized_block_18 or 
	RG_quantized_block_17 or RG_quantized_block_16 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_46 = RG_quantized_block_16 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_46 = RG_quantized_block_17 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_46 = RG_quantized_block_18 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_46 = RG_quantized_block_19 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_46 = RG_quantized_block_20 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_46 = RG_quantized_block_21 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_46 = RG_quantized_block_22 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_46 = RG_quantized_block_23 ;	// line#=../rle.cpp:111
	default :
		TR_46 = 9'hx ;
	endcase
always @ ( RG_quantized_block_31 or RG_quantized_block_30 or RG_quantized_block_29 or 
	RG_quantized_block_28 or RG_quantized_block_27 or RG_quantized_block_26 or 
	RG_quantized_block_25 or RG_quantized_block_24 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_47 = RG_quantized_block_24 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_47 = RG_quantized_block_25 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_47 = RG_quantized_block_26 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_47 = RG_quantized_block_27 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_47 = RG_quantized_block_28 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_47 = RG_quantized_block_29 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_47 = RG_quantized_block_30 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_47 = RG_quantized_block_31 ;	// line#=../rle.cpp:111
	default :
		TR_47 = 9'hx ;
	endcase
always @ ( RG_quantized_block_39 or RG_quantized_block_38 or RG_quantized_block_37 or 
	RG_quantized_block_36 or RG_quantized_block_35 or RG_quantized_block_34 or 
	RG_quantized_block_33 or RG_quantized_block_32 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_48 = RG_quantized_block_32 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_48 = RG_quantized_block_33 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_48 = RG_quantized_block_34 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_48 = RG_quantized_block_35 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_48 = RG_quantized_block_36 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_48 = RG_quantized_block_37 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_48 = RG_quantized_block_38 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_48 = RG_quantized_block_39 ;	// line#=../rle.cpp:111
	default :
		TR_48 = 9'hx ;
	endcase
always @ ( RG_quantized_block_47 or RG_quantized_block_46 or RG_quantized_block_45 or 
	RG_quantized_block_44 or RG_quantized_block_43 or RG_quantized_block_42 or 
	RG_quantized_block_41 or RG_quantized_block_40 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_49 = RG_quantized_block_40 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_49 = RG_quantized_block_41 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_49 = RG_quantized_block_42 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_49 = RG_quantized_block_43 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_49 = RG_quantized_block_44 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_49 = RG_quantized_block_45 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_49 = RG_quantized_block_46 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_49 = RG_quantized_block_47 ;	// line#=../rle.cpp:111
	default :
		TR_49 = 9'hx ;
	endcase
always @ ( RG_quantized_block_55 or RG_quantized_block_54 or RG_quantized_block_53 or 
	RG_quantized_block_52 or RG_quantized_block_51 or RG_quantized_block_50 or 
	RG_quantized_block_49 or RG_quantized_block_48 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_50 = RG_quantized_block_48 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_50 = RG_quantized_block_49 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_50 = RG_quantized_block_50 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_50 = RG_quantized_block_51 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_50 = RG_quantized_block_52 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_50 = RG_quantized_block_53 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_50 = RG_quantized_block_54 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_50 = RG_quantized_block_55 ;	// line#=../rle.cpp:111
	default :
		TR_50 = 9'hx ;
	endcase
always @ ( RG_previous_dc_quantized_block or RG_quantized_block_rl_02_1 or RG_quantized_block_rl_02 or 
	RG_k_quantized_block_02 or RG_quantized_block_59 or RG_quantized_block_58 or 
	RG_quantized_block_57 or RG_quantized_block_56 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_51 = RG_quantized_block_56 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_51 = RG_quantized_block_57 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_51 = RG_quantized_block_58 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_51 = RG_quantized_block_59 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_51 = RG_k_quantized_block_02 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_51 = RG_quantized_block_rl_02 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_51 = RG_quantized_block_rl_02_1 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_51 = RG_previous_dc_quantized_block ;	// line#=../rle.cpp:111
	default :
		TR_51 = 9'hx ;
	endcase
always @ ( U_96 or U_95 or U_94 or U_93 or U_92 or U_91 or U_90 or U_89 or TR_51 or 
	U_14 or TR_50 or U_13 or TR_49 or U_12 or TR_48 or U_11 or TR_47 or U_10 or 
	TR_46 or U_09 or TR_45 or U_08 or TR_44 or U_07 )
	zz_WD2 = ( ( { 9{ U_07 } } & TR_44 )	// line#=../rle.cpp:111
		| ( { 9{ U_08 } } & TR_45 )	// line#=../rle.cpp:111
		| ( { 9{ U_09 } } & TR_46 )	// line#=../rle.cpp:111
		| ( { 9{ U_10 } } & TR_47 )	// line#=../rle.cpp:111
		| ( { 9{ U_11 } } & TR_48 )	// line#=../rle.cpp:111
		| ( { 9{ U_12 } } & TR_49 )	// line#=../rle.cpp:111
		| ( { 9{ U_13 } } & TR_50 )	// line#=../rle.cpp:111
		| ( { 9{ U_14 } } & TR_51 )	// line#=../rle.cpp:111
		| ( { 9{ U_89 } } & TR_44 )	// line#=../rle.cpp:142
		| ( { 9{ U_90 } } & TR_45 )	// line#=../rle.cpp:142
		| ( { 9{ U_91 } } & TR_46 )	// line#=../rle.cpp:142
		| ( { 9{ U_92 } } & TR_47 )	// line#=../rle.cpp:142
		| ( { 9{ U_93 } } & TR_48 )	// line#=../rle.cpp:142
		| ( { 9{ U_94 } } & TR_49 )	// line#=../rle.cpp:142
		| ( { 9{ U_95 } } & TR_50 )	// line#=../rle.cpp:142
		| ( { 9{ U_96 } } & TR_51 )	// line#=../rle.cpp:142
		) ;
assign	M_113 = ~|( RG_i_j_01 [2:0] ^ 3'h1 ) ;	// line#=../rle.cpp:111,142
assign	M_117 = ~|RG_i_j_01 [2:0] ;	// line#=../rle.cpp:111,142
assign	M_122 = ~|( RG_i_j_01 [2:0] ^ 3'h2 ) ;	// line#=../rle.cpp:111,142
assign	M_124 = ~|( RG_i_j_01 [2:0] ^ 3'h7 ) ;	// line#=../rle.cpp:111,142
assign	M_126 = ~|( RG_i_j_01 [2:0] ^ 3'h4 ) ;	// line#=../rle.cpp:111,142
assign	M_128 = ~|( RG_i_j_01 [2:0] ^ 3'h3 ) ;	// line#=../rle.cpp:111,142
assign	M_130 = ~|( RG_i_j_01 [2:0] ^ 3'h5 ) ;	// line#=../rle.cpp:111,142
assign	M_132 = ~|( RG_i_j_01 [2:0] ^ 3'h6 ) ;	// line#=../rle.cpp:111,142
assign	zz_WE2 = ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( U_14 & M_124 ) | ( U_14 & M_132 ) ) | 
	( U_14 & M_130 ) ) | ( U_14 & M_126 ) ) | ( U_14 & M_128 ) ) | ( U_14 & M_122 ) ) | 
	( U_14 & M_113 ) ) | ( U_14 & M_117 ) ) | ( U_13 & M_124 ) ) | ( U_13 & M_132 ) ) | 
	( U_13 & M_130 ) ) | ( U_13 & M_126 ) ) | ( U_13 & M_128 ) ) | ( U_13 & M_122 ) ) | 
	( U_13 & M_113 ) ) | ( U_13 & M_117 ) ) | ( U_12 & M_124 ) ) | ( U_12 & M_132 ) ) | 
	( U_12 & M_130 ) ) | ( U_12 & M_126 ) ) | ( U_12 & M_128 ) ) | ( U_12 & M_122 ) ) | 
	( U_12 & M_113 ) ) | ( U_12 & M_117 ) ) | ( U_11 & M_124 ) ) | ( U_11 & M_132 ) ) | 
	( U_11 & M_130 ) ) | ( U_11 & M_126 ) ) | ( U_11 & M_128 ) ) | ( U_11 & M_122 ) ) | 
	( U_11 & M_113 ) ) | ( U_11 & M_117 ) ) | ( U_10 & M_124 ) ) | ( U_10 & M_132 ) ) | 
	( U_10 & M_130 ) ) | ( U_10 & M_126 ) ) | ( U_10 & M_128 ) ) | ( U_10 & M_122 ) ) | 
	( U_10 & M_113 ) ) | ( U_10 & M_117 ) ) | ( U_09 & M_124 ) ) | ( U_09 & M_132 ) ) | 
	( U_09 & M_130 ) ) | ( U_09 & M_126 ) ) | ( U_09 & M_128 ) ) | ( U_09 & M_122 ) ) | 
	( U_09 & M_113 ) ) | ( U_09 & M_117 ) ) | ( U_08 & M_124 ) ) | ( U_08 & M_132 ) ) | 
	( U_08 & M_130 ) ) | ( U_08 & M_126 ) ) | ( U_08 & M_128 ) ) | ( U_08 & M_122 ) ) | 
	( U_08 & M_113 ) ) | ( U_08 & M_117 ) ) | ( U_07 & M_124 ) ) | ( U_07 & M_132 ) ) | 
	( U_07 & M_130 ) ) | ( U_07 & M_126 ) ) | ( U_07 & M_128 ) ) | ( U_07 & M_122 ) ) | 
	( U_07 & M_113 ) ) | ( U_07 & M_117 ) ) | ( U_96 & M_124 ) ) | ( U_96 & M_132 ) ) | 
	( U_96 & M_130 ) ) | ( U_96 & M_126 ) ) | ( U_96 & M_128 ) ) | ( U_96 & M_122 ) ) | 
	( U_96 & M_113 ) ) | ( U_96 & M_117 ) ) | ( U_95 & M_124 ) ) | ( U_95 & M_132 ) ) | 
	( U_95 & M_130 ) ) | ( U_95 & M_126 ) ) | ( U_95 & M_128 ) ) | ( U_95 & M_122 ) ) | 
	( U_95 & M_113 ) ) | ( U_95 & M_117 ) ) | ( U_94 & M_124 ) ) | ( U_94 & M_132 ) ) | 
	( U_94 & M_130 ) ) | ( U_94 & M_126 ) ) | ( U_94 & M_128 ) ) | ( U_94 & M_122 ) ) | 
	( U_94 & M_113 ) ) | ( U_94 & M_117 ) ) | ( U_93 & M_124 ) ) | ( U_93 & M_132 ) ) | 
	( U_93 & M_130 ) ) | ( U_93 & M_126 ) ) | ( U_93 & M_128 ) ) | ( U_93 & M_122 ) ) | 
	( U_93 & M_113 ) ) | ( U_93 & M_117 ) ) | ( U_92 & M_124 ) ) | ( U_92 & M_132 ) ) | 
	( U_92 & M_130 ) ) | ( U_92 & M_126 ) ) | ( U_92 & M_128 ) ) | ( U_92 & M_122 ) ) | 
	( U_92 & M_113 ) ) | ( U_92 & M_117 ) ) | ( U_91 & M_124 ) ) | ( U_91 & M_132 ) ) | 
	( U_91 & M_130 ) ) | ( U_91 & M_126 ) ) | ( U_91 & M_128 ) ) | ( U_91 & M_122 ) ) | 
	( U_91 & M_113 ) ) | ( U_91 & M_117 ) ) | ( U_90 & M_124 ) ) | ( U_90 & M_132 ) ) | 
	( U_90 & M_130 ) ) | ( U_90 & M_126 ) ) | ( U_90 & M_128 ) ) | ( U_90 & M_122 ) ) | 
	( U_90 & M_113 ) ) | ( U_90 & M_117 ) ) | ( U_89 & M_124 ) ) | ( U_89 & M_132 ) ) | 
	( U_89 & M_130 ) ) | ( U_89 & M_126 ) ) | ( U_89 & M_128 ) ) | ( U_89 & M_122 ) ) | 
	( U_89 & M_113 ) ) | ( U_89 & M_117 ) ) ;
assign	M_137 = ( ST1_05d | ST1_14d ) ;
always @ ( ST1_15d )
	M_172 = ( { 2{ ST1_15d } } & 2'h3 )
		 ;	// line#=../rle.cpp:52
always @ ( ST1_17d )
	TR_17 = ( { 2{ ST1_17d } } & 2'h3 )
		 ;
assign	M_147 = ( ST1_16d | ST1_17d ) ;
always @ ( ST1_18d or TR_17 or M_147 )
	TR_18 = ( ( { 3{ M_147 } } & { 1'h0 , TR_17 } )
		| ( { 3{ ST1_18d } } & 3'h6 ) ) ;
assign	M_144 = ( M_137 | ST1_15d ) ;
always @ ( TR_18 or ST1_18d or M_147 or M_172 or M_144 )
	begin
	TR_06_c1 = ( M_147 | ST1_18d ) ;
	TR_06 = ( ( { 4{ M_144 } } & { 1'h0 , M_172 [1] , 1'h0 , M_172 [0] } )	// line#=../rle.cpp:52
		| ( { 4{ TR_06_c1 } } & { 1'h1 , TR_18 } ) ) ;
	end
always @ ( ST1_21d or ST1_20d or ST1_19d )
	TR_19 = ( ( { 3{ ST1_19d } } & 3'h1 )
		| ( { 3{ ST1_20d } } & 3'h4 )
		| ( { 3{ ST1_21d } } & 3'h7 ) ) ;
always @ ( ST1_23d or ST1_22d )
	TR_32 = ( ( { 3{ ST1_22d } } & 3'h2 )
		| ( { 3{ ST1_23d } } & 3'h5 ) ) ;
assign	M_149 = ( ( ST1_19d | ST1_20d ) | ST1_21d ) ;
always @ ( TR_32 or ST1_23d or ST1_22d or TR_19 or M_149 )
	begin
	TR_20_c1 = ( ST1_22d | ST1_23d ) ;
	TR_20 = ( ( { 4{ M_149 } } & { 1'h0 , TR_19 } )
		| ( { 4{ TR_20_c1 } } & { 1'h1 , TR_32 } ) ) ;
	end
assign	M_146 = ( ( ( M_144 | ST1_16d ) | ST1_17d ) | ST1_18d ) ;
always @ ( TR_20 or ST1_23d or ST1_22d or M_149 or TR_06 or M_146 )
	begin
	TR_07_c1 = ( ( M_149 | ST1_22d ) | ST1_23d ) ;
	TR_07 = ( ( { 5{ M_146 } } & { 1'h0 , TR_06 } )	// line#=../rle.cpp:52
		| ( { 5{ TR_07_c1 } } & { 1'h1 , TR_20 } ) ) ;
	end
always @ ( ST1_25d )
	TR_21 = ( { 2{ ST1_25d } } & 2'h3 )
		 ;
assign	M_150 = ( ST1_24d | ST1_25d ) ;
always @ ( ST1_26d or TR_21 or M_150 )
	TR_22 = ( ( { 3{ M_150 } } & { 1'h0 , TR_21 } )
		| ( { 3{ ST1_26d } } & 3'h6 ) ) ;
always @ ( ST1_29d or ST1_28d or ST1_27d )
	TR_33 = ( ( { 3{ ST1_27d } } & 3'h1 )
		| ( { 3{ ST1_28d } } & 3'h4 )
		| ( { 3{ ST1_29d } } & 3'h7 ) ) ;
assign	M_151 = ( M_150 | ST1_26d ) ;
always @ ( TR_33 or ST1_29d or ST1_28d or ST1_27d or TR_22 or M_151 )
	begin
	TR_23_c1 = ( ( ST1_27d | ST1_28d ) | ST1_29d ) ;
	TR_23 = ( ( { 4{ M_151 } } & { 1'h0 , TR_22 } )
		| ( { 4{ TR_23_c1 } } & { 1'h1 , TR_33 } ) ) ;
	end
always @ ( ST1_31d or ST1_30d )
	TR_34 = ( ( { 3{ ST1_30d } } & 3'h2 )
		| ( { 3{ ST1_31d } } & 3'h5 ) ) ;
always @ ( ST1_33d )
	TR_41 = ( { 2{ ST1_33d } } & 2'h3 )
		 ;
assign	M_154 = ( ST1_32d | ST1_33d ) ;
always @ ( ST1_34d or TR_41 or M_154 )
	TR_42 = ( ( { 3{ M_154 } } & { 1'h0 , TR_41 } )
		| ( { 3{ ST1_34d } } & 3'h6 ) ) ;
assign	M_153 = ( ST1_30d | ST1_31d ) ;
always @ ( TR_42 or ST1_34d or M_154 or TR_34 or M_153 )
	begin
	TR_35_c1 = ( M_154 | ST1_34d ) ;
	TR_35 = ( ( { 4{ M_153 } } & { 1'h0 , TR_34 } )
		| ( { 4{ TR_35_c1 } } & { 1'h1 , TR_42 } ) ) ;
	end
assign	M_152 = ( ( ( M_151 | ST1_27d ) | ST1_28d ) | ST1_29d ) ;
always @ ( TR_35 or ST1_34d or ST1_33d or ST1_32d or M_153 or TR_23 or M_152 )
	begin
	TR_24_c1 = ( ( ( M_153 | ST1_32d ) | ST1_33d ) | ST1_34d ) ;
	TR_24 = ( ( { 5{ M_152 } } & { 1'h0 , TR_23 } )
		| ( { 5{ TR_24_c1 } } & { 1'h1 , TR_35 } ) ) ;
	end
assign	M_148 = ( ( ( ( ( M_146 | ST1_19d ) | ST1_20d ) | ST1_21d ) | ST1_22d ) | 
	ST1_23d ) ;
always @ ( TR_24 or ST1_34d or ST1_33d or ST1_32d or ST1_31d or ST1_30d or M_152 or 
	TR_07 or M_148 )
	begin
	TR_08_c1 = ( ( ( ( ( M_152 | ST1_30d ) | ST1_31d ) | ST1_32d ) | ST1_33d ) | 
		ST1_34d ) ;
	TR_08 = ( ( { 6{ M_148 } } & { 1'h0 , TR_07 } )	// line#=../rle.cpp:52
		| ( { 6{ TR_08_c1 } } & { 1'h1 , TR_24 } ) ) ;
	end
always @ ( ST1_37d or ST1_36d or ST1_35d )
	TR_09 = ( ( { 3{ ST1_35d } } & 3'h1 )
		| ( { 3{ ST1_36d } } & 3'h4 )
		| ( { 3{ ST1_37d } } & 3'h7 ) ) ;
always @ ( ST1_39d or ST1_38d )
	TR_25 = ( ( { 3{ ST1_38d } } & 3'h2 )
		| ( { 3{ ST1_39d } } & 3'h5 ) ) ;
assign	M_155 = ( ( ST1_35d | ST1_36d ) | ST1_37d ) ;
always @ ( TR_25 or ST1_39d or ST1_38d or TR_09 or M_155 )
	begin
	TR_10_c1 = ( ST1_38d | ST1_39d ) ;
	TR_10 = ( ( { 4{ M_155 } } & { 1'h0 , TR_09 } )
		| ( { 4{ TR_10_c1 } } & { 1'h1 , TR_25 } ) ) ;
	end
always @ ( ST1_41d )
	TR_26 = ( { 2{ ST1_41d } } & 2'h3 )
		 ;
assign	M_158 = ( ST1_40d | ST1_41d ) ;
always @ ( ST1_42d or TR_26 or M_158 )
	TR_27 = ( ( { 3{ M_158 } } & { 1'h0 , TR_26 } )
		| ( { 3{ ST1_42d } } & 3'h6 ) ) ;
always @ ( ST1_45d or ST1_44d or ST1_43d )
	TR_36 = ( ( { 3{ ST1_43d } } & 3'h1 )
		| ( { 3{ ST1_44d } } & 3'h4 )
		| ( { 3{ ST1_45d } } & 3'h7 ) ) ;
assign	M_159 = ( M_158 | ST1_42d ) ;
always @ ( TR_36 or ST1_45d or ST1_44d or ST1_43d or TR_27 or M_159 )
	begin
	TR_28_c1 = ( ( ST1_43d | ST1_44d ) | ST1_45d ) ;
	TR_28 = ( ( { 4{ M_159 } } & { 1'h0 , TR_27 } )
		| ( { 4{ TR_28_c1 } } & { 1'h1 , TR_36 } ) ) ;
	end
assign	M_156 = ( ( M_155 | ST1_38d ) | ST1_39d ) ;
always @ ( TR_28 or ST1_45d or ST1_44d or ST1_43d or M_159 or TR_10 or M_156 )
	begin
	TR_11_c1 = ( ( ( M_159 | ST1_43d ) | ST1_44d ) | ST1_45d ) ;
	TR_11 = ( ( { 5{ M_156 } } & { 1'h0 , TR_10 } )
		| ( { 5{ TR_11_c1 } } & { 1'h1 , TR_28 } ) ) ;
	end
always @ ( ST1_47d or ST1_46d )
	TR_29 = ( ( { 3{ ST1_46d } } & 3'h2 )
		| ( { 3{ ST1_47d } } & 3'h5 ) ) ;
always @ ( ST1_49d )
	TR_37 = ( { 2{ ST1_49d } } & 2'h3 )
		 ;
assign	M_162 = ( ST1_48d | ST1_49d ) ;
always @ ( ST1_50d or TR_37 or M_162 )
	TR_38 = ( ( { 3{ M_162 } } & { 1'h0 , TR_37 } )
		| ( { 3{ ST1_50d } } & 3'h6 ) ) ;
assign	M_160 = ( ST1_46d | ST1_47d ) ;
always @ ( TR_38 or ST1_50d or M_162 or TR_29 or M_160 )
	begin
	TR_30_c1 = ( M_162 | ST1_50d ) ;
	TR_30 = ( ( { 4{ M_160 } } & { 1'h0 , TR_29 } )
		| ( { 4{ TR_30_c1 } } & { 1'h1 , TR_38 } ) ) ;
	end
always @ ( ST1_53d or ST1_52d or ST1_51d )
	TR_39 = ( ( { 3{ ST1_51d } } & 3'h1 )
		| ( { 3{ ST1_52d } } & 3'h4 )
		| ( { 3{ ST1_53d } } & 3'h7 ) ) ;
always @ ( ST1_56d or ST1_55d or ST1_54d )
	TR_43 = ( ( { 3{ ST1_54d } } & 3'h2 )
		| ( { 3{ ST1_55d } } & 3'h5 )
		| ( { 3{ ST1_56d } } & 3'h6 ) ) ;
assign	M_163 = ( ( ST1_51d | ST1_52d ) | ST1_53d ) ;
always @ ( TR_43 or ST1_56d or ST1_55d or ST1_54d or TR_39 or M_163 )
	begin
	TR_40_c1 = ( ( ST1_54d | ST1_55d ) | ST1_56d ) ;
	TR_40 = ( ( { 4{ M_163 } } & { 1'h0 , TR_39 } )
		| ( { 4{ TR_40_c1 } } & { 1'h1 , TR_43 } ) ) ;
	end
assign	M_161 = ( ( ( M_160 | ST1_48d ) | ST1_49d ) | ST1_50d ) ;
always @ ( TR_40 or ST1_56d or ST1_55d or ST1_54d or M_163 or TR_30 or M_161 )
	begin
	TR_31_c1 = ( ( ( M_163 | ST1_54d ) | ST1_55d ) | ST1_56d ) ;
	TR_31 = ( ( { 5{ M_161 } } & { 1'h0 , TR_30 } )
		| ( { 5{ TR_31_c1 } } & { 1'h1 , TR_40 } ) ) ;
	end
assign	M_157 = ( ( ( ( ( ( M_156 | ST1_40d ) | ST1_41d ) | ST1_42d ) | ST1_43d ) | 
	ST1_44d ) | ST1_45d ) ;
always @ ( TR_31 or ST1_56d or ST1_55d or ST1_54d or ST1_53d or ST1_52d or ST1_51d or 
	M_161 or TR_11 or M_157 )
	begin
	TR_12_c1 = ( ( ( ( ( ( M_161 | ST1_51d ) | ST1_52d ) | ST1_53d ) | ST1_54d ) | 
		ST1_55d ) | ST1_56d ) ;
	TR_12 = ( ( { 6{ M_157 } } & { 1'h0 , TR_11 } )
		| ( { 6{ TR_12_c1 } } & { 1'h1 , TR_31 } ) ) ;
	end
assign	M_139 = ( ST1_09d | ST1_13d ) ;
always @ ( TR_12 or ST1_56d or ST1_55d or ST1_54d or ST1_53d or ST1_52d or ST1_51d or 
	ST1_50d or ST1_49d or ST1_48d or ST1_47d or ST1_46d or M_157 or RG_75_02 or 
	U_207 or incr8u1ot or M_139 or RG_len_01_1 or ST1_12d or U_173 or TR_08 or 
	ST1_34d or ST1_33d or ST1_32d or ST1_31d or ST1_30d or ST1_29d or ST1_28d or 
	ST1_27d or ST1_26d or ST1_25d or ST1_24d or M_148 )
	begin
	rl_AD1_c1 = ( ( ( ( ( ( ( ( ( ( ( M_148 | ST1_24d ) | ST1_25d ) | ST1_26d ) | 
		ST1_27d ) | ST1_28d ) | ST1_29d ) | ST1_30d ) | ST1_31d ) | ST1_32d ) | 
		ST1_33d ) | ST1_34d ) ;	// line#=../rle.cpp:52
	rl_AD1_c2 = ( U_173 | ST1_12d ) ;	// line#=../rle.cpp:68,73,79
	rl_AD1_c3 = ( ( ( ( ( ( ( ( ( ( ( M_157 | ST1_46d ) | ST1_47d ) | ST1_48d ) | 
		ST1_49d ) | ST1_50d ) | ST1_51d ) | ST1_52d ) | ST1_53d ) | ST1_54d ) | 
		ST1_55d ) | ST1_56d ) ;
	rl_AD1 = ( ( { 7{ rl_AD1_c1 } } & { 1'h0 , TR_08 } )	// line#=../rle.cpp:52
		| ( { 7{ rl_AD1_c2 } } & RG_len_01_1 [6:0] )	// line#=../rle.cpp:68,73,79
		| ( { 7{ M_139 } } & incr8u1ot [6:0] )		// line#=../rle.cpp:68,69,73,74,79,80
		| ( { 7{ U_207 } } & RG_75_02 )			// line#=../rle.cpp:85
		| ( { 7{ rl_AD1_c3 } } & { 1'h1 , TR_12 } ) ) ;
	end
always @ ( zz_RD1 or U_237 or RG_k_quantized_block_02 or U_235 or sub12s_91ot or 
	ST1_05d )
	rl_WD1 = ( ( { 9{ ST1_05d } } & sub12s_91ot )		// line#=../rle.cpp:52
		| ( { 9{ U_235 } } & RG_k_quantized_block_02 )	// line#=../rle.cpp:73
		| ( { 9{ U_237 } } & zz_RD1 )			// line#=../rle.cpp:74
		) ;	// line#=../rle.cpp:68,69,79,80,85
assign	rl_WE1 = ( ( ( ( ( ST1_05d | U_173 ) | ST1_09d ) | U_207 ) | ST1_12d ) | 
	ST1_13d ) ;
always @ ( ST1_54d or ST1_52d or ST1_50d or ST1_48d or ST1_46d or ST1_44d or ST1_42d or 
	ST1_40d or ST1_38d or ST1_36d or ST1_33d or ST1_31d or ST1_29d or ST1_27d or 
	ST1_25d or ST1_23d or ST1_21d or ST1_19d or ST1_17d or ST1_15d or ST1_14d )
	TR_13 = ( ( { 6{ ST1_14d } } & 6'h01 )
		| ( { 6{ ST1_15d } } & 6'h02 )
		| ( { 6{ ST1_17d } } & 6'h05 )
		| ( { 6{ ST1_19d } } & 6'h08 )
		| ( { 6{ ST1_21d } } & 6'h0b )
		| ( { 6{ ST1_23d } } & 6'h0e )
		| ( { 6{ ST1_25d } } & 6'h11 )
		| ( { 6{ ST1_27d } } & 6'h14 )
		| ( { 6{ ST1_29d } } & 6'h17 )
		| ( { 6{ ST1_31d } } & 6'h1a )
		| ( { 6{ ST1_33d } } & 6'h1d )
		| ( { 6{ ST1_36d } } & 6'h21 )
		| ( { 6{ ST1_38d } } & 6'h24 )
		| ( { 6{ ST1_40d } } & 6'h27 )
		| ( { 6{ ST1_42d } } & 6'h2a )
		| ( { 6{ ST1_44d } } & 6'h2d )
		| ( { 6{ ST1_46d } } & 6'h30 )
		| ( { 6{ ST1_48d } } & 6'h33 )
		| ( { 6{ ST1_50d } } & 6'h36 )
		| ( { 6{ ST1_52d } } & 6'h39 )
		| ( { 6{ ST1_54d } } & 6'h3c ) ) ;
always @ ( ST1_56d or ST1_55d or ST1_53d or ST1_51d or ST1_49d or ST1_47d or ST1_45d or 
	ST1_43d or ST1_41d or ST1_39d or ST1_37d or ST1_35d or ST1_34d or ST1_32d or 
	ST1_30d or ST1_28d or ST1_26d or ST1_24d or ST1_22d or ST1_20d or ST1_18d or 
	ST1_16d )
	TR_14 = ( ( { 6{ ST1_16d } } & 6'h03 )
		| ( { 6{ ST1_18d } } & 6'h06 )
		| ( { 6{ ST1_20d } } & 6'h09 )
		| ( { 6{ ST1_22d } } & 6'h0c )
		| ( { 6{ ST1_24d } } & 6'h0f )
		| ( { 6{ ST1_26d } } & 6'h12 )
		| ( { 6{ ST1_28d } } & 6'h15 )
		| ( { 6{ ST1_30d } } & 6'h18 )
		| ( { 6{ ST1_32d } } & 6'h1b )
		| ( { 6{ ST1_34d } } & 6'h1e )
		| ( { 6{ ST1_35d } } & 6'h1f )
		| ( { 6{ ST1_37d } } & 6'h22 )
		| ( { 6{ ST1_39d } } & 6'h25 )
		| ( { 6{ ST1_41d } } & 6'h28 )
		| ( { 6{ ST1_43d } } & 6'h2b )
		| ( { 6{ ST1_45d } } & 6'h2e )
		| ( { 6{ ST1_47d } } & 6'h31 )
		| ( { 6{ ST1_49d } } & 6'h34 )
		| ( { 6{ ST1_51d } } & 6'h37 )
		| ( { 6{ ST1_53d } } & 6'h3a )
		| ( { 6{ ST1_55d } } & 6'h3d )
		| ( { 6{ ST1_56d } } & 6'h3f ) ) ;
always @ ( TR_14 or ST1_56d or M_145 or TR_13 or M_143 or RG_k_01_1 or M_138 )
	begin
	rl_RA2_c1 = ( M_145 | ST1_56d ) ;
	rl_RA2 = ( ( { 7{ M_138 } } & RG_k_01_1 )	// line#=../rle.cpp:77,78,83,84
		| ( { 7{ M_143 } } & { TR_13 , 1'h0 } )
		| ( { 7{ rl_RA2_c1 } } & { TR_14 , 1'h1 } ) ) ;
	end
always @ ( ST1_54d or ST1_52d or ST1_50d or ST1_48d or ST1_46d or ST1_44d or ST1_42d or 
	ST1_40d or ST1_38d or ST1_36d or ST1_33d or ST1_31d or ST1_29d or ST1_27d or 
	ST1_25d or ST1_23d or ST1_21d or ST1_19d or ST1_17d or ST1_15d )
	TR_15 = ( ( { 6{ ST1_15d } } & 6'h01 )
		| ( { 6{ ST1_17d } } & 6'h04 )
		| ( { 6{ ST1_19d } } & 6'h07 )
		| ( { 6{ ST1_21d } } & 6'h0a )
		| ( { 6{ ST1_23d } } & 6'h0d )
		| ( { 6{ ST1_25d } } & 6'h10 )
		| ( { 6{ ST1_27d } } & 6'h13 )
		| ( { 6{ ST1_29d } } & 6'h16 )
		| ( { 6{ ST1_31d } } & 6'h19 )
		| ( { 6{ ST1_33d } } & 6'h1c )
		| ( { 6{ ST1_36d } } & 6'h21 )
		| ( { 6{ ST1_38d } } & 6'h24 )
		| ( { 6{ ST1_40d } } & 6'h27 )
		| ( { 6{ ST1_42d } } & 6'h2a )
		| ( { 6{ ST1_44d } } & 6'h2d )
		| ( { 6{ ST1_46d } } & 6'h30 )
		| ( { 6{ ST1_48d } } & 6'h33 )
		| ( { 6{ ST1_50d } } & 6'h36 )
		| ( { 6{ ST1_52d } } & 6'h39 )
		| ( { 6{ ST1_54d } } & 6'h3c ) ) ;
always @ ( ST1_55d or ST1_53d or ST1_51d or ST1_49d or ST1_47d or ST1_45d or ST1_43d or 
	ST1_41d or ST1_39d or ST1_37d or ST1_35d or ST1_34d or ST1_32d or ST1_30d or 
	ST1_28d or ST1_26d or ST1_24d or ST1_22d or ST1_20d or ST1_18d or ST1_16d )
	TR_16 = ( ( { 6{ ST1_16d } } & 6'h03 )
		| ( { 6{ ST1_18d } } & 6'h06 )
		| ( { 6{ ST1_20d } } & 6'h09 )
		| ( { 6{ ST1_22d } } & 6'h0c )
		| ( { 6{ ST1_24d } } & 6'h0f )
		| ( { 6{ ST1_26d } } & 6'h12 )
		| ( { 6{ ST1_28d } } & 6'h15 )
		| ( { 6{ ST1_30d } } & 6'h18 )
		| ( { 6{ ST1_32d } } & 6'h1b )
		| ( { 6{ ST1_34d } } & 6'h1e )
		| ( { 6{ ST1_35d } } & 6'h20 )
		| ( { 6{ ST1_37d } } & 6'h23 )
		| ( { 6{ ST1_39d } } & 6'h26 )
		| ( { 6{ ST1_41d } } & 6'h29 )
		| ( { 6{ ST1_43d } } & 6'h2c )
		| ( { 6{ ST1_45d } } & 6'h2f )
		| ( { 6{ ST1_47d } } & 6'h32 )
		| ( { 6{ ST1_49d } } & 6'h35 )
		| ( { 6{ ST1_51d } } & 6'h38 )
		| ( { 6{ ST1_53d } } & 6'h3b )
		| ( { 6{ ST1_55d } } & 6'h3e ) ) ;
assign	M_143 = ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ST1_14d | ST1_15d ) | ST1_17d ) | 
	ST1_19d ) | ST1_21d ) | ST1_23d ) | ST1_25d ) | ST1_27d ) | ST1_29d ) | ST1_31d ) | 
	ST1_33d ) | ST1_36d ) | ST1_38d ) | ST1_40d ) | ST1_42d ) | ST1_44d ) | ST1_46d ) | 
	ST1_48d ) | ST1_50d ) | ST1_52d ) | ST1_54d ) ;
assign	M_145 = ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ST1_16d | ST1_18d ) | ST1_20d ) | 
	ST1_22d ) | ST1_24d ) | ST1_26d ) | ST1_28d ) | ST1_30d ) | ST1_32d ) | ST1_34d ) | 
	ST1_35d ) | ST1_37d ) | ST1_39d ) | ST1_41d ) | ST1_43d ) | ST1_45d ) | ST1_47d ) | 
	ST1_49d ) | ST1_51d ) | ST1_53d ) | ST1_55d ) ;
always @ ( TR_16 or M_145 or TR_15 or M_143 or RG_80_01 or M_138 )
	rl_RA3 = ( ( { 7{ M_138 } } & RG_80_01 )
		| ( { 7{ M_143 } } & { TR_15 , 1'h1 } )
		| ( { 7{ M_145 } } & { TR_16 , 1'h0 } ) ) ;

endmodule

module jpeg_sub8u_7_1 ( i1 ,i2 ,o1 );
input	[6:0]	i1 ;
input	[1:0]	i2 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - { 5'h00 , i2 } ) ;

endmodule

module jpeg_sub8u_7 ( i1 ,i2 ,o1 );
input	[6:0]	i1 ;
input	[2:0]	i2 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - { 4'h0 , i2 } ) ;

endmodule

module jpeg_decr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_decr8u_7 ( i1 ,o1 );
input	[6:0]	i1 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_incr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr8u ( i1 ,o1 );
input	[7:0]	i1 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr4s ( i1 ,o1 );
input	[3:0]	i1 ;
output	[3:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_lop8u_1 ( i1 ,i2 ,o1 );
input	[5:0]	i1 ;
input	[5:0]	i2 ;
output		o1 ;
wire		M_01 ;

assign	M_01 = ( i1 < i2 ) ;
assign	o1 = M_01 ;

endmodule

module jpeg_sub12s_9 ( i1 ,i2 ,o1 );
input	[8:0]	i1 ;
input	[8:0]	i2 ;
output	[8:0]	o1 ;

assign	o1 = ( i1 - i2 ) ;

endmodule

module jpeg_sub8u ( i1 ,i2 ,o1 );
input	[7:0]	i1 ;
input	[1:0]	i2 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 - { 6'h00 , i2 } ) ;

endmodule

module jpeg_MEM_rl ( AD1 ,RD1 ,WD1 ,WE1 ,CLK1 ,RA2 ,RD2 ,RA3 ,RD3 );
input	[6:0]	AD1 ;
output	[8:0]	RD1 ;
input	[8:0]	WD1 ;
input		WE1 ;
input		CLK1 ;
input	[6:0]	RA2 ;
output	[8:0]	RD2 ;
input	[6:0]	RA3 ;
output	[8:0]	RD3 ;

jpeg_MEM_rl_subD INST_MEM_rl_subD_1 ( .RD1(RD1) ,.AD1(AD1) ,.WE1(WE1) ,.WD1(WD1) ,
	.CLK1(CLK1) ,.RD2(RD2) ,.RA2(RA2) );
jpeg_MEM_rl_subD INST_MEM_rl_subD_2 ( .RD1() ,.AD1(AD1) ,.WE1(WE1) ,.WD1(WD1) ,.CLK1(CLK1) ,
	.RD2(RD3) ,.RA2(RA3) );

endmodule

(* ram_extract = "yes" *)
module jpeg_MEM_rl_subD ( RD1 ,AD1 ,WE1 ,WD1 ,CLK1 ,RD2 ,RA2 );
output	[8:0]	RD1 ;
input	[6:0]	AD1 ;
input		WE1 ;
input	[8:0]	WD1 ;
input		CLK1 ;
output	[8:0]	RD2 ;
input	[6:0]	RA2 ;
(* ram_style = "distributed" *)reg	[8:0]	rl_r	[0:127] ;

assign	RD1 = rl_r[AD1] ;
assign	RD2 = rl_r[RA2] ;

always @ ( posedge CLK1 )
	begin
	if ( WE1 )
		rl_r [AD1] = WD1 ;
	end

endmodule

module jpeg_MEMB9W64 ( RA1 ,RD1 ,RCLK1 ,WA2 ,WD2 ,WE2 ,WCLK2 );
input	[5:0]	RA1 ;
output	[8:0]	RD1 ;
input		RCLK1 ;
input	[5:0]	WA2 ;
input	[8:0]	WD2 ;
input		WE2 ;
input		WCLK2 ;

jpeg_MEMB9W64_sub INST_MEMB9W64_sub_1 ( .RD1(RD1) ,.WE2(WE2) ,.WD2(WD2) ,.RA1(RA1) ,
	.WA2(WA2) ,.RCLK1(RCLK1) ,.WCLK2(WCLK2) );

endmodule

(* ram_extract = "yes" *)
module jpeg_MEMB9W64_sub ( RD1 ,WE2 ,WD2 ,RA1 ,WA2 ,RCLK1 ,WCLK2 );
output	[8:0]	RD1 ;
input		WE2 ;
input	[8:0]	WD2 ;
input	[5:0]	RA1 ;
input	[5:0]	WA2 ;
input		RCLK1 ;
input		WCLK2 ;
wire		Wen1_wire ;
reg	[8:0]	Rd1_sr	[0:0] ;
(* ram_style = "block" *)reg	[8:0]	MEMB9W64_r	[0:63] ;

assign	RD1 = Rd1_sr[0] ;
assign	Wen1_wire = WE2 ;

always @ ( posedge RCLK1 )
	begin
	Rd1_sr [0] <= MEMB9W64_r[RA1] ;
	end

always @ ( posedge WCLK2 )
	begin
	if ( Wen1_wire )
		begin
		MEMB9W64_r [WA2] <= WD2 ;
		end
	end

endmodule
