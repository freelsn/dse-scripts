// verilog_out version 6.79.2
// options:  veriloggen jpeg_E.IFF
// bdlpars options:  -DDSE ../rle.cpp
// bdltran options:  -c1000 -s -Zresource_fcnt=GENERATE -Zresource_mcnt=GENERATE -lb /home/shuangnan/share/packages/zynq-1.BLIB -lfl /home/shuangnan/share/packages/zynq-1.FLIB jpeg.IFF -OX -a8196 -Zfu_cnt_incr_rate=0 -tcio 
// timestamp_0: 20180213182006_17614_49326
// timestamp_5: 20180213182011_18893_64049
// timestamp_9: 20180213182017_18893_31186
// timestamp_C: 20180213182016_18893_00614
// timestamp_E: 20180213182017_18893_35777
// timestamp_V: 20180213182021_21327_87221

module jpeg ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,jpeg_in_a04 ,
	jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,jpeg_in_a10 ,
	jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,jpeg_in_a16 ,
	jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,jpeg_in_a22 ,
	jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,jpeg_in_a28 ,
	jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,jpeg_in_a34 ,
	jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,jpeg_in_a40 ,
	jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,jpeg_in_a46 ,
	jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,jpeg_in_a52 ,
	jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,jpeg_in_a58 ,
	jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,jpeg_in_a64 ,
	jpeg_in_a65 ,jpeg_in_a66 ,jpeg_in_a67 ,jpeg_in_a68 ,jpeg_in_a69 ,jpeg_in_a70 ,
	jpeg_in_a71 ,jpeg_in_a72 ,jpeg_in_a73 ,jpeg_in_a74 ,jpeg_in_a75 ,jpeg_in_a76 ,
	jpeg_in_a77 ,jpeg_in_a78 ,jpeg_in_a79 ,jpeg_in_a80 ,jpeg_in_a81 ,jpeg_in_a82 ,
	jpeg_in_a83 ,jpeg_in_a84 ,jpeg_in_a85 ,jpeg_in_a86 ,jpeg_in_a87 ,jpeg_in_a88 ,
	jpeg_in_a89 ,jpeg_in_a90 ,jpeg_in_a91 ,jpeg_in_a92 ,jpeg_in_a93 ,jpeg_in_a94 ,
	jpeg_in_a95 ,jpeg_in_a96 ,jpeg_in_a97 ,jpeg_in_a98 ,jpeg_in_a99 ,jpeg_in_a100 ,
	jpeg_in_a101 ,jpeg_in_a102 ,jpeg_in_a103 ,jpeg_in_a104 ,jpeg_in_a105 ,jpeg_in_a106 ,
	jpeg_in_a107 ,jpeg_in_a108 ,jpeg_in_a109 ,jpeg_in_a110 ,jpeg_in_a111 ,jpeg_in_a112 ,
	jpeg_in_a113 ,jpeg_in_a114 ,jpeg_in_a115 ,jpeg_in_a116 ,jpeg_in_a117 ,jpeg_in_a118 ,
	jpeg_in_a119 ,jpeg_in_a120 ,jpeg_in_a121 ,jpeg_in_a122 ,jpeg_in_a123 ,jpeg_in_a124 ,
	jpeg_in_a125 ,jpeg_in_a126 ,jpeg_in_a127 ,jpeg_len_in ,jpeg_out_a00 ,jpeg_out_a01 ,
	jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,jpeg_out_a06 ,jpeg_out_a07 ,
	jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,jpeg_out_a12 ,jpeg_out_a13 ,
	jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,jpeg_out_a18 ,jpeg_out_a19 ,
	jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,jpeg_out_a24 ,jpeg_out_a25 ,
	jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,jpeg_out_a30 ,jpeg_out_a31 ,
	jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,jpeg_out_a36 ,jpeg_out_a37 ,
	jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,jpeg_out_a42 ,jpeg_out_a43 ,
	jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,jpeg_out_a48 ,jpeg_out_a49 ,
	jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,jpeg_out_a54 ,jpeg_out_a55 ,
	jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,jpeg_out_a60 ,jpeg_out_a61 ,
	jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,jpeg_out_a66 ,jpeg_out_a67 ,
	jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,jpeg_out_a72 ,jpeg_out_a73 ,
	jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,jpeg_out_a78 ,jpeg_out_a79 ,
	jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,jpeg_out_a84 ,jpeg_out_a85 ,
	jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,jpeg_out_a90 ,jpeg_out_a91 ,
	jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,jpeg_out_a96 ,jpeg_out_a97 ,
	jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,jpeg_out_a102 ,
	jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,jpeg_out_a107 ,
	jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,jpeg_out_a112 ,
	jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,jpeg_out_a117 ,
	jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,jpeg_out_a122 ,
	jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,jpeg_out_a127 ,
	jpeg_len_out ,valid );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a64 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a65 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a66 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a67 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a68 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a69 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a70 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a71 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a72 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a73 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a74 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a75 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a76 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a77 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a78 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a79 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a80 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a81 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a82 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a83 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a84 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a85 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a86 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a87 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a88 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a89 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a90 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a91 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a92 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a93 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a94 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a95 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a96 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a97 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a98 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a99 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a100 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a101 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a102 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a103 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a104 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a105 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a106 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a107 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a108 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a109 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a110 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a111 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a112 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a113 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a114 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a115 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a116 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a117 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a118 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a119 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a120 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a121 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a122 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a123 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a124 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a125 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a126 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a127 ;	// line#=../rle.h:56
input	[11:0]	jpeg_len_in ;	// line#=../rle.h:57
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
wire		ST1_01d ;
wire		ST1_02d ;
wire		ST1_03d ;
wire		ST1_04d ;
wire		ST1_05d ;
wire		ST1_06d ;
wire		ST1_07d ;
wire		ST1_08d ;
wire		ST1_09d ;
wire		ST1_10d ;
wire		ST1_11d ;
wire		ST1_12d ;
wire		ST1_13d ;
wire		ST1_14d ;
wire		ST1_15d ;
wire		JF_01 ;
wire		FL01_01_Leos_all ;
wire		lop8u_11ot ;
wire		JF_05 ;
wire		FL02_01_Leos_all ;
wire		JF_08 ;
wire		JF_09 ;
wire		JF_10 ;
wire		FL01_02_01_stall ;

jpeg_fsm INST_fsm ( .clk(clk) ,.rst(rst) ,.ST1_15d(ST1_15d) ,.ST1_14d(ST1_14d) ,
	.ST1_13d(ST1_13d) ,.ST1_12d(ST1_12d) ,.ST1_11d(ST1_11d) ,.ST1_10d(ST1_10d) ,
	.ST1_09d(ST1_09d) ,.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,.ST1_06d(ST1_06d) ,
	.ST1_05d(ST1_05d) ,.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,.ST1_02d(ST1_02d) ,
	.ST1_01d(ST1_01d) ,.JF_01(JF_01) ,.FL01_01_Leos_all(FL01_01_Leos_all) ,.lop8u_11ot(lop8u_11ot) ,
	.JF_05(JF_05) ,.FL02_01_Leos_all(FL02_01_Leos_all) ,.JF_08(JF_08) ,.JF_09(JF_09) ,
	.JF_10(JF_10) ,.FL01_02_01_stall(FL01_02_01_stall) );
jpeg_dat INST_dat ( .clk(clk) ,.rst(rst) ,.jpeg_in_a00(jpeg_in_a00) ,.jpeg_in_a01(jpeg_in_a01) ,
	.jpeg_in_a02(jpeg_in_a02) ,.jpeg_in_a03(jpeg_in_a03) ,.jpeg_in_a04(jpeg_in_a04) ,
	.jpeg_in_a05(jpeg_in_a05) ,.jpeg_in_a06(jpeg_in_a06) ,.jpeg_in_a07(jpeg_in_a07) ,
	.jpeg_in_a08(jpeg_in_a08) ,.jpeg_in_a09(jpeg_in_a09) ,.jpeg_in_a10(jpeg_in_a10) ,
	.jpeg_in_a11(jpeg_in_a11) ,.jpeg_in_a12(jpeg_in_a12) ,.jpeg_in_a13(jpeg_in_a13) ,
	.jpeg_in_a14(jpeg_in_a14) ,.jpeg_in_a15(jpeg_in_a15) ,.jpeg_in_a16(jpeg_in_a16) ,
	.jpeg_in_a17(jpeg_in_a17) ,.jpeg_in_a18(jpeg_in_a18) ,.jpeg_in_a19(jpeg_in_a19) ,
	.jpeg_in_a20(jpeg_in_a20) ,.jpeg_in_a21(jpeg_in_a21) ,.jpeg_in_a22(jpeg_in_a22) ,
	.jpeg_in_a23(jpeg_in_a23) ,.jpeg_in_a24(jpeg_in_a24) ,.jpeg_in_a25(jpeg_in_a25) ,
	.jpeg_in_a26(jpeg_in_a26) ,.jpeg_in_a27(jpeg_in_a27) ,.jpeg_in_a28(jpeg_in_a28) ,
	.jpeg_in_a29(jpeg_in_a29) ,.jpeg_in_a30(jpeg_in_a30) ,.jpeg_in_a31(jpeg_in_a31) ,
	.jpeg_in_a32(jpeg_in_a32) ,.jpeg_in_a33(jpeg_in_a33) ,.jpeg_in_a34(jpeg_in_a34) ,
	.jpeg_in_a35(jpeg_in_a35) ,.jpeg_in_a36(jpeg_in_a36) ,.jpeg_in_a37(jpeg_in_a37) ,
	.jpeg_in_a38(jpeg_in_a38) ,.jpeg_in_a39(jpeg_in_a39) ,.jpeg_in_a40(jpeg_in_a40) ,
	.jpeg_in_a41(jpeg_in_a41) ,.jpeg_in_a42(jpeg_in_a42) ,.jpeg_in_a43(jpeg_in_a43) ,
	.jpeg_in_a44(jpeg_in_a44) ,.jpeg_in_a45(jpeg_in_a45) ,.jpeg_in_a46(jpeg_in_a46) ,
	.jpeg_in_a47(jpeg_in_a47) ,.jpeg_in_a48(jpeg_in_a48) ,.jpeg_in_a49(jpeg_in_a49) ,
	.jpeg_in_a50(jpeg_in_a50) ,.jpeg_in_a51(jpeg_in_a51) ,.jpeg_in_a52(jpeg_in_a52) ,
	.jpeg_in_a53(jpeg_in_a53) ,.jpeg_in_a54(jpeg_in_a54) ,.jpeg_in_a55(jpeg_in_a55) ,
	.jpeg_in_a56(jpeg_in_a56) ,.jpeg_in_a57(jpeg_in_a57) ,.jpeg_in_a58(jpeg_in_a58) ,
	.jpeg_in_a59(jpeg_in_a59) ,.jpeg_in_a60(jpeg_in_a60) ,.jpeg_in_a61(jpeg_in_a61) ,
	.jpeg_in_a62(jpeg_in_a62) ,.jpeg_in_a63(jpeg_in_a63) ,.jpeg_in_a64(jpeg_in_a64) ,
	.jpeg_in_a65(jpeg_in_a65) ,.jpeg_in_a66(jpeg_in_a66) ,.jpeg_in_a67(jpeg_in_a67) ,
	.jpeg_in_a68(jpeg_in_a68) ,.jpeg_in_a69(jpeg_in_a69) ,.jpeg_in_a70(jpeg_in_a70) ,
	.jpeg_in_a71(jpeg_in_a71) ,.jpeg_in_a72(jpeg_in_a72) ,.jpeg_in_a73(jpeg_in_a73) ,
	.jpeg_in_a74(jpeg_in_a74) ,.jpeg_in_a75(jpeg_in_a75) ,.jpeg_in_a76(jpeg_in_a76) ,
	.jpeg_in_a77(jpeg_in_a77) ,.jpeg_in_a78(jpeg_in_a78) ,.jpeg_in_a79(jpeg_in_a79) ,
	.jpeg_in_a80(jpeg_in_a80) ,.jpeg_in_a81(jpeg_in_a81) ,.jpeg_in_a82(jpeg_in_a82) ,
	.jpeg_in_a83(jpeg_in_a83) ,.jpeg_in_a84(jpeg_in_a84) ,.jpeg_in_a85(jpeg_in_a85) ,
	.jpeg_in_a86(jpeg_in_a86) ,.jpeg_in_a87(jpeg_in_a87) ,.jpeg_in_a88(jpeg_in_a88) ,
	.jpeg_in_a89(jpeg_in_a89) ,.jpeg_in_a90(jpeg_in_a90) ,.jpeg_in_a91(jpeg_in_a91) ,
	.jpeg_in_a92(jpeg_in_a92) ,.jpeg_in_a93(jpeg_in_a93) ,.jpeg_in_a94(jpeg_in_a94) ,
	.jpeg_in_a95(jpeg_in_a95) ,.jpeg_in_a96(jpeg_in_a96) ,.jpeg_in_a97(jpeg_in_a97) ,
	.jpeg_in_a98(jpeg_in_a98) ,.jpeg_in_a99(jpeg_in_a99) ,.jpeg_in_a100(jpeg_in_a100) ,
	.jpeg_in_a101(jpeg_in_a101) ,.jpeg_in_a102(jpeg_in_a102) ,.jpeg_in_a103(jpeg_in_a103) ,
	.jpeg_in_a104(jpeg_in_a104) ,.jpeg_in_a105(jpeg_in_a105) ,.jpeg_in_a106(jpeg_in_a106) ,
	.jpeg_in_a107(jpeg_in_a107) ,.jpeg_in_a108(jpeg_in_a108) ,.jpeg_in_a109(jpeg_in_a109) ,
	.jpeg_in_a110(jpeg_in_a110) ,.jpeg_in_a111(jpeg_in_a111) ,.jpeg_in_a112(jpeg_in_a112) ,
	.jpeg_in_a113(jpeg_in_a113) ,.jpeg_in_a114(jpeg_in_a114) ,.jpeg_in_a115(jpeg_in_a115) ,
	.jpeg_in_a116(jpeg_in_a116) ,.jpeg_in_a117(jpeg_in_a117) ,.jpeg_in_a118(jpeg_in_a118) ,
	.jpeg_in_a119(jpeg_in_a119) ,.jpeg_in_a120(jpeg_in_a120) ,.jpeg_in_a121(jpeg_in_a121) ,
	.jpeg_in_a122(jpeg_in_a122) ,.jpeg_in_a123(jpeg_in_a123) ,.jpeg_in_a124(jpeg_in_a124) ,
	.jpeg_in_a125(jpeg_in_a125) ,.jpeg_in_a126(jpeg_in_a126) ,.jpeg_in_a127(jpeg_in_a127) ,
	.jpeg_out_a00(jpeg_out_a00) ,.jpeg_out_a01(jpeg_out_a01) ,.jpeg_out_a02(jpeg_out_a02) ,
	.jpeg_out_a03(jpeg_out_a03) ,.jpeg_out_a04(jpeg_out_a04) ,.jpeg_out_a05(jpeg_out_a05) ,
	.jpeg_out_a06(jpeg_out_a06) ,.jpeg_out_a07(jpeg_out_a07) ,.jpeg_out_a08(jpeg_out_a08) ,
	.jpeg_out_a09(jpeg_out_a09) ,.jpeg_out_a10(jpeg_out_a10) ,.jpeg_out_a11(jpeg_out_a11) ,
	.jpeg_out_a12(jpeg_out_a12) ,.jpeg_out_a13(jpeg_out_a13) ,.jpeg_out_a14(jpeg_out_a14) ,
	.jpeg_out_a15(jpeg_out_a15) ,.jpeg_out_a16(jpeg_out_a16) ,.jpeg_out_a17(jpeg_out_a17) ,
	.jpeg_out_a18(jpeg_out_a18) ,.jpeg_out_a19(jpeg_out_a19) ,.jpeg_out_a20(jpeg_out_a20) ,
	.jpeg_out_a21(jpeg_out_a21) ,.jpeg_out_a22(jpeg_out_a22) ,.jpeg_out_a23(jpeg_out_a23) ,
	.jpeg_out_a24(jpeg_out_a24) ,.jpeg_out_a25(jpeg_out_a25) ,.jpeg_out_a26(jpeg_out_a26) ,
	.jpeg_out_a27(jpeg_out_a27) ,.jpeg_out_a28(jpeg_out_a28) ,.jpeg_out_a29(jpeg_out_a29) ,
	.jpeg_out_a30(jpeg_out_a30) ,.jpeg_out_a31(jpeg_out_a31) ,.jpeg_out_a32(jpeg_out_a32) ,
	.jpeg_out_a33(jpeg_out_a33) ,.jpeg_out_a34(jpeg_out_a34) ,.jpeg_out_a35(jpeg_out_a35) ,
	.jpeg_out_a36(jpeg_out_a36) ,.jpeg_out_a37(jpeg_out_a37) ,.jpeg_out_a38(jpeg_out_a38) ,
	.jpeg_out_a39(jpeg_out_a39) ,.jpeg_out_a40(jpeg_out_a40) ,.jpeg_out_a41(jpeg_out_a41) ,
	.jpeg_out_a42(jpeg_out_a42) ,.jpeg_out_a43(jpeg_out_a43) ,.jpeg_out_a44(jpeg_out_a44) ,
	.jpeg_out_a45(jpeg_out_a45) ,.jpeg_out_a46(jpeg_out_a46) ,.jpeg_out_a47(jpeg_out_a47) ,
	.jpeg_out_a48(jpeg_out_a48) ,.jpeg_out_a49(jpeg_out_a49) ,.jpeg_out_a50(jpeg_out_a50) ,
	.jpeg_out_a51(jpeg_out_a51) ,.jpeg_out_a52(jpeg_out_a52) ,.jpeg_out_a53(jpeg_out_a53) ,
	.jpeg_out_a54(jpeg_out_a54) ,.jpeg_out_a55(jpeg_out_a55) ,.jpeg_out_a56(jpeg_out_a56) ,
	.jpeg_out_a57(jpeg_out_a57) ,.jpeg_out_a58(jpeg_out_a58) ,.jpeg_out_a59(jpeg_out_a59) ,
	.jpeg_out_a60(jpeg_out_a60) ,.jpeg_out_a61(jpeg_out_a61) ,.jpeg_out_a62(jpeg_out_a62) ,
	.jpeg_out_a63(jpeg_out_a63) ,.jpeg_out_a64(jpeg_out_a64) ,.jpeg_out_a65(jpeg_out_a65) ,
	.jpeg_out_a66(jpeg_out_a66) ,.jpeg_out_a67(jpeg_out_a67) ,.jpeg_out_a68(jpeg_out_a68) ,
	.jpeg_out_a69(jpeg_out_a69) ,.jpeg_out_a70(jpeg_out_a70) ,.jpeg_out_a71(jpeg_out_a71) ,
	.jpeg_out_a72(jpeg_out_a72) ,.jpeg_out_a73(jpeg_out_a73) ,.jpeg_out_a74(jpeg_out_a74) ,
	.jpeg_out_a75(jpeg_out_a75) ,.jpeg_out_a76(jpeg_out_a76) ,.jpeg_out_a77(jpeg_out_a77) ,
	.jpeg_out_a78(jpeg_out_a78) ,.jpeg_out_a79(jpeg_out_a79) ,.jpeg_out_a80(jpeg_out_a80) ,
	.jpeg_out_a81(jpeg_out_a81) ,.jpeg_out_a82(jpeg_out_a82) ,.jpeg_out_a83(jpeg_out_a83) ,
	.jpeg_out_a84(jpeg_out_a84) ,.jpeg_out_a85(jpeg_out_a85) ,.jpeg_out_a86(jpeg_out_a86) ,
	.jpeg_out_a87(jpeg_out_a87) ,.jpeg_out_a88(jpeg_out_a88) ,.jpeg_out_a89(jpeg_out_a89) ,
	.jpeg_out_a90(jpeg_out_a90) ,.jpeg_out_a91(jpeg_out_a91) ,.jpeg_out_a92(jpeg_out_a92) ,
	.jpeg_out_a93(jpeg_out_a93) ,.jpeg_out_a94(jpeg_out_a94) ,.jpeg_out_a95(jpeg_out_a95) ,
	.jpeg_out_a96(jpeg_out_a96) ,.jpeg_out_a97(jpeg_out_a97) ,.jpeg_out_a98(jpeg_out_a98) ,
	.jpeg_out_a99(jpeg_out_a99) ,.jpeg_out_a100(jpeg_out_a100) ,.jpeg_out_a101(jpeg_out_a101) ,
	.jpeg_out_a102(jpeg_out_a102) ,.jpeg_out_a103(jpeg_out_a103) ,.jpeg_out_a104(jpeg_out_a104) ,
	.jpeg_out_a105(jpeg_out_a105) ,.jpeg_out_a106(jpeg_out_a106) ,.jpeg_out_a107(jpeg_out_a107) ,
	.jpeg_out_a108(jpeg_out_a108) ,.jpeg_out_a109(jpeg_out_a109) ,.jpeg_out_a110(jpeg_out_a110) ,
	.jpeg_out_a111(jpeg_out_a111) ,.jpeg_out_a112(jpeg_out_a112) ,.jpeg_out_a113(jpeg_out_a113) ,
	.jpeg_out_a114(jpeg_out_a114) ,.jpeg_out_a115(jpeg_out_a115) ,.jpeg_out_a116(jpeg_out_a116) ,
	.jpeg_out_a117(jpeg_out_a117) ,.jpeg_out_a118(jpeg_out_a118) ,.jpeg_out_a119(jpeg_out_a119) ,
	.jpeg_out_a120(jpeg_out_a120) ,.jpeg_out_a121(jpeg_out_a121) ,.jpeg_out_a122(jpeg_out_a122) ,
	.jpeg_out_a123(jpeg_out_a123) ,.jpeg_out_a124(jpeg_out_a124) ,.jpeg_out_a125(jpeg_out_a125) ,
	.jpeg_out_a126(jpeg_out_a126) ,.jpeg_out_a127(jpeg_out_a127) ,.jpeg_len_out(jpeg_len_out) ,
	.valid(valid) ,.ST1_15d(ST1_15d) ,.ST1_14d(ST1_14d) ,.ST1_13d(ST1_13d) ,
	.ST1_12d(ST1_12d) ,.ST1_11d(ST1_11d) ,.ST1_10d(ST1_10d) ,.ST1_09d(ST1_09d) ,
	.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,
	.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,
	.JF_01_port(JF_01) ,.FL01_01_Leos_all(FL01_01_Leos_all) ,.lop8u_11ot_port(lop8u_11ot) ,
	.JF_05(JF_05) ,.FL02_01_Leos_all(FL02_01_Leos_all) ,.JF_08(JF_08) ,.JF_09(JF_09) ,
	.JF_10(JF_10) ,.FL01_02_01_stall_port(FL01_02_01_stall) );

endmodule

module jpeg_fsm ( clk ,rst ,ST1_15d ,ST1_14d ,ST1_13d ,ST1_12d ,ST1_11d ,ST1_10d ,
	ST1_09d ,ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,ST1_02d ,
	ST1_01d ,JF_01 ,FL01_01_Leos_all ,lop8u_11ot ,JF_05 ,FL02_01_Leos_all ,JF_08 ,
	JF_09 ,JF_10 ,FL01_02_01_stall );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
output		ST1_15d ;
output		ST1_14d ;
output		ST1_13d ;
output		ST1_12d ;
output		ST1_11d ;
output		ST1_10d ;
output		ST1_09d ;
output		ST1_08d ;
output		ST1_07d ;
output		ST1_06d ;
output		ST1_05d ;
output		ST1_04d ;
output		ST1_03d ;
output		ST1_02d ;
output		ST1_01d ;
input		JF_01 ;
input		FL01_01_Leos_all ;
input		lop8u_11ot ;
input		JF_05 ;
input		FL02_01_Leos_all ;
input		JF_08 ;
input		JF_09 ;
input		JF_10 ;
input		FL01_02_01_stall ;
reg	[3:0]	B01_streg ;

parameter	ST1_01 = 4'h0 ;
parameter	ST1_02 = 4'h1 ;
parameter	ST1_03 = 4'h2 ;
parameter	ST1_04 = 4'h3 ;
parameter	ST1_05 = 4'h4 ;
parameter	ST1_06 = 4'h5 ;
parameter	ST1_07 = 4'h6 ;
parameter	ST1_08 = 4'h7 ;
parameter	ST1_09 = 4'h8 ;
parameter	ST1_10 = 4'h9 ;
parameter	ST1_11 = 4'ha ;
parameter	ST1_12 = 4'hb ;
parameter	ST1_13 = 4'hc ;
parameter	ST1_14 = 4'hd ;
parameter	ST1_15 = 4'he ;

assign	ST1_01d = ( ( B01_streg == ST1_01 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_02d = ( ( B01_streg == ST1_02 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_03d = ( ( B01_streg == ST1_03 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_04d = ( ( B01_streg == ST1_04 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_05d = ( ( B01_streg == ST1_05 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_06d = ( ( B01_streg == ST1_06 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_07d = ( ( B01_streg == ST1_07 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_08d = ( ( B01_streg == ST1_08 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_09d = ( ( B01_streg == ST1_09 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_10d = ( ( B01_streg == ST1_10 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_11d = ( ( B01_streg == ST1_11 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_12d = ( ( B01_streg == ST1_12 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_13d = ( ( B01_streg == ST1_13 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_14d = ( ( B01_streg == ST1_14 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_15d = ( ( B01_streg == ST1_15 ) ? 1'h1 : 1'h0 ) ;
always @ ( posedge clk )
	if ( !rst )
		B01_streg <= ST1_01 ;
	else if ( !FL01_02_01_stall )
		case ( B01_streg )
		ST1_01 :
			B01_streg <= ST1_02 ;
		ST1_02 :
			if ( ( JF_01 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_03 ;
		ST1_03 :
			if ( ( FL01_01_Leos_all != 1'h0 ) )
				B01_streg <= ST1_04 ;
			else
				B01_streg <= ST1_03 ;
		ST1_04 :
			B01_streg <= ST1_05 ;
		ST1_05 :
			if ( ( lop8u_11ot != 1'h0 ) )
				B01_streg <= ST1_05 ;
			else
				B01_streg <= ST1_06 ;
		ST1_06 :
			if ( ( JF_05 != 1'h0 ) )
				B01_streg <= ST1_06 ;
			else
				B01_streg <= ST1_07 ;
		ST1_07 :
			B01_streg <= ST1_08 ;
		ST1_08 :
			if ( ( FL02_01_Leos_all != 1'h0 ) )
				B01_streg <= ST1_09 ;
			else
				B01_streg <= ST1_08 ;
		ST1_09 :
			if ( ( JF_08 != 1'h0 ) )
				B01_streg <= ST1_10 ;
			else
				B01_streg <= ST1_11 ;
		ST1_10 :
			B01_streg <= ST1_11 ;
		ST1_11 :
			if ( ( JF_09 != 1'h0 ) )
				B01_streg <= ST1_12 ;
			else
				B01_streg <= ST1_13 ;
		ST1_12 :
			B01_streg <= ST1_13 ;
		ST1_13 :
			B01_streg <= ST1_14 ;
		ST1_14 :
			if ( ( JF_10 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_15 ;
		ST1_15 :
			B01_streg <= ST1_13 ;
		default :
			B01_streg <= ST1_01 ;
		endcase

endmodule

module jpeg_dat ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,
	jpeg_in_a04 ,jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,
	jpeg_in_a10 ,jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,
	jpeg_in_a16 ,jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,
	jpeg_in_a22 ,jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,
	jpeg_in_a28 ,jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,
	jpeg_in_a34 ,jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,
	jpeg_in_a40 ,jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,
	jpeg_in_a46 ,jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,
	jpeg_in_a52 ,jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,
	jpeg_in_a58 ,jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,
	jpeg_in_a64 ,jpeg_in_a65 ,jpeg_in_a66 ,jpeg_in_a67 ,jpeg_in_a68 ,jpeg_in_a69 ,
	jpeg_in_a70 ,jpeg_in_a71 ,jpeg_in_a72 ,jpeg_in_a73 ,jpeg_in_a74 ,jpeg_in_a75 ,
	jpeg_in_a76 ,jpeg_in_a77 ,jpeg_in_a78 ,jpeg_in_a79 ,jpeg_in_a80 ,jpeg_in_a81 ,
	jpeg_in_a82 ,jpeg_in_a83 ,jpeg_in_a84 ,jpeg_in_a85 ,jpeg_in_a86 ,jpeg_in_a87 ,
	jpeg_in_a88 ,jpeg_in_a89 ,jpeg_in_a90 ,jpeg_in_a91 ,jpeg_in_a92 ,jpeg_in_a93 ,
	jpeg_in_a94 ,jpeg_in_a95 ,jpeg_in_a96 ,jpeg_in_a97 ,jpeg_in_a98 ,jpeg_in_a99 ,
	jpeg_in_a100 ,jpeg_in_a101 ,jpeg_in_a102 ,jpeg_in_a103 ,jpeg_in_a104 ,jpeg_in_a105 ,
	jpeg_in_a106 ,jpeg_in_a107 ,jpeg_in_a108 ,jpeg_in_a109 ,jpeg_in_a110 ,jpeg_in_a111 ,
	jpeg_in_a112 ,jpeg_in_a113 ,jpeg_in_a114 ,jpeg_in_a115 ,jpeg_in_a116 ,jpeg_in_a117 ,
	jpeg_in_a118 ,jpeg_in_a119 ,jpeg_in_a120 ,jpeg_in_a121 ,jpeg_in_a122 ,jpeg_in_a123 ,
	jpeg_in_a124 ,jpeg_in_a125 ,jpeg_in_a126 ,jpeg_in_a127 ,jpeg_out_a00 ,jpeg_out_a01 ,
	jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,jpeg_out_a06 ,jpeg_out_a07 ,
	jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,jpeg_out_a12 ,jpeg_out_a13 ,
	jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,jpeg_out_a18 ,jpeg_out_a19 ,
	jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,jpeg_out_a24 ,jpeg_out_a25 ,
	jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,jpeg_out_a30 ,jpeg_out_a31 ,
	jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,jpeg_out_a36 ,jpeg_out_a37 ,
	jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,jpeg_out_a42 ,jpeg_out_a43 ,
	jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,jpeg_out_a48 ,jpeg_out_a49 ,
	jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,jpeg_out_a54 ,jpeg_out_a55 ,
	jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,jpeg_out_a60 ,jpeg_out_a61 ,
	jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,jpeg_out_a66 ,jpeg_out_a67 ,
	jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,jpeg_out_a72 ,jpeg_out_a73 ,
	jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,jpeg_out_a78 ,jpeg_out_a79 ,
	jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,jpeg_out_a84 ,jpeg_out_a85 ,
	jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,jpeg_out_a90 ,jpeg_out_a91 ,
	jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,jpeg_out_a96 ,jpeg_out_a97 ,
	jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,jpeg_out_a102 ,
	jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,jpeg_out_a107 ,
	jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,jpeg_out_a112 ,
	jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,jpeg_out_a117 ,
	jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,jpeg_out_a122 ,
	jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,jpeg_out_a127 ,
	jpeg_len_out ,valid ,ST1_15d ,ST1_14d ,ST1_13d ,ST1_12d ,ST1_11d ,ST1_10d ,
	ST1_09d ,ST1_08d ,ST1_07d ,ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,ST1_02d ,
	ST1_01d ,JF_01_port ,FL01_01_Leos_all ,lop8u_11ot_port ,JF_05 ,FL02_01_Leos_all ,
	JF_08 ,JF_09 ,JF_10 ,FL01_02_01_stall_port );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a64 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a65 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a66 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a67 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a68 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a69 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a70 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a71 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a72 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a73 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a74 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a75 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a76 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a77 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a78 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a79 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a80 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a81 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a82 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a83 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a84 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a85 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a86 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a87 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a88 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a89 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a90 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a91 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a92 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a93 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a94 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a95 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a96 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a97 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a98 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a99 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a100 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a101 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a102 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a103 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a104 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a105 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a106 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a107 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a108 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a109 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a110 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a111 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a112 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a113 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a114 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a115 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a116 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a117 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a118 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a119 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a120 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a121 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a122 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a123 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a124 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a125 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a126 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a127 ;	// line#=../rle.h:56
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
input		ST1_15d ;
input		ST1_14d ;
input		ST1_13d ;
input		ST1_12d ;
input		ST1_11d ;
input		ST1_10d ;
input		ST1_09d ;
input		ST1_08d ;
input		ST1_07d ;
input		ST1_06d ;
input		ST1_05d ;
input		ST1_04d ;
input		ST1_03d ;
input		ST1_02d ;
input		ST1_01d ;
output		JF_01_port ;
output		FL01_01_Leos_all ;
output		lop8u_11ot_port ;
output		JF_05 ;
output		FL02_01_Leos_all ;
output		JF_08 ;
output		JF_09 ;
output		JF_10 ;
output		FL01_02_01_stall_port ;
wire		M_459 ;
wire		M_458 ;
wire		M_457 ;
wire		M_456 ;
wire		M_455 ;
wire		M_454 ;
wire		M_453 ;
wire		M_452 ;
wire		M_450 ;
wire		M_449 ;
wire		M_447 ;
wire		M_445 ;
wire		M_444 ;
wire		M_443 ;
wire		M_442 ;
wire		M_435 ;
wire		M_432 ;
wire		U_165 ;
wire		U_164 ;
wire		U_159 ;
wire		U_147 ;
wire		U_143 ;
wire		U_140 ;
wire		U_139 ;
wire		U_136 ;
wire		U_135 ;
wire		U_132 ;
wire		U_131 ;
wire		U_130 ;
wire		U_129 ;
wire		U_126 ;
wire		U_125 ;
wire		U_123 ;
wire		U_121 ;
wire		U_118 ;
wire		U_117 ;
wire		U_114 ;
wire		U_112 ;
wire		U_111 ;
wire		U_108 ;
wire		U_107 ;
wire		U_105 ;
wire		U_103 ;
wire		U_102 ;
wire		U_99 ;
wire		U_96 ;
wire		U_95 ;
wire		U_94 ;
wire		U_93 ;
wire		U_92 ;
wire		U_91 ;
wire		U_87 ;
wire		U_85 ;
wire		C_12 ;
wire		U_82 ;
wire		U_79 ;
wire		U_77 ;
wire		U_75 ;
wire		U_74 ;
wire		U_73 ;
wire		U_72 ;
wire		U_70 ;
wire		U_69 ;
wire		U_68 ;
wire		U_67 ;
wire		U_61 ;
wire		U_59 ;
wire		U_58 ;
wire		C_08 ;
wire		U_55 ;
wire		U_54 ;
wire		U_51 ;
wire		U_50 ;
wire		U_49 ;
wire		U_48 ;
wire		U_47 ;
wire		C_06 ;
wire		U_46 ;
wire		U_44 ;
wire		U_41 ;
wire		U_40 ;
wire		U_39 ;
wire		U_38 ;
wire		U_37 ;
wire		C_04 ;
wire		U_36 ;
wire		U_35 ;
wire		U_34 ;
wire		U_28 ;
wire		U_25 ;
wire		U_24 ;
wire		U_21 ;
wire		U_20 ;
wire		U_19 ;
wire		U_17 ;
wire		U_15 ;
wire		U_10 ;
wire		U_06 ;
wire		U_05 ;
wire		U_04 ;
wire		C_01 ;
wire		rl_we02 ;	// line#=../rle.cpp:23
wire		rl_we01 ;	// line#=../rle.cpp:23
wire	[127:0]	rl_d02 ;	// line#=../rle.cpp:23
wire	[127:0]	rl_d01 ;	// line#=../rle.cpp:23
wire	[6:0]	rl_ad02 ;	// line#=../rle.cpp:23
wire	[6:0]	rl_ad01 ;	// line#=../rle.cpp:23
wire	[63:0]	quantized_block_d01 ;	// line#=../rle.cpp:22
wire	[5:0]	quantized_block_ad01 ;	// line#=../rle.cpp:22
wire	[5:0]	incr8u_61i1 ;
wire	[5:0]	incr8u_61ot ;
wire	[5:0]	incr8u_71i1 ;
wire	[6:0]	incr8u_71ot ;
wire	[31:0]	decr32s2i1 ;
wire	[31:0]	decr32s2ot ;
wire	[31:0]	decr32s1i1 ;
wire	[31:0]	decr32s1ot ;
wire	[6:0]	decr8u_71i1 ;
wire	[6:0]	decr8u_71ot ;
wire	[31:0]	incr32s3i1 ;
wire	[31:0]	incr32s3ot ;
wire	[31:0]	incr32s2i1 ;
wire	[31:0]	incr32s2ot ;
wire	[31:0]	incr32s1i1 ;
wire	[31:0]	incr32s1ot ;
wire	[7:0]	incr8u2i1 ;
wire	[7:0]	incr8u2ot ;
wire	[7:0]	incr8u1i1 ;
wire	[7:0]	incr8u1ot ;
wire	[3:0]	incr4s1ot ;
wire	[2:0]	incr3u1i1 ;
wire	[3:0]	incr3u1ot ;
wire	[5:0]	lop8u_11i2 ;
wire	[5:0]	lop8u_11i1 ;
wire		lop8u_11ot ;
wire	[8:0]	sub12s_91i2 ;
wire	[8:0]	sub12s_91i1 ;
wire	[8:0]	sub12s_91ot ;
wire	[7:0]	sub8u1i1 ;
wire	[7:0]	sub8u1ot ;
wire		add3u1i2 ;
wire	[2:0]	add3u1i1 ;
wire	[3:0]	add3u1ot ;
wire		FL02_05_ndat ;
wire		FL02_04_ndat ;
wire		FL02_04_rdy ;
wire		FL02_02_Lndat ;
wire		FL02_02_Lrdy ;
wire		FL02_02_ndat ;
wire		FL02_02_rdy ;
wire		FL02_01_ndat ;
wire		FL02_05_ngo ;
wire		FL02_06_eos ;
wire		FL02_05_eos ;
wire		FL02_04_eos ;
wire		FL02_03_eos ;
wire		FL02_02_eos ;
wire		FL02_01_eos ;
wire		FL02_02_Leos_all ;
wire		FL02_02_Leos ;
wire		FL02_01_Leos_all ;
wire		FJ_11_12 ;
wire		FJ_09_15 ;
wire		FL02_06_01a ;
wire		FL02_05_01a ;
wire		FL02_04_01a ;
wire		FL02_03_01a ;
wire		FL02_02_01a ;
wire		FL02_01_01a ;
wire		FL02_03_break ;
wire		FL02_02_break ;
wire		FL02_01_break ;
wire		FL01_01_ndat ;
wire		FL01_02_01_stall ;
wire		FL01_02_eos ;
wire		FL01_01_eos ;
wire		FL01_01_Leos_all ;
wire		FJ_04_04 ;
wire		FJ_03_05 ;
wire		FL01_02_01a ;
wire		FL01_01_01a ;
wire		FL01_01_break ;
wire		JF_10 ;
wire		JF_09 ;
wire		CT_17 ;
wire		CT_16 ;
wire		CT_14 ;
wire		CT_11 ;
wire		JF_05 ;
wire		CT_06 ;
wire		JF_01 ;
wire		CMPS_FL_C2496_1_DO_v ;
wire		zz_WE2 ;
wire	[8:0]	CMPS_FL_C2603_1_DO_t ;
wire	[8:0]	CMPS_FL_C2496_1_DO_t ;
wire	[8:0]	zz_RD1 ;
wire		RG_previous_dc_en ;
wire		RG_03_02_en ;
wire		FF_j_en ;
wire		RG_i_03_en ;
wire		RG_k_03_en ;
wire		RG_i_02_en ;
wire		RG_k_02_en ;
wire		RG_i_04_en ;
wire		RG_k_04_en ;
wire		RG_i_05_en ;
wire		jpeg_out_a00_r_en ;
wire		jpeg_out_a01_r_en ;
wire		jpeg_out_a02_r_en ;
wire		jpeg_out_a03_r_en ;
wire		jpeg_out_a04_r_en ;
wire		jpeg_out_a05_r_en ;
wire		jpeg_out_a06_r_en ;
wire		jpeg_out_a07_r_en ;
wire		jpeg_out_a08_r_en ;
wire		jpeg_out_a09_r_en ;
wire		jpeg_out_a10_r_en ;
wire		jpeg_out_a11_r_en ;
wire		jpeg_out_a12_r_en ;
wire		jpeg_out_a13_r_en ;
wire		jpeg_out_a14_r_en ;
wire		jpeg_out_a15_r_en ;
wire		jpeg_out_a16_r_en ;
wire		jpeg_out_a17_r_en ;
wire		jpeg_out_a18_r_en ;
wire		jpeg_out_a19_r_en ;
wire		jpeg_out_a20_r_en ;
wire		jpeg_out_a21_r_en ;
wire		jpeg_out_a22_r_en ;
wire		jpeg_out_a23_r_en ;
wire		jpeg_out_a24_r_en ;
wire		jpeg_out_a25_r_en ;
wire		jpeg_out_a26_r_en ;
wire		jpeg_out_a27_r_en ;
wire		jpeg_out_a28_r_en ;
wire		jpeg_out_a29_r_en ;
wire		jpeg_out_a30_r_en ;
wire		jpeg_out_a31_r_en ;
wire		jpeg_out_a32_r_en ;
wire		jpeg_out_a33_r_en ;
wire		jpeg_out_a34_r_en ;
wire		jpeg_out_a35_r_en ;
wire		jpeg_out_a36_r_en ;
wire		jpeg_out_a37_r_en ;
wire		jpeg_out_a38_r_en ;
wire		jpeg_out_a39_r_en ;
wire		jpeg_out_a40_r_en ;
wire		jpeg_out_a41_r_en ;
wire		jpeg_out_a42_r_en ;
wire		jpeg_out_a43_r_en ;
wire		jpeg_out_a44_r_en ;
wire		jpeg_out_a45_r_en ;
wire		jpeg_out_a46_r_en ;
wire		jpeg_out_a47_r_en ;
wire		jpeg_out_a48_r_en ;
wire		jpeg_out_a49_r_en ;
wire		jpeg_out_a50_r_en ;
wire		jpeg_out_a51_r_en ;
wire		jpeg_out_a52_r_en ;
wire		jpeg_out_a53_r_en ;
wire		jpeg_out_a54_r_en ;
wire		jpeg_out_a55_r_en ;
wire		jpeg_out_a56_r_en ;
wire		jpeg_out_a57_r_en ;
wire		jpeg_out_a58_r_en ;
wire		jpeg_out_a59_r_en ;
wire		jpeg_out_a60_r_en ;
wire		jpeg_out_a61_r_en ;
wire		jpeg_out_a62_r_en ;
wire		jpeg_out_a63_r_en ;
wire		jpeg_out_a64_r_en ;
wire		jpeg_out_a65_r_en ;
wire		jpeg_out_a66_r_en ;
wire		jpeg_out_a67_r_en ;
wire		jpeg_out_a68_r_en ;
wire		jpeg_out_a69_r_en ;
wire		jpeg_out_a70_r_en ;
wire		jpeg_out_a71_r_en ;
wire		jpeg_out_a72_r_en ;
wire		jpeg_out_a73_r_en ;
wire		jpeg_out_a74_r_en ;
wire		jpeg_out_a75_r_en ;
wire		jpeg_out_a76_r_en ;
wire		jpeg_out_a77_r_en ;
wire		jpeg_out_a78_r_en ;
wire		jpeg_out_a79_r_en ;
wire		jpeg_out_a80_r_en ;
wire		jpeg_out_a81_r_en ;
wire		jpeg_out_a82_r_en ;
wire		jpeg_out_a83_r_en ;
wire		jpeg_out_a84_r_en ;
wire		jpeg_out_a85_r_en ;
wire		jpeg_out_a86_r_en ;
wire		jpeg_out_a87_r_en ;
wire		jpeg_out_a88_r_en ;
wire		jpeg_out_a89_r_en ;
wire		jpeg_out_a90_r_en ;
wire		jpeg_out_a91_r_en ;
wire		jpeg_out_a92_r_en ;
wire		jpeg_out_a93_r_en ;
wire		jpeg_out_a94_r_en ;
wire		jpeg_out_a95_r_en ;
wire		jpeg_out_a96_r_en ;
wire		jpeg_out_a97_r_en ;
wire		jpeg_out_a98_r_en ;
wire		jpeg_out_a99_r_en ;
wire		jpeg_out_a100_r_en ;
wire		jpeg_out_a101_r_en ;
wire		jpeg_out_a102_r_en ;
wire		jpeg_out_a103_r_en ;
wire		jpeg_out_a104_r_en ;
wire		jpeg_out_a105_r_en ;
wire		jpeg_out_a106_r_en ;
wire		jpeg_out_a107_r_en ;
wire		jpeg_out_a108_r_en ;
wire		jpeg_out_a109_r_en ;
wire		jpeg_out_a110_r_en ;
wire		jpeg_out_a111_r_en ;
wire		jpeg_out_a112_r_en ;
wire		jpeg_out_a113_r_en ;
wire		jpeg_out_a114_r_en ;
wire		jpeg_out_a115_r_en ;
wire		jpeg_out_a116_r_en ;
wire		jpeg_out_a117_r_en ;
wire		jpeg_out_a118_r_en ;
wire		jpeg_out_a119_r_en ;
wire		jpeg_out_a120_r_en ;
wire		jpeg_out_a121_r_en ;
wire		jpeg_out_a122_r_en ;
wire		jpeg_out_a123_r_en ;
wire		jpeg_out_a124_r_en ;
wire		jpeg_out_a125_r_en ;
wire		jpeg_out_a126_r_en ;
wire		jpeg_out_a127_r_en ;
wire		jpeg_len_out_r_en ;
wire		quantized_block_rg00_en ;
wire		quantized_block_rg01_en ;
wire		quantized_block_rg02_en ;
wire		quantized_block_rg03_en ;
wire		quantized_block_rg04_en ;
wire		quantized_block_rg05_en ;
wire		quantized_block_rg06_en ;
wire		quantized_block_rg07_en ;
wire		quantized_block_rg08_en ;
wire		quantized_block_rg09_en ;
wire		quantized_block_rg10_en ;
wire		quantized_block_rg11_en ;
wire		quantized_block_rg12_en ;
wire		quantized_block_rg13_en ;
wire		quantized_block_rg14_en ;
wire		quantized_block_rg15_en ;
wire		quantized_block_rg16_en ;
wire		quantized_block_rg17_en ;
wire		quantized_block_rg18_en ;
wire		quantized_block_rg19_en ;
wire		quantized_block_rg20_en ;
wire		quantized_block_rg21_en ;
wire		quantized_block_rg22_en ;
wire		quantized_block_rg23_en ;
wire		quantized_block_rg24_en ;
wire		quantized_block_rg25_en ;
wire		quantized_block_rg26_en ;
wire		quantized_block_rg27_en ;
wire		quantized_block_rg28_en ;
wire		quantized_block_rg29_en ;
wire		quantized_block_rg30_en ;
wire		quantized_block_rg31_en ;
wire		quantized_block_rg32_en ;
wire		quantized_block_rg33_en ;
wire		quantized_block_rg34_en ;
wire		quantized_block_rg35_en ;
wire		quantized_block_rg36_en ;
wire		quantized_block_rg37_en ;
wire		quantized_block_rg38_en ;
wire		quantized_block_rg39_en ;
wire		quantized_block_rg40_en ;
wire		quantized_block_rg41_en ;
wire		quantized_block_rg42_en ;
wire		quantized_block_rg43_en ;
wire		quantized_block_rg44_en ;
wire		quantized_block_rg45_en ;
wire		quantized_block_rg46_en ;
wire		quantized_block_rg47_en ;
wire		quantized_block_rg48_en ;
wire		quantized_block_rg49_en ;
wire		quantized_block_rg50_en ;
wire		quantized_block_rg51_en ;
wire		quantized_block_rg52_en ;
wire		quantized_block_rg53_en ;
wire		quantized_block_rg54_en ;
wire		quantized_block_rg55_en ;
wire		quantized_block_rg56_en ;
wire		quantized_block_rg57_en ;
wire		quantized_block_rg58_en ;
wire		quantized_block_rg59_en ;
wire		quantized_block_rg60_en ;
wire		quantized_block_rg61_en ;
wire		quantized_block_rg62_en ;
wire		quantized_block_rg63_en ;
wire		M_01 ;
wire		rl_rg00_en ;
wire		rl_rg01_en ;
wire		rl_rg02_en ;
wire		rl_rg03_en ;
wire		rl_rg04_en ;
wire		rl_rg05_en ;
wire		rl_rg06_en ;
wire		rl_rg07_en ;
wire		rl_rg08_en ;
wire		rl_rg09_en ;
wire		rl_rg10_en ;
wire		rl_rg11_en ;
wire		rl_rg12_en ;
wire		rl_rg13_en ;
wire		rl_rg14_en ;
wire		rl_rg15_en ;
wire		rl_rg16_en ;
wire		rl_rg17_en ;
wire		rl_rg18_en ;
wire		rl_rg19_en ;
wire		rl_rg20_en ;
wire		rl_rg21_en ;
wire		rl_rg22_en ;
wire		rl_rg23_en ;
wire		rl_rg24_en ;
wire		rl_rg25_en ;
wire		rl_rg26_en ;
wire		rl_rg27_en ;
wire		rl_rg28_en ;
wire		rl_rg29_en ;
wire		rl_rg30_en ;
wire		rl_rg31_en ;
wire		rl_rg32_en ;
wire		rl_rg33_en ;
wire		rl_rg34_en ;
wire		rl_rg35_en ;
wire		rl_rg36_en ;
wire		rl_rg37_en ;
wire		rl_rg38_en ;
wire		rl_rg39_en ;
wire		rl_rg40_en ;
wire		rl_rg41_en ;
wire		rl_rg42_en ;
wire		rl_rg43_en ;
wire		rl_rg44_en ;
wire		rl_rg45_en ;
wire		rl_rg46_en ;
wire		rl_rg47_en ;
wire		rl_rg48_en ;
wire		rl_rg49_en ;
wire		rl_rg50_en ;
wire		rl_rg51_en ;
wire		rl_rg52_en ;
wire		rl_rg53_en ;
wire		rl_rg54_en ;
wire		rl_rg55_en ;
wire		rl_rg56_en ;
wire		rl_rg57_en ;
wire		rl_rg58_en ;
wire		rl_rg59_en ;
wire		rl_rg60_en ;
wire		rl_rg61_en ;
wire		rl_rg62_en ;
wire		rl_rg63_en ;
wire		rl_rg64_en ;
wire		rl_rg65_en ;
wire		rl_rg66_en ;
wire		rl_rg67_en ;
wire		rl_rg68_en ;
wire		rl_rg69_en ;
wire		rl_rg70_en ;
wire		rl_rg71_en ;
wire		rl_rg72_en ;
wire		rl_rg73_en ;
wire		rl_rg74_en ;
wire		rl_rg75_en ;
wire		rl_rg76_en ;
wire		rl_rg77_en ;
wire		rl_rg78_en ;
wire		rl_rg79_en ;
wire		rl_rg80_en ;
wire		rl_rg81_en ;
wire		rl_rg82_en ;
wire		rl_rg83_en ;
wire		rl_rg84_en ;
wire		rl_rg85_en ;
wire		rl_rg86_en ;
wire		rl_rg87_en ;
wire		rl_rg88_en ;
wire		rl_rg89_en ;
wire		rl_rg90_en ;
wire		rl_rg91_en ;
wire		rl_rg92_en ;
wire		rl_rg93_en ;
wire		rl_rg94_en ;
wire		rl_rg95_en ;
wire		rl_rg96_en ;
wire		rl_rg97_en ;
wire		rl_rg98_en ;
wire		rl_rg99_en ;
wire		rl_rg100_en ;
wire		rl_rg101_en ;
wire		rl_rg102_en ;
wire		rl_rg103_en ;
wire		rl_rg104_en ;
wire		rl_rg105_en ;
wire		rl_rg106_en ;
wire		rl_rg107_en ;
wire		rl_rg108_en ;
wire		rl_rg109_en ;
wire		rl_rg110_en ;
wire		rl_rg111_en ;
wire		rl_rg112_en ;
wire		rl_rg113_en ;
wire		rl_rg114_en ;
wire		rl_rg115_en ;
wire		rl_rg116_en ;
wire		rl_rg117_en ;
wire		rl_rg118_en ;
wire		rl_rg119_en ;
wire		rl_rg120_en ;
wire		rl_rg121_en ;
wire		rl_rg122_en ;
wire		rl_rg123_en ;
wire		rl_rg124_en ;
wire		rl_rg125_en ;
wire		rl_rg126_en ;
wire		rl_rg127_en ;
wire		RG_y_02_en ;
wire		RG_j_x_02_en ;
wire		RG_i_06_en ;
wire		RG_len_05_en ;
wire		RG_i_en ;
wire		RG_j_k_en ;
wire		FF_d_05_en ;
wire		RG_15_02_en ;
wire		RG_k_05_en ;
wire		FL01_01_streg_en ;
wire		FL01_02_streg_en ;
wire		flag_r1_en ;
wire		flag_r2_en ;
wire		flag_r3_en ;
wire		FL02_01_streg_en ;
wire		FL02_02_streg_en ;
wire		FL02_03_streg_en ;
wire		FL02_04_streg_en ;
wire		FL02_05_streg_en ;
wire		FL02_06_streg_en ;
wire		valid_r_en ;
reg	[8:0]	rl_rg127 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg126 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg125 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg124 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg123 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg122 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg121 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg120 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg119 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg118 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg117 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg116 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg115 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg114 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg113 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg112 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg111 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg110 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg109 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg108 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg107 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg106 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg105 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg104 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg103 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg102 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg101 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg100 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg99 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg98 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg97 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg96 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg95 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg94 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg93 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg92 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg91 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg90 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg89 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg88 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg87 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg86 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg85 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg84 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg83 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg82 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg81 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg80 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg79 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg78 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg77 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg76 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg75 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg74 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg73 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg72 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg71 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg70 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg69 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg68 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg67 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg66 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg65 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg64 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg63 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg62 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg61 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg60 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg59 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg58 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg57 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg56 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg55 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg54 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg53 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg52 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg51 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg50 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg49 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg48 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg47 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg46 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg45 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg44 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg43 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg42 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg41 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg40 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg39 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg38 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg37 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg36 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg35 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg34 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg33 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg32 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg31 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg30 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg29 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg28 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg27 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg26 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg25 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg24 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg23 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg22 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg21 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg20 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg19 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg18 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg17 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg16 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg15 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg14 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg13 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg12 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg11 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg10 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg09 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg08 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg07 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg06 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg05 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg04 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg03 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg02 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg01 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg00 ;	// line#=../rle.cpp:23
reg	[8:0]	quantized_block_rg63 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg62 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg61 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg60 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg59 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg58 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg57 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg56 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg55 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg54 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg53 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg52 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg51 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg50 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg49 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg48 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg47 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg46 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg45 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg44 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg43 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg42 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg41 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg40 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg39 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg38 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg37 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg36 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg35 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg34 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg33 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg32 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg31 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg30 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg29 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg28 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg27 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg26 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg25 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg24 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg23 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg22 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg21 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg20 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg19 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg18 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg17 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg16 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg15 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg14 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg13 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg12 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg11 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg10 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg09 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg08 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg07 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg06 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg05 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg04 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg03 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg02 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg01 ;	// line#=../rle.cpp:22
reg	[8:0]	quantized_block_rg00 ;	// line#=../rle.cpp:22
reg	FL02_06_streg ;
reg	FL02_05_streg ;
reg	FL02_04_streg ;
reg	FL02_03_streg ;
reg	[1:0]	FL02_02_streg ;
reg	[1:0]	FL02_01_streg ;
reg	flag_r3 ;
reg	flag_r2 ;
reg	flag_r1 ;
reg	FL01_02_streg ;
reg	FL01_01_streg ;
reg	[8:0]	RG_previous_dc ;	// line#=../rle.h:66
reg	[3:0]	RG_y_02 ;	// line#=../rle.cpp:25
reg	[3:0]	RG_j_x_02 ;	// line#=../rle.cpp:25,27
reg	[2:0]	RG_03_02 ;
reg	[31:0]	RG_i_06 ;	// line#=../rle.cpp:25
reg	[7:0]	RG_len_05 ;	// line#=../rle.cpp:24
reg	FF_j ;	// line#=../rle.cpp:27
reg	[31:0]	RG_i_03 ;	// line#=../rle.cpp:25
reg	[8:0]	RG_k_03 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_i ;	// line#=../rle.cpp:25,105
reg	[31:0]	RG_j_k ;	// line#=../rle.cpp:25,105
reg	[5:0]	RG_k ;	// line#=../rle.cpp:105
reg	FF_d_05 ;	// line#=../rle.cpp:105
reg	[31:0]	RG_i_02 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_k_02 ;	// line#=../rle.cpp:25
reg	RG_15_02 ;
reg	[6:0]	RG_k_05 ;	// line#=../rle.cpp:105
reg	[31:0]	RG_i_04 ;	// line#=../rle.cpp:25
reg	[8:0]	RG_k_04 ;	// line#=../rle.cpp:25
reg	[31:0]	RG_i_05 ;	// line#=../rle.cpp:25
reg	[8:0]	jpeg_out_a00_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a01_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a02_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a03_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a04_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a05_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a06_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a07_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a08_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a09_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a10_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a11_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a12_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a13_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a14_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a15_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a16_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a17_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a18_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a19_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a20_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a21_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a22_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a23_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a24_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a25_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a26_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a27_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a28_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a29_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a30_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a31_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a32_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a33_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a34_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a35_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a36_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a37_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a38_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a39_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a40_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a41_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a42_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a43_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a44_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a45_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a46_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a47_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a48_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a49_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a50_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a51_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a52_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a53_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a54_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a55_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a56_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a57_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a58_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a59_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a60_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a61_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a62_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a63_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a64_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a65_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a66_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a67_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a68_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a69_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a70_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a71_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a72_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a73_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a74_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a75_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a76_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a77_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a78_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a79_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a80_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a81_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a82_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a83_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a84_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a85_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a86_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a87_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a88_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a89_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a90_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a91_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a92_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a93_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a94_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a95_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a96_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a97_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a98_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a99_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a100_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a101_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a102_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a103_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a104_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a105_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a106_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a107_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a108_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a109_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a110_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a111_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a112_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a113_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a114_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a115_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a116_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a117_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a118_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a119_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a120_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a121_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a122_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a123_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a124_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a125_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a126_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a127_r ;	// line#=../rle.h:60
reg	[11:0]	jpeg_len_out_r ;	// line#=../rle.h:61
reg	valid_r ;	// line#=../rle.h:62
reg	FA02_02_gnt ;
reg	FA02_03_gnt ;
reg	[8:0]	quantized_block_rd00 ;	// line#=../rle.cpp:22
reg	[8:0]	rl_rd00 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_rg00_t ;
reg	rl_rg00_t_c1 ;
reg	rl_rg00_t_c2 ;
reg	rl_rg00_t_c3 ;
reg	[8:0]	rl_rg01_t ;
reg	rl_rg01_t_c1 ;
reg	rl_rg01_t_c2 ;
reg	[8:0]	rl_rg02_t ;
reg	rl_rg02_t_c1 ;
reg	rl_rg02_t_c2 ;
reg	[8:0]	rl_rg03_t ;
reg	rl_rg03_t_c1 ;
reg	rl_rg03_t_c2 ;
reg	[8:0]	rl_rg04_t ;
reg	rl_rg04_t_c1 ;
reg	rl_rg04_t_c2 ;
reg	[8:0]	rl_rg05_t ;
reg	rl_rg05_t_c1 ;
reg	rl_rg05_t_c2 ;
reg	[8:0]	rl_rg06_t ;
reg	rl_rg06_t_c1 ;
reg	rl_rg06_t_c2 ;
reg	[8:0]	rl_rg07_t ;
reg	rl_rg07_t_c1 ;
reg	rl_rg07_t_c2 ;
reg	[8:0]	rl_rg08_t ;
reg	rl_rg08_t_c1 ;
reg	rl_rg08_t_c2 ;
reg	[8:0]	rl_rg09_t ;
reg	rl_rg09_t_c1 ;
reg	rl_rg09_t_c2 ;
reg	[8:0]	rl_rg10_t ;
reg	rl_rg10_t_c1 ;
reg	rl_rg10_t_c2 ;
reg	[8:0]	rl_rg11_t ;
reg	rl_rg11_t_c1 ;
reg	rl_rg11_t_c2 ;
reg	[8:0]	rl_rg12_t ;
reg	rl_rg12_t_c1 ;
reg	rl_rg12_t_c2 ;
reg	[8:0]	rl_rg13_t ;
reg	rl_rg13_t_c1 ;
reg	rl_rg13_t_c2 ;
reg	[8:0]	rl_rg14_t ;
reg	rl_rg14_t_c1 ;
reg	rl_rg14_t_c2 ;
reg	[8:0]	rl_rg15_t ;
reg	rl_rg15_t_c1 ;
reg	rl_rg15_t_c2 ;
reg	[8:0]	rl_rg16_t ;
reg	rl_rg16_t_c1 ;
reg	rl_rg16_t_c2 ;
reg	[8:0]	rl_rg17_t ;
reg	rl_rg17_t_c1 ;
reg	rl_rg17_t_c2 ;
reg	[8:0]	rl_rg18_t ;
reg	rl_rg18_t_c1 ;
reg	rl_rg18_t_c2 ;
reg	[8:0]	rl_rg19_t ;
reg	rl_rg19_t_c1 ;
reg	rl_rg19_t_c2 ;
reg	[8:0]	rl_rg20_t ;
reg	rl_rg20_t_c1 ;
reg	rl_rg20_t_c2 ;
reg	[8:0]	rl_rg21_t ;
reg	rl_rg21_t_c1 ;
reg	rl_rg21_t_c2 ;
reg	[8:0]	rl_rg22_t ;
reg	rl_rg22_t_c1 ;
reg	rl_rg22_t_c2 ;
reg	[8:0]	rl_rg23_t ;
reg	rl_rg23_t_c1 ;
reg	rl_rg23_t_c2 ;
reg	[8:0]	rl_rg24_t ;
reg	rl_rg24_t_c1 ;
reg	rl_rg24_t_c2 ;
reg	[8:0]	rl_rg25_t ;
reg	rl_rg25_t_c1 ;
reg	rl_rg25_t_c2 ;
reg	[8:0]	rl_rg26_t ;
reg	rl_rg26_t_c1 ;
reg	rl_rg26_t_c2 ;
reg	[8:0]	rl_rg27_t ;
reg	rl_rg27_t_c1 ;
reg	rl_rg27_t_c2 ;
reg	[8:0]	rl_rg28_t ;
reg	rl_rg28_t_c1 ;
reg	rl_rg28_t_c2 ;
reg	[8:0]	rl_rg29_t ;
reg	rl_rg29_t_c1 ;
reg	rl_rg29_t_c2 ;
reg	[8:0]	rl_rg30_t ;
reg	rl_rg30_t_c1 ;
reg	rl_rg30_t_c2 ;
reg	[8:0]	rl_rg31_t ;
reg	rl_rg31_t_c1 ;
reg	rl_rg31_t_c2 ;
reg	[8:0]	rl_rg32_t ;
reg	rl_rg32_t_c1 ;
reg	rl_rg32_t_c2 ;
reg	[8:0]	rl_rg33_t ;
reg	rl_rg33_t_c1 ;
reg	rl_rg33_t_c2 ;
reg	[8:0]	rl_rg34_t ;
reg	rl_rg34_t_c1 ;
reg	rl_rg34_t_c2 ;
reg	[8:0]	rl_rg35_t ;
reg	rl_rg35_t_c1 ;
reg	rl_rg35_t_c2 ;
reg	[8:0]	rl_rg36_t ;
reg	rl_rg36_t_c1 ;
reg	rl_rg36_t_c2 ;
reg	[8:0]	rl_rg37_t ;
reg	rl_rg37_t_c1 ;
reg	rl_rg37_t_c2 ;
reg	[8:0]	rl_rg38_t ;
reg	rl_rg38_t_c1 ;
reg	rl_rg38_t_c2 ;
reg	[8:0]	rl_rg39_t ;
reg	rl_rg39_t_c1 ;
reg	rl_rg39_t_c2 ;
reg	[8:0]	rl_rg40_t ;
reg	rl_rg40_t_c1 ;
reg	rl_rg40_t_c2 ;
reg	[8:0]	rl_rg41_t ;
reg	rl_rg41_t_c1 ;
reg	rl_rg41_t_c2 ;
reg	[8:0]	rl_rg42_t ;
reg	rl_rg42_t_c1 ;
reg	rl_rg42_t_c2 ;
reg	[8:0]	rl_rg43_t ;
reg	rl_rg43_t_c1 ;
reg	rl_rg43_t_c2 ;
reg	[8:0]	rl_rg44_t ;
reg	rl_rg44_t_c1 ;
reg	rl_rg44_t_c2 ;
reg	[8:0]	rl_rg45_t ;
reg	rl_rg45_t_c1 ;
reg	rl_rg45_t_c2 ;
reg	[8:0]	rl_rg46_t ;
reg	rl_rg46_t_c1 ;
reg	rl_rg46_t_c2 ;
reg	[8:0]	rl_rg47_t ;
reg	rl_rg47_t_c1 ;
reg	rl_rg47_t_c2 ;
reg	[8:0]	rl_rg48_t ;
reg	rl_rg48_t_c1 ;
reg	rl_rg48_t_c2 ;
reg	[8:0]	rl_rg49_t ;
reg	rl_rg49_t_c1 ;
reg	rl_rg49_t_c2 ;
reg	[8:0]	rl_rg50_t ;
reg	rl_rg50_t_c1 ;
reg	rl_rg50_t_c2 ;
reg	[8:0]	rl_rg51_t ;
reg	rl_rg51_t_c1 ;
reg	rl_rg51_t_c2 ;
reg	[8:0]	rl_rg52_t ;
reg	rl_rg52_t_c1 ;
reg	rl_rg52_t_c2 ;
reg	[8:0]	rl_rg53_t ;
reg	rl_rg53_t_c1 ;
reg	rl_rg53_t_c2 ;
reg	[8:0]	rl_rg54_t ;
reg	rl_rg54_t_c1 ;
reg	rl_rg54_t_c2 ;
reg	[8:0]	rl_rg55_t ;
reg	rl_rg55_t_c1 ;
reg	rl_rg55_t_c2 ;
reg	[8:0]	rl_rg56_t ;
reg	rl_rg56_t_c1 ;
reg	rl_rg56_t_c2 ;
reg	[8:0]	rl_rg57_t ;
reg	rl_rg57_t_c1 ;
reg	rl_rg57_t_c2 ;
reg	[8:0]	rl_rg58_t ;
reg	rl_rg58_t_c1 ;
reg	rl_rg58_t_c2 ;
reg	[8:0]	rl_rg59_t ;
reg	rl_rg59_t_c1 ;
reg	rl_rg59_t_c2 ;
reg	[8:0]	rl_rg60_t ;
reg	rl_rg60_t_c1 ;
reg	rl_rg60_t_c2 ;
reg	[8:0]	rl_rg61_t ;
reg	rl_rg61_t_c1 ;
reg	rl_rg61_t_c2 ;
reg	[8:0]	rl_rg62_t ;
reg	rl_rg62_t_c1 ;
reg	rl_rg62_t_c2 ;
reg	[8:0]	rl_rg63_t ;
reg	rl_rg63_t_c1 ;
reg	rl_rg63_t_c2 ;
reg	[8:0]	rl_rg64_t ;
reg	rl_rg64_t_c1 ;
reg	rl_rg64_t_c2 ;
reg	[8:0]	rl_rg65_t ;
reg	rl_rg65_t_c1 ;
reg	rl_rg65_t_c2 ;
reg	[8:0]	rl_rg66_t ;
reg	rl_rg66_t_c1 ;
reg	rl_rg66_t_c2 ;
reg	[8:0]	rl_rg67_t ;
reg	rl_rg67_t_c1 ;
reg	rl_rg67_t_c2 ;
reg	[8:0]	rl_rg68_t ;
reg	rl_rg68_t_c1 ;
reg	rl_rg68_t_c2 ;
reg	[8:0]	rl_rg69_t ;
reg	rl_rg69_t_c1 ;
reg	rl_rg69_t_c2 ;
reg	[8:0]	rl_rg70_t ;
reg	rl_rg70_t_c1 ;
reg	rl_rg70_t_c2 ;
reg	[8:0]	rl_rg71_t ;
reg	rl_rg71_t_c1 ;
reg	rl_rg71_t_c2 ;
reg	[8:0]	rl_rg72_t ;
reg	rl_rg72_t_c1 ;
reg	rl_rg72_t_c2 ;
reg	[8:0]	rl_rg73_t ;
reg	rl_rg73_t_c1 ;
reg	rl_rg73_t_c2 ;
reg	[8:0]	rl_rg74_t ;
reg	rl_rg74_t_c1 ;
reg	rl_rg74_t_c2 ;
reg	[8:0]	rl_rg75_t ;
reg	rl_rg75_t_c1 ;
reg	rl_rg75_t_c2 ;
reg	[8:0]	rl_rg76_t ;
reg	rl_rg76_t_c1 ;
reg	rl_rg76_t_c2 ;
reg	[8:0]	rl_rg77_t ;
reg	rl_rg77_t_c1 ;
reg	rl_rg77_t_c2 ;
reg	[8:0]	rl_rg78_t ;
reg	rl_rg78_t_c1 ;
reg	rl_rg78_t_c2 ;
reg	[8:0]	rl_rg79_t ;
reg	rl_rg79_t_c1 ;
reg	rl_rg79_t_c2 ;
reg	[8:0]	rl_rg80_t ;
reg	rl_rg80_t_c1 ;
reg	rl_rg80_t_c2 ;
reg	[8:0]	rl_rg81_t ;
reg	rl_rg81_t_c1 ;
reg	rl_rg81_t_c2 ;
reg	[8:0]	rl_rg82_t ;
reg	rl_rg82_t_c1 ;
reg	rl_rg82_t_c2 ;
reg	[8:0]	rl_rg83_t ;
reg	rl_rg83_t_c1 ;
reg	rl_rg83_t_c2 ;
reg	[8:0]	rl_rg84_t ;
reg	rl_rg84_t_c1 ;
reg	rl_rg84_t_c2 ;
reg	[8:0]	rl_rg85_t ;
reg	rl_rg85_t_c1 ;
reg	rl_rg85_t_c2 ;
reg	[8:0]	rl_rg86_t ;
reg	rl_rg86_t_c1 ;
reg	rl_rg86_t_c2 ;
reg	[8:0]	rl_rg87_t ;
reg	rl_rg87_t_c1 ;
reg	rl_rg87_t_c2 ;
reg	[8:0]	rl_rg88_t ;
reg	rl_rg88_t_c1 ;
reg	rl_rg88_t_c2 ;
reg	[8:0]	rl_rg89_t ;
reg	rl_rg89_t_c1 ;
reg	rl_rg89_t_c2 ;
reg	[8:0]	rl_rg90_t ;
reg	rl_rg90_t_c1 ;
reg	rl_rg90_t_c2 ;
reg	[8:0]	rl_rg91_t ;
reg	rl_rg91_t_c1 ;
reg	rl_rg91_t_c2 ;
reg	[8:0]	rl_rg92_t ;
reg	rl_rg92_t_c1 ;
reg	rl_rg92_t_c2 ;
reg	[8:0]	rl_rg93_t ;
reg	rl_rg93_t_c1 ;
reg	rl_rg93_t_c2 ;
reg	[8:0]	rl_rg94_t ;
reg	rl_rg94_t_c1 ;
reg	rl_rg94_t_c2 ;
reg	[8:0]	rl_rg95_t ;
reg	rl_rg95_t_c1 ;
reg	rl_rg95_t_c2 ;
reg	[8:0]	rl_rg96_t ;
reg	rl_rg96_t_c1 ;
reg	rl_rg96_t_c2 ;
reg	[8:0]	rl_rg97_t ;
reg	rl_rg97_t_c1 ;
reg	rl_rg97_t_c2 ;
reg	[8:0]	rl_rg98_t ;
reg	rl_rg98_t_c1 ;
reg	rl_rg98_t_c2 ;
reg	[8:0]	rl_rg99_t ;
reg	rl_rg99_t_c1 ;
reg	rl_rg99_t_c2 ;
reg	[8:0]	rl_rg100_t ;
reg	rl_rg100_t_c1 ;
reg	rl_rg100_t_c2 ;
reg	[8:0]	rl_rg101_t ;
reg	rl_rg101_t_c1 ;
reg	rl_rg101_t_c2 ;
reg	[8:0]	rl_rg102_t ;
reg	rl_rg102_t_c1 ;
reg	rl_rg102_t_c2 ;
reg	[8:0]	rl_rg103_t ;
reg	rl_rg103_t_c1 ;
reg	rl_rg103_t_c2 ;
reg	[8:0]	rl_rg104_t ;
reg	rl_rg104_t_c1 ;
reg	rl_rg104_t_c2 ;
reg	[8:0]	rl_rg105_t ;
reg	rl_rg105_t_c1 ;
reg	rl_rg105_t_c2 ;
reg	[8:0]	rl_rg106_t ;
reg	rl_rg106_t_c1 ;
reg	rl_rg106_t_c2 ;
reg	[8:0]	rl_rg107_t ;
reg	rl_rg107_t_c1 ;
reg	rl_rg107_t_c2 ;
reg	[8:0]	rl_rg108_t ;
reg	rl_rg108_t_c1 ;
reg	rl_rg108_t_c2 ;
reg	[8:0]	rl_rg109_t ;
reg	rl_rg109_t_c1 ;
reg	rl_rg109_t_c2 ;
reg	[8:0]	rl_rg110_t ;
reg	rl_rg110_t_c1 ;
reg	rl_rg110_t_c2 ;
reg	[8:0]	rl_rg111_t ;
reg	rl_rg111_t_c1 ;
reg	rl_rg111_t_c2 ;
reg	[8:0]	rl_rg112_t ;
reg	rl_rg112_t_c1 ;
reg	rl_rg112_t_c2 ;
reg	[8:0]	rl_rg113_t ;
reg	rl_rg113_t_c1 ;
reg	rl_rg113_t_c2 ;
reg	[8:0]	rl_rg114_t ;
reg	rl_rg114_t_c1 ;
reg	rl_rg114_t_c2 ;
reg	[8:0]	rl_rg115_t ;
reg	rl_rg115_t_c1 ;
reg	rl_rg115_t_c2 ;
reg	[8:0]	rl_rg116_t ;
reg	rl_rg116_t_c1 ;
reg	rl_rg116_t_c2 ;
reg	[8:0]	rl_rg117_t ;
reg	rl_rg117_t_c1 ;
reg	rl_rg117_t_c2 ;
reg	[8:0]	rl_rg118_t ;
reg	rl_rg118_t_c1 ;
reg	rl_rg118_t_c2 ;
reg	[8:0]	rl_rg119_t ;
reg	rl_rg119_t_c1 ;
reg	rl_rg119_t_c2 ;
reg	[8:0]	rl_rg120_t ;
reg	rl_rg120_t_c1 ;
reg	rl_rg120_t_c2 ;
reg	[8:0]	rl_rg121_t ;
reg	rl_rg121_t_c1 ;
reg	rl_rg121_t_c2 ;
reg	[8:0]	rl_rg122_t ;
reg	rl_rg122_t_c1 ;
reg	rl_rg122_t_c2 ;
reg	[8:0]	rl_rg123_t ;
reg	rl_rg123_t_c1 ;
reg	rl_rg123_t_c2 ;
reg	[8:0]	rl_rg124_t ;
reg	rl_rg124_t_c1 ;
reg	rl_rg124_t_c2 ;
reg	[8:0]	rl_rg125_t ;
reg	rl_rg125_t_c1 ;
reg	rl_rg125_t_c2 ;
reg	[8:0]	rl_rg126_t ;
reg	rl_rg126_t_c1 ;
reg	rl_rg126_t_c2 ;
reg	[8:0]	rl_rg127_t ;
reg	rl_rg127_t_c1 ;
reg	rl_rg127_t_c2 ;
reg	M_01_t1 ;
reg	JF_08 ;
reg	CT_20 ;
reg	[8:0]	quantized_block_wd01 ;	// line#=../rle.cpp:22
reg	[3:0]	RG_y_02_t ;
reg	RG_y_02_t_c1 ;
reg	RG_y_02_t_c2 ;
reg	[3:0]	RG_j_x_02_t ;
reg	RG_j_x_02_t_c1 ;
reg	RG_j_x_02_t_c2 ;
reg	[31:0]	RG_i_06_t ;
reg	RG_i_06_t_c1 ;
reg	RG_i_06_t_c2 ;
reg	[7:0]	RG_len_05_t ;
reg	RG_len_05_t_c1 ;
reg	[2:0]	TR_02 ;
reg	[31:0]	RG_i_t ;
reg	RG_i_t_c1 ;
reg	RG_i_t_c2 ;
reg	[31:0]	RG_j_k_t ;
reg	RG_j_k_t_c1 ;
reg	RG_j_k_t_c2 ;
reg	RG_j_k_t_c3 ;
reg	[5:0]	RG_k_t ;
reg	FF_d_05_t ;
reg	FF_d_05_t_c1 ;
reg	FF_d_05_t_c2 ;
reg	RG_15_02_t ;
reg	[6:0]	RG_k_05_t ;
reg	FL01_01_streg_t ;
reg	FL01_01_streg_t_c1 ;
reg	FL01_01_streg_t_c2 ;
reg	FL01_02_streg_t ;
reg	FL01_02_streg_t_c1 ;
reg	FL01_02_streg_t_c2 ;
reg	flag_r1_t ;
reg	flag_r1_t_c1 ;
reg	flag_r2_t ;
reg	flag_r2_t_c1 ;
reg	flag_r3_t ;
reg	flag_r3_t_c1 ;
reg	[1:0]	FL02_01_streg_t ;
reg	FL02_01_streg_t_c1 ;
reg	FL02_01_streg_t_c2 ;
reg	[1:0]	FL02_02_streg_t ;
reg	FL02_02_streg_t_c1 ;
reg	FL02_02_streg_t_c2 ;
reg	[1:0]	FL02_02_streg_t1 ;
reg	FL02_02_streg_t1_c1 ;
reg	FL02_02_streg_t1_c2 ;
reg	FL02_02_streg_t1_c3 ;
reg	FL02_03_streg_t ;
reg	FL02_03_streg_t_c1 ;
reg	FL02_03_streg_t_c2 ;
reg	FL02_04_streg_t ;
reg	FL02_04_streg_t_c1 ;
reg	FL02_04_streg_t_c2 ;
reg	FL02_05_streg_t ;
reg	FL02_05_streg_t_c1 ;
reg	FL02_05_streg_t_c2 ;
reg	FL02_06_streg_t ;
reg	FL02_06_streg_t_c1 ;
reg	FL02_06_streg_t_c2 ;
reg	valid_r_t ;
reg	[2:0]	sub8u1i2 ;
reg	sub8u1i2_c1 ;
reg	[3:0]	incr4s1i1 ;
reg	[5:0]	zz_RA1 ;
reg	[5:0]	zz_WA2 ;
reg	[6:0]	rl_ad00 ;	// line#=../rle.cpp:23
reg	rl_ad00_c1 ;
reg	[8:0]	rl_wd01 ;	// line#=../rle.cpp:23
reg	[8:0]	rl_wd02 ;	// line#=../rle.cpp:23

jpeg_incr8u_6 INST_incr8u_6_1 ( .i1(incr8u_61i1) ,.o1(incr8u_61ot) );	// line#=../rle.cpp:111
jpeg_incr8u_7 INST_incr8u_7_1 ( .i1(incr8u_71i1) ,.o1(incr8u_71ot) );	// line#=../rle.cpp:142
jpeg_decr32s INST_decr32s_1 ( .i1(decr32s1i1) ,.o1(decr32s1ot) );	// line#=../rle.cpp:124,155
jpeg_decr32s INST_decr32s_2 ( .i1(decr32s2i1) ,.o1(decr32s2ot) );	// line#=../rle.cpp:130,161
jpeg_decr8u_7 INST_decr8u_7_1 ( .i1(decr8u_71i1) ,.o1(decr8u_71ot) );	// line#=../rle.cpp:77,78
jpeg_incr32s INST_incr32s_1 ( .i1(incr32s1i1) ,.o1(incr32s1ot) );	// line#=../rle.cpp:64,114,125,145,156
jpeg_incr32s INST_incr32s_2 ( .i1(incr32s2i1) ,.o1(incr32s2ot) );	// line#=../rle.cpp:61,62,63,119,129,150
									// ,160
jpeg_incr32s INST_incr32s_3 ( .i1(incr32s3i1) ,.o1(incr32s3ot) );	// line#=../rle.cpp:74
jpeg_incr8u INST_incr8u_1 ( .i1(incr8u1i1) ,.o1(incr8u1ot) );	// line#=../rle.cpp:68,73,79,80
jpeg_incr8u INST_incr8u_2 ( .i1(incr8u2i1) ,.o1(incr8u2ot) );	// line#=../rle.cpp:69,74
jpeg_incr4s INST_incr4s_1 ( .i1(incr4s1i1) ,.o1(incr4s1ot) );	// line#=../rle.cpp:34,44
jpeg_incr3u INST_incr3u_1 ( .i1(incr3u1i1) ,.o1(incr3u1ot) );	// line#=../rle.cpp:42
jpeg_lop8u_1 INST_lop8u_1_1 ( .i1(lop8u_11i1) ,.i2(lop8u_11i2) ,.o1(lop8u_11ot) );	// line#=../rle.cpp:109,110
assign	lop8u_11ot_port = lop8u_11ot ;
jpeg_sub12s_9 INST_sub12s_9_1 ( .i1(sub12s_91i1) ,.i2(sub12s_91i2) ,.o1(sub12s_91ot) );	// line#=../rle.cpp:52
jpeg_sub8u INST_sub8u_1 ( .i1(sub8u1i1) ,.i2(sub8u1i2) ,.o1(sub8u1ot) );	// line#=../rle.cpp:77,78,83,84,86
jpeg_add3u INST_add3u_1 ( .i1(add3u1i1) ,.i2(add3u1i2) ,.o1(add3u1ot) );	// line#=../rle.cpp:45
always @ ( U_103 or U_129 )
	FA02_02_gnt = ( { 1{ ~U_129 } } & U_103 )
		 ;
always @ ( U_108 or U_136 )
	FA02_03_gnt = ( { 1{ ~U_136 } } & U_108 )
		 ;
jpeg_MEMB9W64 zz ( .RA1(zz_RA1) ,.RD1(zz_RD1) ,.RCLK1(clk) ,.WA2(zz_WA2) ,.WD2(quantized_block_rd00) ,
	.WE2(zz_WE2) ,.WCLK2(clk) );	// line#=../rle.h:65
assign	jpeg_out_a00 = jpeg_out_a00_r ;	// line#=../rle.h:60
assign	jpeg_out_a01 = jpeg_out_a01_r ;	// line#=../rle.h:60
assign	jpeg_out_a02 = jpeg_out_a02_r ;	// line#=../rle.h:60
assign	jpeg_out_a03 = jpeg_out_a03_r ;	// line#=../rle.h:60
assign	jpeg_out_a04 = jpeg_out_a04_r ;	// line#=../rle.h:60
assign	jpeg_out_a05 = jpeg_out_a05_r ;	// line#=../rle.h:60
assign	jpeg_out_a06 = jpeg_out_a06_r ;	// line#=../rle.h:60
assign	jpeg_out_a07 = jpeg_out_a07_r ;	// line#=../rle.h:60
assign	jpeg_out_a08 = jpeg_out_a08_r ;	// line#=../rle.h:60
assign	jpeg_out_a09 = jpeg_out_a09_r ;	// line#=../rle.h:60
assign	jpeg_out_a10 = jpeg_out_a10_r ;	// line#=../rle.h:60
assign	jpeg_out_a11 = jpeg_out_a11_r ;	// line#=../rle.h:60
assign	jpeg_out_a12 = jpeg_out_a12_r ;	// line#=../rle.h:60
assign	jpeg_out_a13 = jpeg_out_a13_r ;	// line#=../rle.h:60
assign	jpeg_out_a14 = jpeg_out_a14_r ;	// line#=../rle.h:60
assign	jpeg_out_a15 = jpeg_out_a15_r ;	// line#=../rle.h:60
assign	jpeg_out_a16 = jpeg_out_a16_r ;	// line#=../rle.h:60
assign	jpeg_out_a17 = jpeg_out_a17_r ;	// line#=../rle.h:60
assign	jpeg_out_a18 = jpeg_out_a18_r ;	// line#=../rle.h:60
assign	jpeg_out_a19 = jpeg_out_a19_r ;	// line#=../rle.h:60
assign	jpeg_out_a20 = jpeg_out_a20_r ;	// line#=../rle.h:60
assign	jpeg_out_a21 = jpeg_out_a21_r ;	// line#=../rle.h:60
assign	jpeg_out_a22 = jpeg_out_a22_r ;	// line#=../rle.h:60
assign	jpeg_out_a23 = jpeg_out_a23_r ;	// line#=../rle.h:60
assign	jpeg_out_a24 = jpeg_out_a24_r ;	// line#=../rle.h:60
assign	jpeg_out_a25 = jpeg_out_a25_r ;	// line#=../rle.h:60
assign	jpeg_out_a26 = jpeg_out_a26_r ;	// line#=../rle.h:60
assign	jpeg_out_a27 = jpeg_out_a27_r ;	// line#=../rle.h:60
assign	jpeg_out_a28 = jpeg_out_a28_r ;	// line#=../rle.h:60
assign	jpeg_out_a29 = jpeg_out_a29_r ;	// line#=../rle.h:60
assign	jpeg_out_a30 = jpeg_out_a30_r ;	// line#=../rle.h:60
assign	jpeg_out_a31 = jpeg_out_a31_r ;	// line#=../rle.h:60
assign	jpeg_out_a32 = jpeg_out_a32_r ;	// line#=../rle.h:60
assign	jpeg_out_a33 = jpeg_out_a33_r ;	// line#=../rle.h:60
assign	jpeg_out_a34 = jpeg_out_a34_r ;	// line#=../rle.h:60
assign	jpeg_out_a35 = jpeg_out_a35_r ;	// line#=../rle.h:60
assign	jpeg_out_a36 = jpeg_out_a36_r ;	// line#=../rle.h:60
assign	jpeg_out_a37 = jpeg_out_a37_r ;	// line#=../rle.h:60
assign	jpeg_out_a38 = jpeg_out_a38_r ;	// line#=../rle.h:60
assign	jpeg_out_a39 = jpeg_out_a39_r ;	// line#=../rle.h:60
assign	jpeg_out_a40 = jpeg_out_a40_r ;	// line#=../rle.h:60
assign	jpeg_out_a41 = jpeg_out_a41_r ;	// line#=../rle.h:60
assign	jpeg_out_a42 = jpeg_out_a42_r ;	// line#=../rle.h:60
assign	jpeg_out_a43 = jpeg_out_a43_r ;	// line#=../rle.h:60
assign	jpeg_out_a44 = jpeg_out_a44_r ;	// line#=../rle.h:60
assign	jpeg_out_a45 = jpeg_out_a45_r ;	// line#=../rle.h:60
assign	jpeg_out_a46 = jpeg_out_a46_r ;	// line#=../rle.h:60
assign	jpeg_out_a47 = jpeg_out_a47_r ;	// line#=../rle.h:60
assign	jpeg_out_a48 = jpeg_out_a48_r ;	// line#=../rle.h:60
assign	jpeg_out_a49 = jpeg_out_a49_r ;	// line#=../rle.h:60
assign	jpeg_out_a50 = jpeg_out_a50_r ;	// line#=../rle.h:60
assign	jpeg_out_a51 = jpeg_out_a51_r ;	// line#=../rle.h:60
assign	jpeg_out_a52 = jpeg_out_a52_r ;	// line#=../rle.h:60
assign	jpeg_out_a53 = jpeg_out_a53_r ;	// line#=../rle.h:60
assign	jpeg_out_a54 = jpeg_out_a54_r ;	// line#=../rle.h:60
assign	jpeg_out_a55 = jpeg_out_a55_r ;	// line#=../rle.h:60
assign	jpeg_out_a56 = jpeg_out_a56_r ;	// line#=../rle.h:60
assign	jpeg_out_a57 = jpeg_out_a57_r ;	// line#=../rle.h:60
assign	jpeg_out_a58 = jpeg_out_a58_r ;	// line#=../rle.h:60
assign	jpeg_out_a59 = jpeg_out_a59_r ;	// line#=../rle.h:60
assign	jpeg_out_a60 = jpeg_out_a60_r ;	// line#=../rle.h:60
assign	jpeg_out_a61 = jpeg_out_a61_r ;	// line#=../rle.h:60
assign	jpeg_out_a62 = jpeg_out_a62_r ;	// line#=../rle.h:60
assign	jpeg_out_a63 = jpeg_out_a63_r ;	// line#=../rle.h:60
assign	jpeg_out_a64 = jpeg_out_a64_r ;	// line#=../rle.h:60
assign	jpeg_out_a65 = jpeg_out_a65_r ;	// line#=../rle.h:60
assign	jpeg_out_a66 = jpeg_out_a66_r ;	// line#=../rle.h:60
assign	jpeg_out_a67 = jpeg_out_a67_r ;	// line#=../rle.h:60
assign	jpeg_out_a68 = jpeg_out_a68_r ;	// line#=../rle.h:60
assign	jpeg_out_a69 = jpeg_out_a69_r ;	// line#=../rle.h:60
assign	jpeg_out_a70 = jpeg_out_a70_r ;	// line#=../rle.h:60
assign	jpeg_out_a71 = jpeg_out_a71_r ;	// line#=../rle.h:60
assign	jpeg_out_a72 = jpeg_out_a72_r ;	// line#=../rle.h:60
assign	jpeg_out_a73 = jpeg_out_a73_r ;	// line#=../rle.h:60
assign	jpeg_out_a74 = jpeg_out_a74_r ;	// line#=../rle.h:60
assign	jpeg_out_a75 = jpeg_out_a75_r ;	// line#=../rle.h:60
assign	jpeg_out_a76 = jpeg_out_a76_r ;	// line#=../rle.h:60
assign	jpeg_out_a77 = jpeg_out_a77_r ;	// line#=../rle.h:60
assign	jpeg_out_a78 = jpeg_out_a78_r ;	// line#=../rle.h:60
assign	jpeg_out_a79 = jpeg_out_a79_r ;	// line#=../rle.h:60
assign	jpeg_out_a80 = jpeg_out_a80_r ;	// line#=../rle.h:60
assign	jpeg_out_a81 = jpeg_out_a81_r ;	// line#=../rle.h:60
assign	jpeg_out_a82 = jpeg_out_a82_r ;	// line#=../rle.h:60
assign	jpeg_out_a83 = jpeg_out_a83_r ;	// line#=../rle.h:60
assign	jpeg_out_a84 = jpeg_out_a84_r ;	// line#=../rle.h:60
assign	jpeg_out_a85 = jpeg_out_a85_r ;	// line#=../rle.h:60
assign	jpeg_out_a86 = jpeg_out_a86_r ;	// line#=../rle.h:60
assign	jpeg_out_a87 = jpeg_out_a87_r ;	// line#=../rle.h:60
assign	jpeg_out_a88 = jpeg_out_a88_r ;	// line#=../rle.h:60
assign	jpeg_out_a89 = jpeg_out_a89_r ;	// line#=../rle.h:60
assign	jpeg_out_a90 = jpeg_out_a90_r ;	// line#=../rle.h:60
assign	jpeg_out_a91 = jpeg_out_a91_r ;	// line#=../rle.h:60
assign	jpeg_out_a92 = jpeg_out_a92_r ;	// line#=../rle.h:60
assign	jpeg_out_a93 = jpeg_out_a93_r ;	// line#=../rle.h:60
assign	jpeg_out_a94 = jpeg_out_a94_r ;	// line#=../rle.h:60
assign	jpeg_out_a95 = jpeg_out_a95_r ;	// line#=../rle.h:60
assign	jpeg_out_a96 = jpeg_out_a96_r ;	// line#=../rle.h:60
assign	jpeg_out_a97 = jpeg_out_a97_r ;	// line#=../rle.h:60
assign	jpeg_out_a98 = jpeg_out_a98_r ;	// line#=../rle.h:60
assign	jpeg_out_a99 = jpeg_out_a99_r ;	// line#=../rle.h:60
assign	jpeg_out_a100 = jpeg_out_a100_r ;	// line#=../rle.h:60
assign	jpeg_out_a101 = jpeg_out_a101_r ;	// line#=../rle.h:60
assign	jpeg_out_a102 = jpeg_out_a102_r ;	// line#=../rle.h:60
assign	jpeg_out_a103 = jpeg_out_a103_r ;	// line#=../rle.h:60
assign	jpeg_out_a104 = jpeg_out_a104_r ;	// line#=../rle.h:60
assign	jpeg_out_a105 = jpeg_out_a105_r ;	// line#=../rle.h:60
assign	jpeg_out_a106 = jpeg_out_a106_r ;	// line#=../rle.h:60
assign	jpeg_out_a107 = jpeg_out_a107_r ;	// line#=../rle.h:60
assign	jpeg_out_a108 = jpeg_out_a108_r ;	// line#=../rle.h:60
assign	jpeg_out_a109 = jpeg_out_a109_r ;	// line#=../rle.h:60
assign	jpeg_out_a110 = jpeg_out_a110_r ;	// line#=../rle.h:60
assign	jpeg_out_a111 = jpeg_out_a111_r ;	// line#=../rle.h:60
assign	jpeg_out_a112 = jpeg_out_a112_r ;	// line#=../rle.h:60
assign	jpeg_out_a113 = jpeg_out_a113_r ;	// line#=../rle.h:60
assign	jpeg_out_a114 = jpeg_out_a114_r ;	// line#=../rle.h:60
assign	jpeg_out_a115 = jpeg_out_a115_r ;	// line#=../rle.h:60
assign	jpeg_out_a116 = jpeg_out_a116_r ;	// line#=../rle.h:60
assign	jpeg_out_a117 = jpeg_out_a117_r ;	// line#=../rle.h:60
assign	jpeg_out_a118 = jpeg_out_a118_r ;	// line#=../rle.h:60
assign	jpeg_out_a119 = jpeg_out_a119_r ;	// line#=../rle.h:60
assign	jpeg_out_a120 = jpeg_out_a120_r ;	// line#=../rle.h:60
assign	jpeg_out_a121 = jpeg_out_a121_r ;	// line#=../rle.h:60
assign	jpeg_out_a122 = jpeg_out_a122_r ;	// line#=../rle.h:60
assign	jpeg_out_a123 = jpeg_out_a123_r ;	// line#=../rle.h:60
assign	jpeg_out_a124 = jpeg_out_a124_r ;	// line#=../rle.h:60
assign	jpeg_out_a125 = jpeg_out_a125_r ;	// line#=../rle.h:60
assign	jpeg_out_a126 = jpeg_out_a126_r ;	// line#=../rle.h:60
assign	jpeg_out_a127 = jpeg_out_a127_r ;	// line#=../rle.h:60
assign	jpeg_len_out = jpeg_len_out_r ;	// line#=../rle.h:61
assign	valid = valid_r ;	// line#=../rle.h:62
jpeg_decoder_6to64 INST_decoder_6to64_1 ( .DECODER_in(quantized_block_ad01) ,.DECODER_out(quantized_block_d01) );	// line#=../rle.cpp:22
always @ ( quantized_block_rg63 or quantized_block_rg62 or quantized_block_rg61 or 
	quantized_block_rg60 or quantized_block_rg59 or quantized_block_rg58 or 
	quantized_block_rg57 or quantized_block_rg56 or quantized_block_rg55 or 
	quantized_block_rg54 or quantized_block_rg53 or quantized_block_rg52 or 
	quantized_block_rg51 or quantized_block_rg50 or quantized_block_rg49 or 
	quantized_block_rg48 or quantized_block_rg47 or quantized_block_rg46 or 
	quantized_block_rg45 or quantized_block_rg44 or quantized_block_rg43 or 
	quantized_block_rg42 or quantized_block_rg41 or quantized_block_rg40 or 
	quantized_block_rg39 or quantized_block_rg38 or quantized_block_rg37 or 
	quantized_block_rg36 or quantized_block_rg35 or quantized_block_rg34 or 
	quantized_block_rg33 or quantized_block_rg32 or quantized_block_rg31 or 
	quantized_block_rg30 or quantized_block_rg29 or quantized_block_rg28 or 
	quantized_block_rg27 or quantized_block_rg26 or quantized_block_rg25 or 
	quantized_block_rg24 or quantized_block_rg23 or quantized_block_rg22 or 
	quantized_block_rg21 or quantized_block_rg20 or quantized_block_rg19 or 
	quantized_block_rg18 or quantized_block_rg17 or quantized_block_rg16 or 
	quantized_block_rg15 or quantized_block_rg14 or quantized_block_rg13 or 
	quantized_block_rg12 or quantized_block_rg11 or quantized_block_rg10 or 
	quantized_block_rg09 or quantized_block_rg08 or quantized_block_rg07 or 
	quantized_block_rg06 or quantized_block_rg05 or quantized_block_rg04 or 
	quantized_block_rg03 or quantized_block_rg02 or quantized_block_rg01 or 
	quantized_block_rg00 or RG_j_k or RG_i )	// line#=../rle.cpp:22,111,142
	case ( { RG_i [2:0] , RG_j_k [2:0] } )
	6'h00 :
		quantized_block_rd00 = quantized_block_rg00 ;
	6'h01 :
		quantized_block_rd00 = quantized_block_rg01 ;
	6'h02 :
		quantized_block_rd00 = quantized_block_rg02 ;
	6'h03 :
		quantized_block_rd00 = quantized_block_rg03 ;
	6'h04 :
		quantized_block_rd00 = quantized_block_rg04 ;
	6'h05 :
		quantized_block_rd00 = quantized_block_rg05 ;
	6'h06 :
		quantized_block_rd00 = quantized_block_rg06 ;
	6'h07 :
		quantized_block_rd00 = quantized_block_rg07 ;
	6'h08 :
		quantized_block_rd00 = quantized_block_rg08 ;
	6'h09 :
		quantized_block_rd00 = quantized_block_rg09 ;
	6'h0a :
		quantized_block_rd00 = quantized_block_rg10 ;
	6'h0b :
		quantized_block_rd00 = quantized_block_rg11 ;
	6'h0c :
		quantized_block_rd00 = quantized_block_rg12 ;
	6'h0d :
		quantized_block_rd00 = quantized_block_rg13 ;
	6'h0e :
		quantized_block_rd00 = quantized_block_rg14 ;
	6'h0f :
		quantized_block_rd00 = quantized_block_rg15 ;
	6'h10 :
		quantized_block_rd00 = quantized_block_rg16 ;
	6'h11 :
		quantized_block_rd00 = quantized_block_rg17 ;
	6'h12 :
		quantized_block_rd00 = quantized_block_rg18 ;
	6'h13 :
		quantized_block_rd00 = quantized_block_rg19 ;
	6'h14 :
		quantized_block_rd00 = quantized_block_rg20 ;
	6'h15 :
		quantized_block_rd00 = quantized_block_rg21 ;
	6'h16 :
		quantized_block_rd00 = quantized_block_rg22 ;
	6'h17 :
		quantized_block_rd00 = quantized_block_rg23 ;
	6'h18 :
		quantized_block_rd00 = quantized_block_rg24 ;
	6'h19 :
		quantized_block_rd00 = quantized_block_rg25 ;
	6'h1a :
		quantized_block_rd00 = quantized_block_rg26 ;
	6'h1b :
		quantized_block_rd00 = quantized_block_rg27 ;
	6'h1c :
		quantized_block_rd00 = quantized_block_rg28 ;
	6'h1d :
		quantized_block_rd00 = quantized_block_rg29 ;
	6'h1e :
		quantized_block_rd00 = quantized_block_rg30 ;
	6'h1f :
		quantized_block_rd00 = quantized_block_rg31 ;
	6'h20 :
		quantized_block_rd00 = quantized_block_rg32 ;
	6'h21 :
		quantized_block_rd00 = quantized_block_rg33 ;
	6'h22 :
		quantized_block_rd00 = quantized_block_rg34 ;
	6'h23 :
		quantized_block_rd00 = quantized_block_rg35 ;
	6'h24 :
		quantized_block_rd00 = quantized_block_rg36 ;
	6'h25 :
		quantized_block_rd00 = quantized_block_rg37 ;
	6'h26 :
		quantized_block_rd00 = quantized_block_rg38 ;
	6'h27 :
		quantized_block_rd00 = quantized_block_rg39 ;
	6'h28 :
		quantized_block_rd00 = quantized_block_rg40 ;
	6'h29 :
		quantized_block_rd00 = quantized_block_rg41 ;
	6'h2a :
		quantized_block_rd00 = quantized_block_rg42 ;
	6'h2b :
		quantized_block_rd00 = quantized_block_rg43 ;
	6'h2c :
		quantized_block_rd00 = quantized_block_rg44 ;
	6'h2d :
		quantized_block_rd00 = quantized_block_rg45 ;
	6'h2e :
		quantized_block_rd00 = quantized_block_rg46 ;
	6'h2f :
		quantized_block_rd00 = quantized_block_rg47 ;
	6'h30 :
		quantized_block_rd00 = quantized_block_rg48 ;
	6'h31 :
		quantized_block_rd00 = quantized_block_rg49 ;
	6'h32 :
		quantized_block_rd00 = quantized_block_rg50 ;
	6'h33 :
		quantized_block_rd00 = quantized_block_rg51 ;
	6'h34 :
		quantized_block_rd00 = quantized_block_rg52 ;
	6'h35 :
		quantized_block_rd00 = quantized_block_rg53 ;
	6'h36 :
		quantized_block_rd00 = quantized_block_rg54 ;
	6'h37 :
		quantized_block_rd00 = quantized_block_rg55 ;
	6'h38 :
		quantized_block_rd00 = quantized_block_rg56 ;
	6'h39 :
		quantized_block_rd00 = quantized_block_rg57 ;
	6'h3a :
		quantized_block_rd00 = quantized_block_rg58 ;
	6'h3b :
		quantized_block_rd00 = quantized_block_rg59 ;
	6'h3c :
		quantized_block_rd00 = quantized_block_rg60 ;
	6'h3d :
		quantized_block_rd00 = quantized_block_rg61 ;
	6'h3e :
		quantized_block_rd00 = quantized_block_rg62 ;
	6'h3f :
		quantized_block_rd00 = quantized_block_rg63 ;
	default :
		quantized_block_rd00 = 9'hx ;
	endcase
assign	quantized_block_rg00_en = ( U_10 & quantized_block_d01 [63] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg00 <= 9'h000 ;
	else if ( quantized_block_rg00_en )
		quantized_block_rg00 <= quantized_block_wd01 ;
assign	quantized_block_rg01_en = ( U_10 & quantized_block_d01 [62] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg01 <= 9'h000 ;
	else if ( quantized_block_rg01_en )
		quantized_block_rg01 <= quantized_block_wd01 ;
assign	quantized_block_rg02_en = ( U_10 & quantized_block_d01 [61] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg02 <= 9'h000 ;
	else if ( quantized_block_rg02_en )
		quantized_block_rg02 <= quantized_block_wd01 ;
assign	quantized_block_rg03_en = ( U_10 & quantized_block_d01 [60] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg03 <= 9'h000 ;
	else if ( quantized_block_rg03_en )
		quantized_block_rg03 <= quantized_block_wd01 ;
assign	quantized_block_rg04_en = ( U_10 & quantized_block_d01 [59] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg04 <= 9'h000 ;
	else if ( quantized_block_rg04_en )
		quantized_block_rg04 <= quantized_block_wd01 ;
assign	quantized_block_rg05_en = ( U_10 & quantized_block_d01 [58] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg05 <= 9'h000 ;
	else if ( quantized_block_rg05_en )
		quantized_block_rg05 <= quantized_block_wd01 ;
assign	quantized_block_rg06_en = ( U_10 & quantized_block_d01 [57] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg06 <= 9'h000 ;
	else if ( quantized_block_rg06_en )
		quantized_block_rg06 <= quantized_block_wd01 ;
assign	quantized_block_rg07_en = ( U_10 & quantized_block_d01 [56] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg07 <= 9'h000 ;
	else if ( quantized_block_rg07_en )
		quantized_block_rg07 <= quantized_block_wd01 ;
assign	quantized_block_rg08_en = ( U_10 & quantized_block_d01 [55] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg08 <= 9'h000 ;
	else if ( quantized_block_rg08_en )
		quantized_block_rg08 <= quantized_block_wd01 ;
assign	quantized_block_rg09_en = ( U_10 & quantized_block_d01 [54] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg09 <= 9'h000 ;
	else if ( quantized_block_rg09_en )
		quantized_block_rg09 <= quantized_block_wd01 ;
assign	quantized_block_rg10_en = ( U_10 & quantized_block_d01 [53] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg10 <= 9'h000 ;
	else if ( quantized_block_rg10_en )
		quantized_block_rg10 <= quantized_block_wd01 ;
assign	quantized_block_rg11_en = ( U_10 & quantized_block_d01 [52] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg11 <= 9'h000 ;
	else if ( quantized_block_rg11_en )
		quantized_block_rg11 <= quantized_block_wd01 ;
assign	quantized_block_rg12_en = ( U_10 & quantized_block_d01 [51] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg12 <= 9'h000 ;
	else if ( quantized_block_rg12_en )
		quantized_block_rg12 <= quantized_block_wd01 ;
assign	quantized_block_rg13_en = ( U_10 & quantized_block_d01 [50] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg13 <= 9'h000 ;
	else if ( quantized_block_rg13_en )
		quantized_block_rg13 <= quantized_block_wd01 ;
assign	quantized_block_rg14_en = ( U_10 & quantized_block_d01 [49] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg14 <= 9'h000 ;
	else if ( quantized_block_rg14_en )
		quantized_block_rg14 <= quantized_block_wd01 ;
assign	quantized_block_rg15_en = ( U_10 & quantized_block_d01 [48] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg15 <= 9'h000 ;
	else if ( quantized_block_rg15_en )
		quantized_block_rg15 <= quantized_block_wd01 ;
assign	quantized_block_rg16_en = ( U_10 & quantized_block_d01 [47] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg16 <= 9'h000 ;
	else if ( quantized_block_rg16_en )
		quantized_block_rg16 <= quantized_block_wd01 ;
assign	quantized_block_rg17_en = ( U_10 & quantized_block_d01 [46] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg17 <= 9'h000 ;
	else if ( quantized_block_rg17_en )
		quantized_block_rg17 <= quantized_block_wd01 ;
assign	quantized_block_rg18_en = ( U_10 & quantized_block_d01 [45] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg18 <= 9'h000 ;
	else if ( quantized_block_rg18_en )
		quantized_block_rg18 <= quantized_block_wd01 ;
assign	quantized_block_rg19_en = ( U_10 & quantized_block_d01 [44] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg19 <= 9'h000 ;
	else if ( quantized_block_rg19_en )
		quantized_block_rg19 <= quantized_block_wd01 ;
assign	quantized_block_rg20_en = ( U_10 & quantized_block_d01 [43] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg20 <= 9'h000 ;
	else if ( quantized_block_rg20_en )
		quantized_block_rg20 <= quantized_block_wd01 ;
assign	quantized_block_rg21_en = ( U_10 & quantized_block_d01 [42] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg21 <= 9'h000 ;
	else if ( quantized_block_rg21_en )
		quantized_block_rg21 <= quantized_block_wd01 ;
assign	quantized_block_rg22_en = ( U_10 & quantized_block_d01 [41] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg22 <= 9'h000 ;
	else if ( quantized_block_rg22_en )
		quantized_block_rg22 <= quantized_block_wd01 ;
assign	quantized_block_rg23_en = ( U_10 & quantized_block_d01 [40] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg23 <= 9'h000 ;
	else if ( quantized_block_rg23_en )
		quantized_block_rg23 <= quantized_block_wd01 ;
assign	quantized_block_rg24_en = ( U_10 & quantized_block_d01 [39] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg24 <= 9'h000 ;
	else if ( quantized_block_rg24_en )
		quantized_block_rg24 <= quantized_block_wd01 ;
assign	quantized_block_rg25_en = ( U_10 & quantized_block_d01 [38] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg25 <= 9'h000 ;
	else if ( quantized_block_rg25_en )
		quantized_block_rg25 <= quantized_block_wd01 ;
assign	quantized_block_rg26_en = ( U_10 & quantized_block_d01 [37] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg26 <= 9'h000 ;
	else if ( quantized_block_rg26_en )
		quantized_block_rg26 <= quantized_block_wd01 ;
assign	quantized_block_rg27_en = ( U_10 & quantized_block_d01 [36] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg27 <= 9'h000 ;
	else if ( quantized_block_rg27_en )
		quantized_block_rg27 <= quantized_block_wd01 ;
assign	quantized_block_rg28_en = ( U_10 & quantized_block_d01 [35] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg28 <= 9'h000 ;
	else if ( quantized_block_rg28_en )
		quantized_block_rg28 <= quantized_block_wd01 ;
assign	quantized_block_rg29_en = ( U_10 & quantized_block_d01 [34] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg29 <= 9'h000 ;
	else if ( quantized_block_rg29_en )
		quantized_block_rg29 <= quantized_block_wd01 ;
assign	quantized_block_rg30_en = ( U_10 & quantized_block_d01 [33] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg30 <= 9'h000 ;
	else if ( quantized_block_rg30_en )
		quantized_block_rg30 <= quantized_block_wd01 ;
assign	quantized_block_rg31_en = ( U_10 & quantized_block_d01 [32] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg31 <= 9'h000 ;
	else if ( quantized_block_rg31_en )
		quantized_block_rg31 <= quantized_block_wd01 ;
assign	quantized_block_rg32_en = ( U_10 & quantized_block_d01 [31] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg32 <= 9'h000 ;
	else if ( quantized_block_rg32_en )
		quantized_block_rg32 <= quantized_block_wd01 ;
assign	quantized_block_rg33_en = ( U_10 & quantized_block_d01 [30] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg33 <= 9'h000 ;
	else if ( quantized_block_rg33_en )
		quantized_block_rg33 <= quantized_block_wd01 ;
assign	quantized_block_rg34_en = ( U_10 & quantized_block_d01 [29] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg34 <= 9'h000 ;
	else if ( quantized_block_rg34_en )
		quantized_block_rg34 <= quantized_block_wd01 ;
assign	quantized_block_rg35_en = ( U_10 & quantized_block_d01 [28] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg35 <= 9'h000 ;
	else if ( quantized_block_rg35_en )
		quantized_block_rg35 <= quantized_block_wd01 ;
assign	quantized_block_rg36_en = ( U_10 & quantized_block_d01 [27] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg36 <= 9'h000 ;
	else if ( quantized_block_rg36_en )
		quantized_block_rg36 <= quantized_block_wd01 ;
assign	quantized_block_rg37_en = ( U_10 & quantized_block_d01 [26] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg37 <= 9'h000 ;
	else if ( quantized_block_rg37_en )
		quantized_block_rg37 <= quantized_block_wd01 ;
assign	quantized_block_rg38_en = ( U_10 & quantized_block_d01 [25] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg38 <= 9'h000 ;
	else if ( quantized_block_rg38_en )
		quantized_block_rg38 <= quantized_block_wd01 ;
assign	quantized_block_rg39_en = ( U_10 & quantized_block_d01 [24] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg39 <= 9'h000 ;
	else if ( quantized_block_rg39_en )
		quantized_block_rg39 <= quantized_block_wd01 ;
assign	quantized_block_rg40_en = ( U_10 & quantized_block_d01 [23] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg40 <= 9'h000 ;
	else if ( quantized_block_rg40_en )
		quantized_block_rg40 <= quantized_block_wd01 ;
assign	quantized_block_rg41_en = ( U_10 & quantized_block_d01 [22] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg41 <= 9'h000 ;
	else if ( quantized_block_rg41_en )
		quantized_block_rg41 <= quantized_block_wd01 ;
assign	quantized_block_rg42_en = ( U_10 & quantized_block_d01 [21] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg42 <= 9'h000 ;
	else if ( quantized_block_rg42_en )
		quantized_block_rg42 <= quantized_block_wd01 ;
assign	quantized_block_rg43_en = ( U_10 & quantized_block_d01 [20] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg43 <= 9'h000 ;
	else if ( quantized_block_rg43_en )
		quantized_block_rg43 <= quantized_block_wd01 ;
assign	quantized_block_rg44_en = ( U_10 & quantized_block_d01 [19] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg44 <= 9'h000 ;
	else if ( quantized_block_rg44_en )
		quantized_block_rg44 <= quantized_block_wd01 ;
assign	quantized_block_rg45_en = ( U_10 & quantized_block_d01 [18] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg45 <= 9'h000 ;
	else if ( quantized_block_rg45_en )
		quantized_block_rg45 <= quantized_block_wd01 ;
assign	quantized_block_rg46_en = ( U_10 & quantized_block_d01 [17] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg46 <= 9'h000 ;
	else if ( quantized_block_rg46_en )
		quantized_block_rg46 <= quantized_block_wd01 ;
assign	quantized_block_rg47_en = ( U_10 & quantized_block_d01 [16] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg47 <= 9'h000 ;
	else if ( quantized_block_rg47_en )
		quantized_block_rg47 <= quantized_block_wd01 ;
assign	quantized_block_rg48_en = ( U_10 & quantized_block_d01 [15] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg48 <= 9'h000 ;
	else if ( quantized_block_rg48_en )
		quantized_block_rg48 <= quantized_block_wd01 ;
assign	quantized_block_rg49_en = ( U_10 & quantized_block_d01 [14] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg49 <= 9'h000 ;
	else if ( quantized_block_rg49_en )
		quantized_block_rg49 <= quantized_block_wd01 ;
assign	quantized_block_rg50_en = ( U_10 & quantized_block_d01 [13] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg50 <= 9'h000 ;
	else if ( quantized_block_rg50_en )
		quantized_block_rg50 <= quantized_block_wd01 ;
assign	quantized_block_rg51_en = ( U_10 & quantized_block_d01 [12] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg51 <= 9'h000 ;
	else if ( quantized_block_rg51_en )
		quantized_block_rg51 <= quantized_block_wd01 ;
assign	quantized_block_rg52_en = ( U_10 & quantized_block_d01 [11] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg52 <= 9'h000 ;
	else if ( quantized_block_rg52_en )
		quantized_block_rg52 <= quantized_block_wd01 ;
assign	quantized_block_rg53_en = ( U_10 & quantized_block_d01 [10] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg53 <= 9'h000 ;
	else if ( quantized_block_rg53_en )
		quantized_block_rg53 <= quantized_block_wd01 ;
assign	quantized_block_rg54_en = ( U_10 & quantized_block_d01 [9] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg54 <= 9'h000 ;
	else if ( quantized_block_rg54_en )
		quantized_block_rg54 <= quantized_block_wd01 ;
assign	quantized_block_rg55_en = ( U_10 & quantized_block_d01 [8] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg55 <= 9'h000 ;
	else if ( quantized_block_rg55_en )
		quantized_block_rg55 <= quantized_block_wd01 ;
assign	quantized_block_rg56_en = ( U_10 & quantized_block_d01 [7] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg56 <= 9'h000 ;
	else if ( quantized_block_rg56_en )
		quantized_block_rg56 <= quantized_block_wd01 ;
assign	quantized_block_rg57_en = ( U_10 & quantized_block_d01 [6] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg57 <= 9'h000 ;
	else if ( quantized_block_rg57_en )
		quantized_block_rg57 <= quantized_block_wd01 ;
assign	quantized_block_rg58_en = ( U_10 & quantized_block_d01 [5] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg58 <= 9'h000 ;
	else if ( quantized_block_rg58_en )
		quantized_block_rg58 <= quantized_block_wd01 ;
assign	quantized_block_rg59_en = ( U_10 & quantized_block_d01 [4] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg59 <= 9'h000 ;
	else if ( quantized_block_rg59_en )
		quantized_block_rg59 <= quantized_block_wd01 ;
assign	quantized_block_rg60_en = ( U_10 & quantized_block_d01 [3] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg60 <= 9'h000 ;
	else if ( quantized_block_rg60_en )
		quantized_block_rg60 <= quantized_block_wd01 ;
assign	quantized_block_rg61_en = ( U_10 & quantized_block_d01 [2] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg61 <= 9'h000 ;
	else if ( quantized_block_rg61_en )
		quantized_block_rg61 <= quantized_block_wd01 ;
assign	quantized_block_rg62_en = ( U_10 & quantized_block_d01 [1] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg62 <= 9'h000 ;
	else if ( quantized_block_rg62_en )
		quantized_block_rg62 <= quantized_block_wd01 ;
assign	quantized_block_rg63_en = ( U_10 & quantized_block_d01 [0] ) ;
always @ ( posedge clk )	// line#=../rle.cpp:22,45
	if ( !rst )
		quantized_block_rg63 <= 9'h000 ;
	else if ( quantized_block_rg63_en )
		quantized_block_rg63 <= quantized_block_wd01 ;
jpeg_decoder_7to128 INST_decoder_7to128_1 ( .DECODER_in(rl_ad01) ,.DECODER_out(rl_d01) );	// line#=../rle.cpp:23
jpeg_decoder_7to128 INST_decoder_7to128_2 ( .DECODER_in(rl_ad02) ,.DECODER_out(rl_d02) );	// line#=../rle.cpp:23
always @ ( rl_rg127 or rl_rg126 or rl_rg125 or rl_rg124 or rl_rg123 or rl_rg122 or 
	rl_rg121 or rl_rg120 or rl_rg119 or rl_rg118 or rl_rg117 or rl_rg116 or 
	rl_rg115 or rl_rg114 or rl_rg113 or rl_rg112 or rl_rg111 or rl_rg110 or 
	rl_rg109 or rl_rg108 or rl_rg107 or rl_rg106 or rl_rg105 or rl_rg104 or 
	rl_rg103 or rl_rg102 or rl_rg101 or rl_rg100 or rl_rg99 or rl_rg98 or rl_rg97 or 
	rl_rg96 or rl_rg95 or rl_rg94 or rl_rg93 or rl_rg92 or rl_rg91 or rl_rg90 or 
	rl_rg89 or rl_rg88 or rl_rg87 or rl_rg86 or rl_rg85 or rl_rg84 or rl_rg83 or 
	rl_rg82 or rl_rg81 or rl_rg80 or rl_rg79 or rl_rg78 or rl_rg77 or rl_rg76 or 
	rl_rg75 or rl_rg74 or rl_rg73 or rl_rg72 or rl_rg71 or rl_rg70 or rl_rg69 or 
	rl_rg68 or rl_rg67 or rl_rg66 or rl_rg65 or rl_rg64 or rl_rg63 or rl_rg62 or 
	rl_rg61 or rl_rg60 or rl_rg59 or rl_rg58 or rl_rg57 or rl_rg56 or rl_rg55 or 
	rl_rg54 or rl_rg53 or rl_rg52 or rl_rg51 or rl_rg50 or rl_rg49 or rl_rg48 or 
	rl_rg47 or rl_rg46 or rl_rg45 or rl_rg44 or rl_rg43 or rl_rg42 or rl_rg41 or 
	rl_rg40 or rl_rg39 or rl_rg38 or rl_rg37 or rl_rg36 or rl_rg35 or rl_rg34 or 
	rl_rg33 or rl_rg32 or rl_rg31 or rl_rg30 or rl_rg29 or rl_rg28 or rl_rg27 or 
	rl_rg26 or rl_rg25 or rl_rg24 or rl_rg23 or rl_rg22 or rl_rg21 or rl_rg20 or 
	rl_rg19 or rl_rg18 or rl_rg17 or rl_rg16 or rl_rg15 or rl_rg14 or rl_rg13 or 
	rl_rg12 or rl_rg11 or rl_rg10 or rl_rg09 or rl_rg08 or rl_rg07 or rl_rg06 or 
	rl_rg05 or rl_rg04 or rl_rg03 or rl_rg02 or rl_rg01 or rl_rg00 or rl_ad00 )	// line#=../rle.cpp:23
	case ( rl_ad00 )
	7'h00 :
		rl_rd00 = rl_rg00 ;
	7'h01 :
		rl_rd00 = rl_rg01 ;
	7'h02 :
		rl_rd00 = rl_rg02 ;
	7'h03 :
		rl_rd00 = rl_rg03 ;
	7'h04 :
		rl_rd00 = rl_rg04 ;
	7'h05 :
		rl_rd00 = rl_rg05 ;
	7'h06 :
		rl_rd00 = rl_rg06 ;
	7'h07 :
		rl_rd00 = rl_rg07 ;
	7'h08 :
		rl_rd00 = rl_rg08 ;
	7'h09 :
		rl_rd00 = rl_rg09 ;
	7'h0a :
		rl_rd00 = rl_rg10 ;
	7'h0b :
		rl_rd00 = rl_rg11 ;
	7'h0c :
		rl_rd00 = rl_rg12 ;
	7'h0d :
		rl_rd00 = rl_rg13 ;
	7'h0e :
		rl_rd00 = rl_rg14 ;
	7'h0f :
		rl_rd00 = rl_rg15 ;
	7'h10 :
		rl_rd00 = rl_rg16 ;
	7'h11 :
		rl_rd00 = rl_rg17 ;
	7'h12 :
		rl_rd00 = rl_rg18 ;
	7'h13 :
		rl_rd00 = rl_rg19 ;
	7'h14 :
		rl_rd00 = rl_rg20 ;
	7'h15 :
		rl_rd00 = rl_rg21 ;
	7'h16 :
		rl_rd00 = rl_rg22 ;
	7'h17 :
		rl_rd00 = rl_rg23 ;
	7'h18 :
		rl_rd00 = rl_rg24 ;
	7'h19 :
		rl_rd00 = rl_rg25 ;
	7'h1a :
		rl_rd00 = rl_rg26 ;
	7'h1b :
		rl_rd00 = rl_rg27 ;
	7'h1c :
		rl_rd00 = rl_rg28 ;
	7'h1d :
		rl_rd00 = rl_rg29 ;
	7'h1e :
		rl_rd00 = rl_rg30 ;
	7'h1f :
		rl_rd00 = rl_rg31 ;
	7'h20 :
		rl_rd00 = rl_rg32 ;
	7'h21 :
		rl_rd00 = rl_rg33 ;
	7'h22 :
		rl_rd00 = rl_rg34 ;
	7'h23 :
		rl_rd00 = rl_rg35 ;
	7'h24 :
		rl_rd00 = rl_rg36 ;
	7'h25 :
		rl_rd00 = rl_rg37 ;
	7'h26 :
		rl_rd00 = rl_rg38 ;
	7'h27 :
		rl_rd00 = rl_rg39 ;
	7'h28 :
		rl_rd00 = rl_rg40 ;
	7'h29 :
		rl_rd00 = rl_rg41 ;
	7'h2a :
		rl_rd00 = rl_rg42 ;
	7'h2b :
		rl_rd00 = rl_rg43 ;
	7'h2c :
		rl_rd00 = rl_rg44 ;
	7'h2d :
		rl_rd00 = rl_rg45 ;
	7'h2e :
		rl_rd00 = rl_rg46 ;
	7'h2f :
		rl_rd00 = rl_rg47 ;
	7'h30 :
		rl_rd00 = rl_rg48 ;
	7'h31 :
		rl_rd00 = rl_rg49 ;
	7'h32 :
		rl_rd00 = rl_rg50 ;
	7'h33 :
		rl_rd00 = rl_rg51 ;
	7'h34 :
		rl_rd00 = rl_rg52 ;
	7'h35 :
		rl_rd00 = rl_rg53 ;
	7'h36 :
		rl_rd00 = rl_rg54 ;
	7'h37 :
		rl_rd00 = rl_rg55 ;
	7'h38 :
		rl_rd00 = rl_rg56 ;
	7'h39 :
		rl_rd00 = rl_rg57 ;
	7'h3a :
		rl_rd00 = rl_rg58 ;
	7'h3b :
		rl_rd00 = rl_rg59 ;
	7'h3c :
		rl_rd00 = rl_rg60 ;
	7'h3d :
		rl_rd00 = rl_rg61 ;
	7'h3e :
		rl_rd00 = rl_rg62 ;
	7'h3f :
		rl_rd00 = rl_rg63 ;
	7'h40 :
		rl_rd00 = rl_rg64 ;
	7'h41 :
		rl_rd00 = rl_rg65 ;
	7'h42 :
		rl_rd00 = rl_rg66 ;
	7'h43 :
		rl_rd00 = rl_rg67 ;
	7'h44 :
		rl_rd00 = rl_rg68 ;
	7'h45 :
		rl_rd00 = rl_rg69 ;
	7'h46 :
		rl_rd00 = rl_rg70 ;
	7'h47 :
		rl_rd00 = rl_rg71 ;
	7'h48 :
		rl_rd00 = rl_rg72 ;
	7'h49 :
		rl_rd00 = rl_rg73 ;
	7'h4a :
		rl_rd00 = rl_rg74 ;
	7'h4b :
		rl_rd00 = rl_rg75 ;
	7'h4c :
		rl_rd00 = rl_rg76 ;
	7'h4d :
		rl_rd00 = rl_rg77 ;
	7'h4e :
		rl_rd00 = rl_rg78 ;
	7'h4f :
		rl_rd00 = rl_rg79 ;
	7'h50 :
		rl_rd00 = rl_rg80 ;
	7'h51 :
		rl_rd00 = rl_rg81 ;
	7'h52 :
		rl_rd00 = rl_rg82 ;
	7'h53 :
		rl_rd00 = rl_rg83 ;
	7'h54 :
		rl_rd00 = rl_rg84 ;
	7'h55 :
		rl_rd00 = rl_rg85 ;
	7'h56 :
		rl_rd00 = rl_rg86 ;
	7'h57 :
		rl_rd00 = rl_rg87 ;
	7'h58 :
		rl_rd00 = rl_rg88 ;
	7'h59 :
		rl_rd00 = rl_rg89 ;
	7'h5a :
		rl_rd00 = rl_rg90 ;
	7'h5b :
		rl_rd00 = rl_rg91 ;
	7'h5c :
		rl_rd00 = rl_rg92 ;
	7'h5d :
		rl_rd00 = rl_rg93 ;
	7'h5e :
		rl_rd00 = rl_rg94 ;
	7'h5f :
		rl_rd00 = rl_rg95 ;
	7'h60 :
		rl_rd00 = rl_rg96 ;
	7'h61 :
		rl_rd00 = rl_rg97 ;
	7'h62 :
		rl_rd00 = rl_rg98 ;
	7'h63 :
		rl_rd00 = rl_rg99 ;
	7'h64 :
		rl_rd00 = rl_rg100 ;
	7'h65 :
		rl_rd00 = rl_rg101 ;
	7'h66 :
		rl_rd00 = rl_rg102 ;
	7'h67 :
		rl_rd00 = rl_rg103 ;
	7'h68 :
		rl_rd00 = rl_rg104 ;
	7'h69 :
		rl_rd00 = rl_rg105 ;
	7'h6a :
		rl_rd00 = rl_rg106 ;
	7'h6b :
		rl_rd00 = rl_rg107 ;
	7'h6c :
		rl_rd00 = rl_rg108 ;
	7'h6d :
		rl_rd00 = rl_rg109 ;
	7'h6e :
		rl_rd00 = rl_rg110 ;
	7'h6f :
		rl_rd00 = rl_rg111 ;
	7'h70 :
		rl_rd00 = rl_rg112 ;
	7'h71 :
		rl_rd00 = rl_rg113 ;
	7'h72 :
		rl_rd00 = rl_rg114 ;
	7'h73 :
		rl_rd00 = rl_rg115 ;
	7'h74 :
		rl_rd00 = rl_rg116 ;
	7'h75 :
		rl_rd00 = rl_rg117 ;
	7'h76 :
		rl_rd00 = rl_rg118 ;
	7'h77 :
		rl_rd00 = rl_rg119 ;
	7'h78 :
		rl_rd00 = rl_rg120 ;
	7'h79 :
		rl_rd00 = rl_rg121 ;
	7'h7a :
		rl_rd00 = rl_rg122 ;
	7'h7b :
		rl_rd00 = rl_rg123 ;
	7'h7c :
		rl_rd00 = rl_rg124 ;
	7'h7d :
		rl_rd00 = rl_rg125 ;
	7'h7e :
		rl_rd00 = rl_rg126 ;
	7'h7f :
		rl_rd00 = rl_rg127 ;
	default :
		rl_rd00 = 9'hx ;
	endcase
assign	M_01 = ~( ( rl_we01 & rl_d01 [127] ) | ( rl_we02 & rl_d02 [127] ) ) ;
always @ ( sub12s_91ot or M_01 or ST1_07d or rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or 
	rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg00_t_c1 = ( rl_we01 & rl_d01 [127] ) ;
	rl_rg00_t_c2 = ( rl_we02 & rl_d02 [127] ) ;
	rl_rg00_t_c3 = ( ST1_07d & M_01 ) ;	// line#=../rle.cpp:52
	rl_rg00_t = ( ( { 9{ rl_rg00_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg00_t_c2 } } & rl_wd02 )
		| ( { 9{ rl_rg00_t_c3 } } & sub12s_91ot )	// line#=../rle.cpp:52
		) ;
	end
assign	rl_rg00_en = ( rl_rg00_t_c1 | rl_rg00_t_c2 | rl_rg00_t_c3 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg00 <= 9'h000 ;
	else if ( rl_rg00_en )
		rl_rg00 <= rl_rg00_t ;	// line#=../rle.cpp:23,52
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg01_t_c1 = ( rl_we01 & rl_d01 [126] ) ;
	rl_rg01_t_c2 = ( rl_we02 & rl_d02 [126] ) ;
	rl_rg01_t = ( ( { 9{ rl_rg01_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg01_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg01_en = ( rl_rg01_t_c1 | rl_rg01_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg01 <= 9'h000 ;
	else if ( rl_rg01_en )
		rl_rg01 <= rl_rg01_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg02_t_c1 = ( rl_we01 & rl_d01 [125] ) ;
	rl_rg02_t_c2 = ( rl_we02 & rl_d02 [125] ) ;
	rl_rg02_t = ( ( { 9{ rl_rg02_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg02_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg02_en = ( rl_rg02_t_c1 | rl_rg02_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg02 <= 9'h000 ;
	else if ( rl_rg02_en )
		rl_rg02 <= rl_rg02_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg03_t_c1 = ( rl_we01 & rl_d01 [124] ) ;
	rl_rg03_t_c2 = ( rl_we02 & rl_d02 [124] ) ;
	rl_rg03_t = ( ( { 9{ rl_rg03_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg03_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg03_en = ( rl_rg03_t_c1 | rl_rg03_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg03 <= 9'h000 ;
	else if ( rl_rg03_en )
		rl_rg03 <= rl_rg03_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg04_t_c1 = ( rl_we01 & rl_d01 [123] ) ;
	rl_rg04_t_c2 = ( rl_we02 & rl_d02 [123] ) ;
	rl_rg04_t = ( ( { 9{ rl_rg04_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg04_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg04_en = ( rl_rg04_t_c1 | rl_rg04_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg04 <= 9'h000 ;
	else if ( rl_rg04_en )
		rl_rg04 <= rl_rg04_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg05_t_c1 = ( rl_we01 & rl_d01 [122] ) ;
	rl_rg05_t_c2 = ( rl_we02 & rl_d02 [122] ) ;
	rl_rg05_t = ( ( { 9{ rl_rg05_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg05_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg05_en = ( rl_rg05_t_c1 | rl_rg05_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg05 <= 9'h000 ;
	else if ( rl_rg05_en )
		rl_rg05 <= rl_rg05_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg06_t_c1 = ( rl_we01 & rl_d01 [121] ) ;
	rl_rg06_t_c2 = ( rl_we02 & rl_d02 [121] ) ;
	rl_rg06_t = ( ( { 9{ rl_rg06_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg06_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg06_en = ( rl_rg06_t_c1 | rl_rg06_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg06 <= 9'h000 ;
	else if ( rl_rg06_en )
		rl_rg06 <= rl_rg06_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg07_t_c1 = ( rl_we01 & rl_d01 [120] ) ;
	rl_rg07_t_c2 = ( rl_we02 & rl_d02 [120] ) ;
	rl_rg07_t = ( ( { 9{ rl_rg07_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg07_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg07_en = ( rl_rg07_t_c1 | rl_rg07_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg07 <= 9'h000 ;
	else if ( rl_rg07_en )
		rl_rg07 <= rl_rg07_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg08_t_c1 = ( rl_we01 & rl_d01 [119] ) ;
	rl_rg08_t_c2 = ( rl_we02 & rl_d02 [119] ) ;
	rl_rg08_t = ( ( { 9{ rl_rg08_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg08_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg08_en = ( rl_rg08_t_c1 | rl_rg08_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg08 <= 9'h000 ;
	else if ( rl_rg08_en )
		rl_rg08 <= rl_rg08_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg09_t_c1 = ( rl_we01 & rl_d01 [118] ) ;
	rl_rg09_t_c2 = ( rl_we02 & rl_d02 [118] ) ;
	rl_rg09_t = ( ( { 9{ rl_rg09_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg09_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg09_en = ( rl_rg09_t_c1 | rl_rg09_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg09 <= 9'h000 ;
	else if ( rl_rg09_en )
		rl_rg09 <= rl_rg09_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg10_t_c1 = ( rl_we01 & rl_d01 [117] ) ;
	rl_rg10_t_c2 = ( rl_we02 & rl_d02 [117] ) ;
	rl_rg10_t = ( ( { 9{ rl_rg10_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg10_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg10_en = ( rl_rg10_t_c1 | rl_rg10_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg10 <= 9'h000 ;
	else if ( rl_rg10_en )
		rl_rg10 <= rl_rg10_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg11_t_c1 = ( rl_we01 & rl_d01 [116] ) ;
	rl_rg11_t_c2 = ( rl_we02 & rl_d02 [116] ) ;
	rl_rg11_t = ( ( { 9{ rl_rg11_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg11_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg11_en = ( rl_rg11_t_c1 | rl_rg11_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg11 <= 9'h000 ;
	else if ( rl_rg11_en )
		rl_rg11 <= rl_rg11_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg12_t_c1 = ( rl_we01 & rl_d01 [115] ) ;
	rl_rg12_t_c2 = ( rl_we02 & rl_d02 [115] ) ;
	rl_rg12_t = ( ( { 9{ rl_rg12_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg12_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg12_en = ( rl_rg12_t_c1 | rl_rg12_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg12 <= 9'h000 ;
	else if ( rl_rg12_en )
		rl_rg12 <= rl_rg12_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg13_t_c1 = ( rl_we01 & rl_d01 [114] ) ;
	rl_rg13_t_c2 = ( rl_we02 & rl_d02 [114] ) ;
	rl_rg13_t = ( ( { 9{ rl_rg13_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg13_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg13_en = ( rl_rg13_t_c1 | rl_rg13_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg13 <= 9'h000 ;
	else if ( rl_rg13_en )
		rl_rg13 <= rl_rg13_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg14_t_c1 = ( rl_we01 & rl_d01 [113] ) ;
	rl_rg14_t_c2 = ( rl_we02 & rl_d02 [113] ) ;
	rl_rg14_t = ( ( { 9{ rl_rg14_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg14_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg14_en = ( rl_rg14_t_c1 | rl_rg14_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg14 <= 9'h000 ;
	else if ( rl_rg14_en )
		rl_rg14 <= rl_rg14_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg15_t_c1 = ( rl_we01 & rl_d01 [112] ) ;
	rl_rg15_t_c2 = ( rl_we02 & rl_d02 [112] ) ;
	rl_rg15_t = ( ( { 9{ rl_rg15_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg15_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg15_en = ( rl_rg15_t_c1 | rl_rg15_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg15 <= 9'h000 ;
	else if ( rl_rg15_en )
		rl_rg15 <= rl_rg15_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg16_t_c1 = ( rl_we01 & rl_d01 [111] ) ;
	rl_rg16_t_c2 = ( rl_we02 & rl_d02 [111] ) ;
	rl_rg16_t = ( ( { 9{ rl_rg16_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg16_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg16_en = ( rl_rg16_t_c1 | rl_rg16_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg16 <= 9'h000 ;
	else if ( rl_rg16_en )
		rl_rg16 <= rl_rg16_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg17_t_c1 = ( rl_we01 & rl_d01 [110] ) ;
	rl_rg17_t_c2 = ( rl_we02 & rl_d02 [110] ) ;
	rl_rg17_t = ( ( { 9{ rl_rg17_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg17_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg17_en = ( rl_rg17_t_c1 | rl_rg17_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg17 <= 9'h000 ;
	else if ( rl_rg17_en )
		rl_rg17 <= rl_rg17_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg18_t_c1 = ( rl_we01 & rl_d01 [109] ) ;
	rl_rg18_t_c2 = ( rl_we02 & rl_d02 [109] ) ;
	rl_rg18_t = ( ( { 9{ rl_rg18_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg18_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg18_en = ( rl_rg18_t_c1 | rl_rg18_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg18 <= 9'h000 ;
	else if ( rl_rg18_en )
		rl_rg18 <= rl_rg18_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg19_t_c1 = ( rl_we01 & rl_d01 [108] ) ;
	rl_rg19_t_c2 = ( rl_we02 & rl_d02 [108] ) ;
	rl_rg19_t = ( ( { 9{ rl_rg19_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg19_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg19_en = ( rl_rg19_t_c1 | rl_rg19_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg19 <= 9'h000 ;
	else if ( rl_rg19_en )
		rl_rg19 <= rl_rg19_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg20_t_c1 = ( rl_we01 & rl_d01 [107] ) ;
	rl_rg20_t_c2 = ( rl_we02 & rl_d02 [107] ) ;
	rl_rg20_t = ( ( { 9{ rl_rg20_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg20_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg20_en = ( rl_rg20_t_c1 | rl_rg20_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg20 <= 9'h000 ;
	else if ( rl_rg20_en )
		rl_rg20 <= rl_rg20_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg21_t_c1 = ( rl_we01 & rl_d01 [106] ) ;
	rl_rg21_t_c2 = ( rl_we02 & rl_d02 [106] ) ;
	rl_rg21_t = ( ( { 9{ rl_rg21_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg21_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg21_en = ( rl_rg21_t_c1 | rl_rg21_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg21 <= 9'h000 ;
	else if ( rl_rg21_en )
		rl_rg21 <= rl_rg21_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg22_t_c1 = ( rl_we01 & rl_d01 [105] ) ;
	rl_rg22_t_c2 = ( rl_we02 & rl_d02 [105] ) ;
	rl_rg22_t = ( ( { 9{ rl_rg22_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg22_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg22_en = ( rl_rg22_t_c1 | rl_rg22_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg22 <= 9'h000 ;
	else if ( rl_rg22_en )
		rl_rg22 <= rl_rg22_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg23_t_c1 = ( rl_we01 & rl_d01 [104] ) ;
	rl_rg23_t_c2 = ( rl_we02 & rl_d02 [104] ) ;
	rl_rg23_t = ( ( { 9{ rl_rg23_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg23_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg23_en = ( rl_rg23_t_c1 | rl_rg23_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg23 <= 9'h000 ;
	else if ( rl_rg23_en )
		rl_rg23 <= rl_rg23_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg24_t_c1 = ( rl_we01 & rl_d01 [103] ) ;
	rl_rg24_t_c2 = ( rl_we02 & rl_d02 [103] ) ;
	rl_rg24_t = ( ( { 9{ rl_rg24_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg24_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg24_en = ( rl_rg24_t_c1 | rl_rg24_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg24 <= 9'h000 ;
	else if ( rl_rg24_en )
		rl_rg24 <= rl_rg24_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg25_t_c1 = ( rl_we01 & rl_d01 [102] ) ;
	rl_rg25_t_c2 = ( rl_we02 & rl_d02 [102] ) ;
	rl_rg25_t = ( ( { 9{ rl_rg25_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg25_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg25_en = ( rl_rg25_t_c1 | rl_rg25_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg25 <= 9'h000 ;
	else if ( rl_rg25_en )
		rl_rg25 <= rl_rg25_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg26_t_c1 = ( rl_we01 & rl_d01 [101] ) ;
	rl_rg26_t_c2 = ( rl_we02 & rl_d02 [101] ) ;
	rl_rg26_t = ( ( { 9{ rl_rg26_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg26_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg26_en = ( rl_rg26_t_c1 | rl_rg26_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg26 <= 9'h000 ;
	else if ( rl_rg26_en )
		rl_rg26 <= rl_rg26_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg27_t_c1 = ( rl_we01 & rl_d01 [100] ) ;
	rl_rg27_t_c2 = ( rl_we02 & rl_d02 [100] ) ;
	rl_rg27_t = ( ( { 9{ rl_rg27_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg27_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg27_en = ( rl_rg27_t_c1 | rl_rg27_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg27 <= 9'h000 ;
	else if ( rl_rg27_en )
		rl_rg27 <= rl_rg27_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg28_t_c1 = ( rl_we01 & rl_d01 [99] ) ;
	rl_rg28_t_c2 = ( rl_we02 & rl_d02 [99] ) ;
	rl_rg28_t = ( ( { 9{ rl_rg28_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg28_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg28_en = ( rl_rg28_t_c1 | rl_rg28_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg28 <= 9'h000 ;
	else if ( rl_rg28_en )
		rl_rg28 <= rl_rg28_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg29_t_c1 = ( rl_we01 & rl_d01 [98] ) ;
	rl_rg29_t_c2 = ( rl_we02 & rl_d02 [98] ) ;
	rl_rg29_t = ( ( { 9{ rl_rg29_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg29_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg29_en = ( rl_rg29_t_c1 | rl_rg29_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg29 <= 9'h000 ;
	else if ( rl_rg29_en )
		rl_rg29 <= rl_rg29_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg30_t_c1 = ( rl_we01 & rl_d01 [97] ) ;
	rl_rg30_t_c2 = ( rl_we02 & rl_d02 [97] ) ;
	rl_rg30_t = ( ( { 9{ rl_rg30_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg30_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg30_en = ( rl_rg30_t_c1 | rl_rg30_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg30 <= 9'h000 ;
	else if ( rl_rg30_en )
		rl_rg30 <= rl_rg30_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg31_t_c1 = ( rl_we01 & rl_d01 [96] ) ;
	rl_rg31_t_c2 = ( rl_we02 & rl_d02 [96] ) ;
	rl_rg31_t = ( ( { 9{ rl_rg31_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg31_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg31_en = ( rl_rg31_t_c1 | rl_rg31_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg31 <= 9'h000 ;
	else if ( rl_rg31_en )
		rl_rg31 <= rl_rg31_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg32_t_c1 = ( rl_we01 & rl_d01 [95] ) ;
	rl_rg32_t_c2 = ( rl_we02 & rl_d02 [95] ) ;
	rl_rg32_t = ( ( { 9{ rl_rg32_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg32_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg32_en = ( rl_rg32_t_c1 | rl_rg32_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg32 <= 9'h000 ;
	else if ( rl_rg32_en )
		rl_rg32 <= rl_rg32_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg33_t_c1 = ( rl_we01 & rl_d01 [94] ) ;
	rl_rg33_t_c2 = ( rl_we02 & rl_d02 [94] ) ;
	rl_rg33_t = ( ( { 9{ rl_rg33_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg33_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg33_en = ( rl_rg33_t_c1 | rl_rg33_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg33 <= 9'h000 ;
	else if ( rl_rg33_en )
		rl_rg33 <= rl_rg33_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg34_t_c1 = ( rl_we01 & rl_d01 [93] ) ;
	rl_rg34_t_c2 = ( rl_we02 & rl_d02 [93] ) ;
	rl_rg34_t = ( ( { 9{ rl_rg34_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg34_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg34_en = ( rl_rg34_t_c1 | rl_rg34_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg34 <= 9'h000 ;
	else if ( rl_rg34_en )
		rl_rg34 <= rl_rg34_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg35_t_c1 = ( rl_we01 & rl_d01 [92] ) ;
	rl_rg35_t_c2 = ( rl_we02 & rl_d02 [92] ) ;
	rl_rg35_t = ( ( { 9{ rl_rg35_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg35_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg35_en = ( rl_rg35_t_c1 | rl_rg35_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg35 <= 9'h000 ;
	else if ( rl_rg35_en )
		rl_rg35 <= rl_rg35_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg36_t_c1 = ( rl_we01 & rl_d01 [91] ) ;
	rl_rg36_t_c2 = ( rl_we02 & rl_d02 [91] ) ;
	rl_rg36_t = ( ( { 9{ rl_rg36_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg36_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg36_en = ( rl_rg36_t_c1 | rl_rg36_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg36 <= 9'h000 ;
	else if ( rl_rg36_en )
		rl_rg36 <= rl_rg36_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg37_t_c1 = ( rl_we01 & rl_d01 [90] ) ;
	rl_rg37_t_c2 = ( rl_we02 & rl_d02 [90] ) ;
	rl_rg37_t = ( ( { 9{ rl_rg37_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg37_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg37_en = ( rl_rg37_t_c1 | rl_rg37_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg37 <= 9'h000 ;
	else if ( rl_rg37_en )
		rl_rg37 <= rl_rg37_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg38_t_c1 = ( rl_we01 & rl_d01 [89] ) ;
	rl_rg38_t_c2 = ( rl_we02 & rl_d02 [89] ) ;
	rl_rg38_t = ( ( { 9{ rl_rg38_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg38_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg38_en = ( rl_rg38_t_c1 | rl_rg38_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg38 <= 9'h000 ;
	else if ( rl_rg38_en )
		rl_rg38 <= rl_rg38_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg39_t_c1 = ( rl_we01 & rl_d01 [88] ) ;
	rl_rg39_t_c2 = ( rl_we02 & rl_d02 [88] ) ;
	rl_rg39_t = ( ( { 9{ rl_rg39_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg39_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg39_en = ( rl_rg39_t_c1 | rl_rg39_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg39 <= 9'h000 ;
	else if ( rl_rg39_en )
		rl_rg39 <= rl_rg39_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg40_t_c1 = ( rl_we01 & rl_d01 [87] ) ;
	rl_rg40_t_c2 = ( rl_we02 & rl_d02 [87] ) ;
	rl_rg40_t = ( ( { 9{ rl_rg40_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg40_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg40_en = ( rl_rg40_t_c1 | rl_rg40_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg40 <= 9'h000 ;
	else if ( rl_rg40_en )
		rl_rg40 <= rl_rg40_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg41_t_c1 = ( rl_we01 & rl_d01 [86] ) ;
	rl_rg41_t_c2 = ( rl_we02 & rl_d02 [86] ) ;
	rl_rg41_t = ( ( { 9{ rl_rg41_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg41_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg41_en = ( rl_rg41_t_c1 | rl_rg41_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg41 <= 9'h000 ;
	else if ( rl_rg41_en )
		rl_rg41 <= rl_rg41_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg42_t_c1 = ( rl_we01 & rl_d01 [85] ) ;
	rl_rg42_t_c2 = ( rl_we02 & rl_d02 [85] ) ;
	rl_rg42_t = ( ( { 9{ rl_rg42_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg42_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg42_en = ( rl_rg42_t_c1 | rl_rg42_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg42 <= 9'h000 ;
	else if ( rl_rg42_en )
		rl_rg42 <= rl_rg42_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg43_t_c1 = ( rl_we01 & rl_d01 [84] ) ;
	rl_rg43_t_c2 = ( rl_we02 & rl_d02 [84] ) ;
	rl_rg43_t = ( ( { 9{ rl_rg43_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg43_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg43_en = ( rl_rg43_t_c1 | rl_rg43_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg43 <= 9'h000 ;
	else if ( rl_rg43_en )
		rl_rg43 <= rl_rg43_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg44_t_c1 = ( rl_we01 & rl_d01 [83] ) ;
	rl_rg44_t_c2 = ( rl_we02 & rl_d02 [83] ) ;
	rl_rg44_t = ( ( { 9{ rl_rg44_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg44_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg44_en = ( rl_rg44_t_c1 | rl_rg44_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg44 <= 9'h000 ;
	else if ( rl_rg44_en )
		rl_rg44 <= rl_rg44_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg45_t_c1 = ( rl_we01 & rl_d01 [82] ) ;
	rl_rg45_t_c2 = ( rl_we02 & rl_d02 [82] ) ;
	rl_rg45_t = ( ( { 9{ rl_rg45_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg45_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg45_en = ( rl_rg45_t_c1 | rl_rg45_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg45 <= 9'h000 ;
	else if ( rl_rg45_en )
		rl_rg45 <= rl_rg45_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg46_t_c1 = ( rl_we01 & rl_d01 [81] ) ;
	rl_rg46_t_c2 = ( rl_we02 & rl_d02 [81] ) ;
	rl_rg46_t = ( ( { 9{ rl_rg46_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg46_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg46_en = ( rl_rg46_t_c1 | rl_rg46_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg46 <= 9'h000 ;
	else if ( rl_rg46_en )
		rl_rg46 <= rl_rg46_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg47_t_c1 = ( rl_we01 & rl_d01 [80] ) ;
	rl_rg47_t_c2 = ( rl_we02 & rl_d02 [80] ) ;
	rl_rg47_t = ( ( { 9{ rl_rg47_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg47_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg47_en = ( rl_rg47_t_c1 | rl_rg47_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg47 <= 9'h000 ;
	else if ( rl_rg47_en )
		rl_rg47 <= rl_rg47_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg48_t_c1 = ( rl_we01 & rl_d01 [79] ) ;
	rl_rg48_t_c2 = ( rl_we02 & rl_d02 [79] ) ;
	rl_rg48_t = ( ( { 9{ rl_rg48_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg48_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg48_en = ( rl_rg48_t_c1 | rl_rg48_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg48 <= 9'h000 ;
	else if ( rl_rg48_en )
		rl_rg48 <= rl_rg48_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg49_t_c1 = ( rl_we01 & rl_d01 [78] ) ;
	rl_rg49_t_c2 = ( rl_we02 & rl_d02 [78] ) ;
	rl_rg49_t = ( ( { 9{ rl_rg49_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg49_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg49_en = ( rl_rg49_t_c1 | rl_rg49_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg49 <= 9'h000 ;
	else if ( rl_rg49_en )
		rl_rg49 <= rl_rg49_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg50_t_c1 = ( rl_we01 & rl_d01 [77] ) ;
	rl_rg50_t_c2 = ( rl_we02 & rl_d02 [77] ) ;
	rl_rg50_t = ( ( { 9{ rl_rg50_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg50_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg50_en = ( rl_rg50_t_c1 | rl_rg50_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg50 <= 9'h000 ;
	else if ( rl_rg50_en )
		rl_rg50 <= rl_rg50_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg51_t_c1 = ( rl_we01 & rl_d01 [76] ) ;
	rl_rg51_t_c2 = ( rl_we02 & rl_d02 [76] ) ;
	rl_rg51_t = ( ( { 9{ rl_rg51_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg51_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg51_en = ( rl_rg51_t_c1 | rl_rg51_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg51 <= 9'h000 ;
	else if ( rl_rg51_en )
		rl_rg51 <= rl_rg51_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg52_t_c1 = ( rl_we01 & rl_d01 [75] ) ;
	rl_rg52_t_c2 = ( rl_we02 & rl_d02 [75] ) ;
	rl_rg52_t = ( ( { 9{ rl_rg52_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg52_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg52_en = ( rl_rg52_t_c1 | rl_rg52_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg52 <= 9'h000 ;
	else if ( rl_rg52_en )
		rl_rg52 <= rl_rg52_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg53_t_c1 = ( rl_we01 & rl_d01 [74] ) ;
	rl_rg53_t_c2 = ( rl_we02 & rl_d02 [74] ) ;
	rl_rg53_t = ( ( { 9{ rl_rg53_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg53_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg53_en = ( rl_rg53_t_c1 | rl_rg53_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg53 <= 9'h000 ;
	else if ( rl_rg53_en )
		rl_rg53 <= rl_rg53_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg54_t_c1 = ( rl_we01 & rl_d01 [73] ) ;
	rl_rg54_t_c2 = ( rl_we02 & rl_d02 [73] ) ;
	rl_rg54_t = ( ( { 9{ rl_rg54_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg54_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg54_en = ( rl_rg54_t_c1 | rl_rg54_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg54 <= 9'h000 ;
	else if ( rl_rg54_en )
		rl_rg54 <= rl_rg54_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg55_t_c1 = ( rl_we01 & rl_d01 [72] ) ;
	rl_rg55_t_c2 = ( rl_we02 & rl_d02 [72] ) ;
	rl_rg55_t = ( ( { 9{ rl_rg55_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg55_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg55_en = ( rl_rg55_t_c1 | rl_rg55_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg55 <= 9'h000 ;
	else if ( rl_rg55_en )
		rl_rg55 <= rl_rg55_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg56_t_c1 = ( rl_we01 & rl_d01 [71] ) ;
	rl_rg56_t_c2 = ( rl_we02 & rl_d02 [71] ) ;
	rl_rg56_t = ( ( { 9{ rl_rg56_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg56_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg56_en = ( rl_rg56_t_c1 | rl_rg56_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg56 <= 9'h000 ;
	else if ( rl_rg56_en )
		rl_rg56 <= rl_rg56_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg57_t_c1 = ( rl_we01 & rl_d01 [70] ) ;
	rl_rg57_t_c2 = ( rl_we02 & rl_d02 [70] ) ;
	rl_rg57_t = ( ( { 9{ rl_rg57_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg57_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg57_en = ( rl_rg57_t_c1 | rl_rg57_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg57 <= 9'h000 ;
	else if ( rl_rg57_en )
		rl_rg57 <= rl_rg57_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg58_t_c1 = ( rl_we01 & rl_d01 [69] ) ;
	rl_rg58_t_c2 = ( rl_we02 & rl_d02 [69] ) ;
	rl_rg58_t = ( ( { 9{ rl_rg58_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg58_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg58_en = ( rl_rg58_t_c1 | rl_rg58_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg58 <= 9'h000 ;
	else if ( rl_rg58_en )
		rl_rg58 <= rl_rg58_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg59_t_c1 = ( rl_we01 & rl_d01 [68] ) ;
	rl_rg59_t_c2 = ( rl_we02 & rl_d02 [68] ) ;
	rl_rg59_t = ( ( { 9{ rl_rg59_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg59_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg59_en = ( rl_rg59_t_c1 | rl_rg59_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg59 <= 9'h000 ;
	else if ( rl_rg59_en )
		rl_rg59 <= rl_rg59_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg60_t_c1 = ( rl_we01 & rl_d01 [67] ) ;
	rl_rg60_t_c2 = ( rl_we02 & rl_d02 [67] ) ;
	rl_rg60_t = ( ( { 9{ rl_rg60_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg60_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg60_en = ( rl_rg60_t_c1 | rl_rg60_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg60 <= 9'h000 ;
	else if ( rl_rg60_en )
		rl_rg60 <= rl_rg60_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg61_t_c1 = ( rl_we01 & rl_d01 [66] ) ;
	rl_rg61_t_c2 = ( rl_we02 & rl_d02 [66] ) ;
	rl_rg61_t = ( ( { 9{ rl_rg61_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg61_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg61_en = ( rl_rg61_t_c1 | rl_rg61_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg61 <= 9'h000 ;
	else if ( rl_rg61_en )
		rl_rg61 <= rl_rg61_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg62_t_c1 = ( rl_we01 & rl_d01 [65] ) ;
	rl_rg62_t_c2 = ( rl_we02 & rl_d02 [65] ) ;
	rl_rg62_t = ( ( { 9{ rl_rg62_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg62_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg62_en = ( rl_rg62_t_c1 | rl_rg62_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg62 <= 9'h000 ;
	else if ( rl_rg62_en )
		rl_rg62 <= rl_rg62_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg63_t_c1 = ( rl_we01 & rl_d01 [64] ) ;
	rl_rg63_t_c2 = ( rl_we02 & rl_d02 [64] ) ;
	rl_rg63_t = ( ( { 9{ rl_rg63_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg63_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg63_en = ( rl_rg63_t_c1 | rl_rg63_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg63 <= 9'h000 ;
	else if ( rl_rg63_en )
		rl_rg63 <= rl_rg63_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg64_t_c1 = ( rl_we01 & rl_d01 [63] ) ;
	rl_rg64_t_c2 = ( rl_we02 & rl_d02 [63] ) ;
	rl_rg64_t = ( ( { 9{ rl_rg64_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg64_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg64_en = ( rl_rg64_t_c1 | rl_rg64_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg64 <= 9'h000 ;
	else if ( rl_rg64_en )
		rl_rg64 <= rl_rg64_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg65_t_c1 = ( rl_we01 & rl_d01 [62] ) ;
	rl_rg65_t_c2 = ( rl_we02 & rl_d02 [62] ) ;
	rl_rg65_t = ( ( { 9{ rl_rg65_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg65_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg65_en = ( rl_rg65_t_c1 | rl_rg65_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg65 <= 9'h000 ;
	else if ( rl_rg65_en )
		rl_rg65 <= rl_rg65_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg66_t_c1 = ( rl_we01 & rl_d01 [61] ) ;
	rl_rg66_t_c2 = ( rl_we02 & rl_d02 [61] ) ;
	rl_rg66_t = ( ( { 9{ rl_rg66_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg66_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg66_en = ( rl_rg66_t_c1 | rl_rg66_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg66 <= 9'h000 ;
	else if ( rl_rg66_en )
		rl_rg66 <= rl_rg66_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg67_t_c1 = ( rl_we01 & rl_d01 [60] ) ;
	rl_rg67_t_c2 = ( rl_we02 & rl_d02 [60] ) ;
	rl_rg67_t = ( ( { 9{ rl_rg67_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg67_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg67_en = ( rl_rg67_t_c1 | rl_rg67_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg67 <= 9'h000 ;
	else if ( rl_rg67_en )
		rl_rg67 <= rl_rg67_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg68_t_c1 = ( rl_we01 & rl_d01 [59] ) ;
	rl_rg68_t_c2 = ( rl_we02 & rl_d02 [59] ) ;
	rl_rg68_t = ( ( { 9{ rl_rg68_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg68_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg68_en = ( rl_rg68_t_c1 | rl_rg68_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg68 <= 9'h000 ;
	else if ( rl_rg68_en )
		rl_rg68 <= rl_rg68_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg69_t_c1 = ( rl_we01 & rl_d01 [58] ) ;
	rl_rg69_t_c2 = ( rl_we02 & rl_d02 [58] ) ;
	rl_rg69_t = ( ( { 9{ rl_rg69_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg69_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg69_en = ( rl_rg69_t_c1 | rl_rg69_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg69 <= 9'h000 ;
	else if ( rl_rg69_en )
		rl_rg69 <= rl_rg69_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg70_t_c1 = ( rl_we01 & rl_d01 [57] ) ;
	rl_rg70_t_c2 = ( rl_we02 & rl_d02 [57] ) ;
	rl_rg70_t = ( ( { 9{ rl_rg70_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg70_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg70_en = ( rl_rg70_t_c1 | rl_rg70_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg70 <= 9'h000 ;
	else if ( rl_rg70_en )
		rl_rg70 <= rl_rg70_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg71_t_c1 = ( rl_we01 & rl_d01 [56] ) ;
	rl_rg71_t_c2 = ( rl_we02 & rl_d02 [56] ) ;
	rl_rg71_t = ( ( { 9{ rl_rg71_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg71_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg71_en = ( rl_rg71_t_c1 | rl_rg71_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg71 <= 9'h000 ;
	else if ( rl_rg71_en )
		rl_rg71 <= rl_rg71_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg72_t_c1 = ( rl_we01 & rl_d01 [55] ) ;
	rl_rg72_t_c2 = ( rl_we02 & rl_d02 [55] ) ;
	rl_rg72_t = ( ( { 9{ rl_rg72_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg72_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg72_en = ( rl_rg72_t_c1 | rl_rg72_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg72 <= 9'h000 ;
	else if ( rl_rg72_en )
		rl_rg72 <= rl_rg72_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg73_t_c1 = ( rl_we01 & rl_d01 [54] ) ;
	rl_rg73_t_c2 = ( rl_we02 & rl_d02 [54] ) ;
	rl_rg73_t = ( ( { 9{ rl_rg73_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg73_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg73_en = ( rl_rg73_t_c1 | rl_rg73_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg73 <= 9'h000 ;
	else if ( rl_rg73_en )
		rl_rg73 <= rl_rg73_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg74_t_c1 = ( rl_we01 & rl_d01 [53] ) ;
	rl_rg74_t_c2 = ( rl_we02 & rl_d02 [53] ) ;
	rl_rg74_t = ( ( { 9{ rl_rg74_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg74_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg74_en = ( rl_rg74_t_c1 | rl_rg74_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg74 <= 9'h000 ;
	else if ( rl_rg74_en )
		rl_rg74 <= rl_rg74_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg75_t_c1 = ( rl_we01 & rl_d01 [52] ) ;
	rl_rg75_t_c2 = ( rl_we02 & rl_d02 [52] ) ;
	rl_rg75_t = ( ( { 9{ rl_rg75_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg75_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg75_en = ( rl_rg75_t_c1 | rl_rg75_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg75 <= 9'h000 ;
	else if ( rl_rg75_en )
		rl_rg75 <= rl_rg75_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg76_t_c1 = ( rl_we01 & rl_d01 [51] ) ;
	rl_rg76_t_c2 = ( rl_we02 & rl_d02 [51] ) ;
	rl_rg76_t = ( ( { 9{ rl_rg76_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg76_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg76_en = ( rl_rg76_t_c1 | rl_rg76_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg76 <= 9'h000 ;
	else if ( rl_rg76_en )
		rl_rg76 <= rl_rg76_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg77_t_c1 = ( rl_we01 & rl_d01 [50] ) ;
	rl_rg77_t_c2 = ( rl_we02 & rl_d02 [50] ) ;
	rl_rg77_t = ( ( { 9{ rl_rg77_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg77_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg77_en = ( rl_rg77_t_c1 | rl_rg77_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg77 <= 9'h000 ;
	else if ( rl_rg77_en )
		rl_rg77 <= rl_rg77_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg78_t_c1 = ( rl_we01 & rl_d01 [49] ) ;
	rl_rg78_t_c2 = ( rl_we02 & rl_d02 [49] ) ;
	rl_rg78_t = ( ( { 9{ rl_rg78_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg78_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg78_en = ( rl_rg78_t_c1 | rl_rg78_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg78 <= 9'h000 ;
	else if ( rl_rg78_en )
		rl_rg78 <= rl_rg78_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg79_t_c1 = ( rl_we01 & rl_d01 [48] ) ;
	rl_rg79_t_c2 = ( rl_we02 & rl_d02 [48] ) ;
	rl_rg79_t = ( ( { 9{ rl_rg79_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg79_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg79_en = ( rl_rg79_t_c1 | rl_rg79_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg79 <= 9'h000 ;
	else if ( rl_rg79_en )
		rl_rg79 <= rl_rg79_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg80_t_c1 = ( rl_we01 & rl_d01 [47] ) ;
	rl_rg80_t_c2 = ( rl_we02 & rl_d02 [47] ) ;
	rl_rg80_t = ( ( { 9{ rl_rg80_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg80_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg80_en = ( rl_rg80_t_c1 | rl_rg80_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg80 <= 9'h000 ;
	else if ( rl_rg80_en )
		rl_rg80 <= rl_rg80_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg81_t_c1 = ( rl_we01 & rl_d01 [46] ) ;
	rl_rg81_t_c2 = ( rl_we02 & rl_d02 [46] ) ;
	rl_rg81_t = ( ( { 9{ rl_rg81_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg81_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg81_en = ( rl_rg81_t_c1 | rl_rg81_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg81 <= 9'h000 ;
	else if ( rl_rg81_en )
		rl_rg81 <= rl_rg81_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg82_t_c1 = ( rl_we01 & rl_d01 [45] ) ;
	rl_rg82_t_c2 = ( rl_we02 & rl_d02 [45] ) ;
	rl_rg82_t = ( ( { 9{ rl_rg82_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg82_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg82_en = ( rl_rg82_t_c1 | rl_rg82_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg82 <= 9'h000 ;
	else if ( rl_rg82_en )
		rl_rg82 <= rl_rg82_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg83_t_c1 = ( rl_we01 & rl_d01 [44] ) ;
	rl_rg83_t_c2 = ( rl_we02 & rl_d02 [44] ) ;
	rl_rg83_t = ( ( { 9{ rl_rg83_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg83_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg83_en = ( rl_rg83_t_c1 | rl_rg83_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg83 <= 9'h000 ;
	else if ( rl_rg83_en )
		rl_rg83 <= rl_rg83_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg84_t_c1 = ( rl_we01 & rl_d01 [43] ) ;
	rl_rg84_t_c2 = ( rl_we02 & rl_d02 [43] ) ;
	rl_rg84_t = ( ( { 9{ rl_rg84_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg84_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg84_en = ( rl_rg84_t_c1 | rl_rg84_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg84 <= 9'h000 ;
	else if ( rl_rg84_en )
		rl_rg84 <= rl_rg84_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg85_t_c1 = ( rl_we01 & rl_d01 [42] ) ;
	rl_rg85_t_c2 = ( rl_we02 & rl_d02 [42] ) ;
	rl_rg85_t = ( ( { 9{ rl_rg85_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg85_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg85_en = ( rl_rg85_t_c1 | rl_rg85_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg85 <= 9'h000 ;
	else if ( rl_rg85_en )
		rl_rg85 <= rl_rg85_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg86_t_c1 = ( rl_we01 & rl_d01 [41] ) ;
	rl_rg86_t_c2 = ( rl_we02 & rl_d02 [41] ) ;
	rl_rg86_t = ( ( { 9{ rl_rg86_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg86_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg86_en = ( rl_rg86_t_c1 | rl_rg86_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg86 <= 9'h000 ;
	else if ( rl_rg86_en )
		rl_rg86 <= rl_rg86_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg87_t_c1 = ( rl_we01 & rl_d01 [40] ) ;
	rl_rg87_t_c2 = ( rl_we02 & rl_d02 [40] ) ;
	rl_rg87_t = ( ( { 9{ rl_rg87_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg87_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg87_en = ( rl_rg87_t_c1 | rl_rg87_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg87 <= 9'h000 ;
	else if ( rl_rg87_en )
		rl_rg87 <= rl_rg87_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg88_t_c1 = ( rl_we01 & rl_d01 [39] ) ;
	rl_rg88_t_c2 = ( rl_we02 & rl_d02 [39] ) ;
	rl_rg88_t = ( ( { 9{ rl_rg88_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg88_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg88_en = ( rl_rg88_t_c1 | rl_rg88_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg88 <= 9'h000 ;
	else if ( rl_rg88_en )
		rl_rg88 <= rl_rg88_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg89_t_c1 = ( rl_we01 & rl_d01 [38] ) ;
	rl_rg89_t_c2 = ( rl_we02 & rl_d02 [38] ) ;
	rl_rg89_t = ( ( { 9{ rl_rg89_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg89_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg89_en = ( rl_rg89_t_c1 | rl_rg89_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg89 <= 9'h000 ;
	else if ( rl_rg89_en )
		rl_rg89 <= rl_rg89_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg90_t_c1 = ( rl_we01 & rl_d01 [37] ) ;
	rl_rg90_t_c2 = ( rl_we02 & rl_d02 [37] ) ;
	rl_rg90_t = ( ( { 9{ rl_rg90_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg90_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg90_en = ( rl_rg90_t_c1 | rl_rg90_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg90 <= 9'h000 ;
	else if ( rl_rg90_en )
		rl_rg90 <= rl_rg90_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg91_t_c1 = ( rl_we01 & rl_d01 [36] ) ;
	rl_rg91_t_c2 = ( rl_we02 & rl_d02 [36] ) ;
	rl_rg91_t = ( ( { 9{ rl_rg91_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg91_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg91_en = ( rl_rg91_t_c1 | rl_rg91_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg91 <= 9'h000 ;
	else if ( rl_rg91_en )
		rl_rg91 <= rl_rg91_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg92_t_c1 = ( rl_we01 & rl_d01 [35] ) ;
	rl_rg92_t_c2 = ( rl_we02 & rl_d02 [35] ) ;
	rl_rg92_t = ( ( { 9{ rl_rg92_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg92_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg92_en = ( rl_rg92_t_c1 | rl_rg92_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg92 <= 9'h000 ;
	else if ( rl_rg92_en )
		rl_rg92 <= rl_rg92_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg93_t_c1 = ( rl_we01 & rl_d01 [34] ) ;
	rl_rg93_t_c2 = ( rl_we02 & rl_d02 [34] ) ;
	rl_rg93_t = ( ( { 9{ rl_rg93_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg93_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg93_en = ( rl_rg93_t_c1 | rl_rg93_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg93 <= 9'h000 ;
	else if ( rl_rg93_en )
		rl_rg93 <= rl_rg93_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg94_t_c1 = ( rl_we01 & rl_d01 [33] ) ;
	rl_rg94_t_c2 = ( rl_we02 & rl_d02 [33] ) ;
	rl_rg94_t = ( ( { 9{ rl_rg94_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg94_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg94_en = ( rl_rg94_t_c1 | rl_rg94_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg94 <= 9'h000 ;
	else if ( rl_rg94_en )
		rl_rg94 <= rl_rg94_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg95_t_c1 = ( rl_we01 & rl_d01 [32] ) ;
	rl_rg95_t_c2 = ( rl_we02 & rl_d02 [32] ) ;
	rl_rg95_t = ( ( { 9{ rl_rg95_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg95_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg95_en = ( rl_rg95_t_c1 | rl_rg95_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg95 <= 9'h000 ;
	else if ( rl_rg95_en )
		rl_rg95 <= rl_rg95_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg96_t_c1 = ( rl_we01 & rl_d01 [31] ) ;
	rl_rg96_t_c2 = ( rl_we02 & rl_d02 [31] ) ;
	rl_rg96_t = ( ( { 9{ rl_rg96_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg96_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg96_en = ( rl_rg96_t_c1 | rl_rg96_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg96 <= 9'h000 ;
	else if ( rl_rg96_en )
		rl_rg96 <= rl_rg96_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg97_t_c1 = ( rl_we01 & rl_d01 [30] ) ;
	rl_rg97_t_c2 = ( rl_we02 & rl_d02 [30] ) ;
	rl_rg97_t = ( ( { 9{ rl_rg97_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg97_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg97_en = ( rl_rg97_t_c1 | rl_rg97_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg97 <= 9'h000 ;
	else if ( rl_rg97_en )
		rl_rg97 <= rl_rg97_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg98_t_c1 = ( rl_we01 & rl_d01 [29] ) ;
	rl_rg98_t_c2 = ( rl_we02 & rl_d02 [29] ) ;
	rl_rg98_t = ( ( { 9{ rl_rg98_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg98_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg98_en = ( rl_rg98_t_c1 | rl_rg98_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg98 <= 9'h000 ;
	else if ( rl_rg98_en )
		rl_rg98 <= rl_rg98_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg99_t_c1 = ( rl_we01 & rl_d01 [28] ) ;
	rl_rg99_t_c2 = ( rl_we02 & rl_d02 [28] ) ;
	rl_rg99_t = ( ( { 9{ rl_rg99_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg99_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg99_en = ( rl_rg99_t_c1 | rl_rg99_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg99 <= 9'h000 ;
	else if ( rl_rg99_en )
		rl_rg99 <= rl_rg99_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg100_t_c1 = ( rl_we01 & rl_d01 [27] ) ;
	rl_rg100_t_c2 = ( rl_we02 & rl_d02 [27] ) ;
	rl_rg100_t = ( ( { 9{ rl_rg100_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg100_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg100_en = ( rl_rg100_t_c1 | rl_rg100_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg100 <= 9'h000 ;
	else if ( rl_rg100_en )
		rl_rg100 <= rl_rg100_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg101_t_c1 = ( rl_we01 & rl_d01 [26] ) ;
	rl_rg101_t_c2 = ( rl_we02 & rl_d02 [26] ) ;
	rl_rg101_t = ( ( { 9{ rl_rg101_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg101_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg101_en = ( rl_rg101_t_c1 | rl_rg101_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg101 <= 9'h000 ;
	else if ( rl_rg101_en )
		rl_rg101 <= rl_rg101_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg102_t_c1 = ( rl_we01 & rl_d01 [25] ) ;
	rl_rg102_t_c2 = ( rl_we02 & rl_d02 [25] ) ;
	rl_rg102_t = ( ( { 9{ rl_rg102_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg102_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg102_en = ( rl_rg102_t_c1 | rl_rg102_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg102 <= 9'h000 ;
	else if ( rl_rg102_en )
		rl_rg102 <= rl_rg102_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg103_t_c1 = ( rl_we01 & rl_d01 [24] ) ;
	rl_rg103_t_c2 = ( rl_we02 & rl_d02 [24] ) ;
	rl_rg103_t = ( ( { 9{ rl_rg103_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg103_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg103_en = ( rl_rg103_t_c1 | rl_rg103_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg103 <= 9'h000 ;
	else if ( rl_rg103_en )
		rl_rg103 <= rl_rg103_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg104_t_c1 = ( rl_we01 & rl_d01 [23] ) ;
	rl_rg104_t_c2 = ( rl_we02 & rl_d02 [23] ) ;
	rl_rg104_t = ( ( { 9{ rl_rg104_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg104_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg104_en = ( rl_rg104_t_c1 | rl_rg104_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg104 <= 9'h000 ;
	else if ( rl_rg104_en )
		rl_rg104 <= rl_rg104_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg105_t_c1 = ( rl_we01 & rl_d01 [22] ) ;
	rl_rg105_t_c2 = ( rl_we02 & rl_d02 [22] ) ;
	rl_rg105_t = ( ( { 9{ rl_rg105_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg105_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg105_en = ( rl_rg105_t_c1 | rl_rg105_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg105 <= 9'h000 ;
	else if ( rl_rg105_en )
		rl_rg105 <= rl_rg105_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg106_t_c1 = ( rl_we01 & rl_d01 [21] ) ;
	rl_rg106_t_c2 = ( rl_we02 & rl_d02 [21] ) ;
	rl_rg106_t = ( ( { 9{ rl_rg106_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg106_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg106_en = ( rl_rg106_t_c1 | rl_rg106_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg106 <= 9'h000 ;
	else if ( rl_rg106_en )
		rl_rg106 <= rl_rg106_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg107_t_c1 = ( rl_we01 & rl_d01 [20] ) ;
	rl_rg107_t_c2 = ( rl_we02 & rl_d02 [20] ) ;
	rl_rg107_t = ( ( { 9{ rl_rg107_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg107_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg107_en = ( rl_rg107_t_c1 | rl_rg107_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg107 <= 9'h000 ;
	else if ( rl_rg107_en )
		rl_rg107 <= rl_rg107_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg108_t_c1 = ( rl_we01 & rl_d01 [19] ) ;
	rl_rg108_t_c2 = ( rl_we02 & rl_d02 [19] ) ;
	rl_rg108_t = ( ( { 9{ rl_rg108_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg108_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg108_en = ( rl_rg108_t_c1 | rl_rg108_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg108 <= 9'h000 ;
	else if ( rl_rg108_en )
		rl_rg108 <= rl_rg108_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg109_t_c1 = ( rl_we01 & rl_d01 [18] ) ;
	rl_rg109_t_c2 = ( rl_we02 & rl_d02 [18] ) ;
	rl_rg109_t = ( ( { 9{ rl_rg109_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg109_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg109_en = ( rl_rg109_t_c1 | rl_rg109_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg109 <= 9'h000 ;
	else if ( rl_rg109_en )
		rl_rg109 <= rl_rg109_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg110_t_c1 = ( rl_we01 & rl_d01 [17] ) ;
	rl_rg110_t_c2 = ( rl_we02 & rl_d02 [17] ) ;
	rl_rg110_t = ( ( { 9{ rl_rg110_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg110_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg110_en = ( rl_rg110_t_c1 | rl_rg110_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg110 <= 9'h000 ;
	else if ( rl_rg110_en )
		rl_rg110 <= rl_rg110_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg111_t_c1 = ( rl_we01 & rl_d01 [16] ) ;
	rl_rg111_t_c2 = ( rl_we02 & rl_d02 [16] ) ;
	rl_rg111_t = ( ( { 9{ rl_rg111_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg111_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg111_en = ( rl_rg111_t_c1 | rl_rg111_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg111 <= 9'h000 ;
	else if ( rl_rg111_en )
		rl_rg111 <= rl_rg111_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg112_t_c1 = ( rl_we01 & rl_d01 [15] ) ;
	rl_rg112_t_c2 = ( rl_we02 & rl_d02 [15] ) ;
	rl_rg112_t = ( ( { 9{ rl_rg112_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg112_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg112_en = ( rl_rg112_t_c1 | rl_rg112_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg112 <= 9'h000 ;
	else if ( rl_rg112_en )
		rl_rg112 <= rl_rg112_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg113_t_c1 = ( rl_we01 & rl_d01 [14] ) ;
	rl_rg113_t_c2 = ( rl_we02 & rl_d02 [14] ) ;
	rl_rg113_t = ( ( { 9{ rl_rg113_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg113_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg113_en = ( rl_rg113_t_c1 | rl_rg113_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg113 <= 9'h000 ;
	else if ( rl_rg113_en )
		rl_rg113 <= rl_rg113_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg114_t_c1 = ( rl_we01 & rl_d01 [13] ) ;
	rl_rg114_t_c2 = ( rl_we02 & rl_d02 [13] ) ;
	rl_rg114_t = ( ( { 9{ rl_rg114_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg114_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg114_en = ( rl_rg114_t_c1 | rl_rg114_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg114 <= 9'h000 ;
	else if ( rl_rg114_en )
		rl_rg114 <= rl_rg114_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg115_t_c1 = ( rl_we01 & rl_d01 [12] ) ;
	rl_rg115_t_c2 = ( rl_we02 & rl_d02 [12] ) ;
	rl_rg115_t = ( ( { 9{ rl_rg115_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg115_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg115_en = ( rl_rg115_t_c1 | rl_rg115_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg115 <= 9'h000 ;
	else if ( rl_rg115_en )
		rl_rg115 <= rl_rg115_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg116_t_c1 = ( rl_we01 & rl_d01 [11] ) ;
	rl_rg116_t_c2 = ( rl_we02 & rl_d02 [11] ) ;
	rl_rg116_t = ( ( { 9{ rl_rg116_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg116_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg116_en = ( rl_rg116_t_c1 | rl_rg116_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg116 <= 9'h000 ;
	else if ( rl_rg116_en )
		rl_rg116 <= rl_rg116_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg117_t_c1 = ( rl_we01 & rl_d01 [10] ) ;
	rl_rg117_t_c2 = ( rl_we02 & rl_d02 [10] ) ;
	rl_rg117_t = ( ( { 9{ rl_rg117_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg117_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg117_en = ( rl_rg117_t_c1 | rl_rg117_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg117 <= 9'h000 ;
	else if ( rl_rg117_en )
		rl_rg117 <= rl_rg117_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg118_t_c1 = ( rl_we01 & rl_d01 [9] ) ;
	rl_rg118_t_c2 = ( rl_we02 & rl_d02 [9] ) ;
	rl_rg118_t = ( ( { 9{ rl_rg118_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg118_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg118_en = ( rl_rg118_t_c1 | rl_rg118_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg118 <= 9'h000 ;
	else if ( rl_rg118_en )
		rl_rg118 <= rl_rg118_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg119_t_c1 = ( rl_we01 & rl_d01 [8] ) ;
	rl_rg119_t_c2 = ( rl_we02 & rl_d02 [8] ) ;
	rl_rg119_t = ( ( { 9{ rl_rg119_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg119_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg119_en = ( rl_rg119_t_c1 | rl_rg119_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg119 <= 9'h000 ;
	else if ( rl_rg119_en )
		rl_rg119 <= rl_rg119_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg120_t_c1 = ( rl_we01 & rl_d01 [7] ) ;
	rl_rg120_t_c2 = ( rl_we02 & rl_d02 [7] ) ;
	rl_rg120_t = ( ( { 9{ rl_rg120_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg120_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg120_en = ( rl_rg120_t_c1 | rl_rg120_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg120 <= 9'h000 ;
	else if ( rl_rg120_en )
		rl_rg120 <= rl_rg120_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg121_t_c1 = ( rl_we01 & rl_d01 [6] ) ;
	rl_rg121_t_c2 = ( rl_we02 & rl_d02 [6] ) ;
	rl_rg121_t = ( ( { 9{ rl_rg121_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg121_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg121_en = ( rl_rg121_t_c1 | rl_rg121_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg121 <= 9'h000 ;
	else if ( rl_rg121_en )
		rl_rg121 <= rl_rg121_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg122_t_c1 = ( rl_we01 & rl_d01 [5] ) ;
	rl_rg122_t_c2 = ( rl_we02 & rl_d02 [5] ) ;
	rl_rg122_t = ( ( { 9{ rl_rg122_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg122_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg122_en = ( rl_rg122_t_c1 | rl_rg122_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg122 <= 9'h000 ;
	else if ( rl_rg122_en )
		rl_rg122 <= rl_rg122_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg123_t_c1 = ( rl_we01 & rl_d01 [4] ) ;
	rl_rg123_t_c2 = ( rl_we02 & rl_d02 [4] ) ;
	rl_rg123_t = ( ( { 9{ rl_rg123_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg123_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg123_en = ( rl_rg123_t_c1 | rl_rg123_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg123 <= 9'h000 ;
	else if ( rl_rg123_en )
		rl_rg123 <= rl_rg123_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg124_t_c1 = ( rl_we01 & rl_d01 [3] ) ;
	rl_rg124_t_c2 = ( rl_we02 & rl_d02 [3] ) ;
	rl_rg124_t = ( ( { 9{ rl_rg124_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg124_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg124_en = ( rl_rg124_t_c1 | rl_rg124_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg124 <= 9'h000 ;
	else if ( rl_rg124_en )
		rl_rg124 <= rl_rg124_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg125_t_c1 = ( rl_we01 & rl_d01 [2] ) ;
	rl_rg125_t_c2 = ( rl_we02 & rl_d02 [2] ) ;
	rl_rg125_t = ( ( { 9{ rl_rg125_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg125_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg125_en = ( rl_rg125_t_c1 | rl_rg125_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg125 <= 9'h000 ;
	else if ( rl_rg125_en )
		rl_rg125 <= rl_rg125_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg126_t_c1 = ( rl_we01 & rl_d01 [1] ) ;
	rl_rg126_t_c2 = ( rl_we02 & rl_d02 [1] ) ;
	rl_rg126_t = ( ( { 9{ rl_rg126_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg126_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg126_en = ( rl_rg126_t_c1 | rl_rg126_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg126 <= 9'h000 ;
	else if ( rl_rg126_en )
		rl_rg126 <= rl_rg126_t ;	// line#=../rle.cpp:23
always @ ( rl_wd02 or rl_d02 or rl_we02 or rl_wd01 or rl_d01 or rl_we01 )	// line#=../rle.cpp:23
	begin
	rl_rg127_t_c1 = ( rl_we01 & rl_d01 [0] ) ;
	rl_rg127_t_c2 = ( rl_we02 & rl_d02 [0] ) ;
	rl_rg127_t = ( ( { 9{ rl_rg127_t_c1 } } & rl_wd01 )
		| ( { 9{ rl_rg127_t_c2 } } & rl_wd02 ) ) ;
	end
assign	rl_rg127_en = ( rl_rg127_t_c1 | rl_rg127_t_c2 ) ;	// line#=../rle.cpp:23
always @ ( posedge clk )	// line#=../rle.cpp:23
	if ( !rst )
		rl_rg127 <= 9'h000 ;
	else if ( rl_rg127_en )
		rl_rg127 <= rl_rg127_t ;	// line#=../rle.cpp:23
assign	CT_06 = ( ( ~|RG_j_k ) & M_432 ) ;	// line#=../rle.cpp:117,118
assign	M_432 = ~|{ ( RG_i [31] & RG_i [0] ) , ~RG_i [0] } ;	// line#=../rle.cpp:117,118,148,149
assign	CT_11 = ( ( ~|{ RG_j_k [31:3] , ~RG_j_k [2:0] } ) & M_432 ) ;	// line#=../rle.cpp:148,149
assign	CT_14 = ( RG_i [31] | ( ~|RG_i [30:6] ) ) ;	// line#=../rle.cpp:61,62
jpeg_CMPS_FL_C2496 #(9) CMPS_FL_C2496_1 ( .CLOCK(clk) ,.RESET(rst) ,.DO(zz_RD1) ,
	.DO_v(CMPS_FL_C2496_1_DO_v) ,.AD_v(U_59) ,.FL_RESET(ST1_07d) ,.DO_t(CMPS_FL_C2496_1_DO_t) );
always @ ( CMPS_FL_C2496_1_DO_t or RG_15_02 )	// line#=../rle.cpp:61,62
	case ( RG_15_02 )
	1'h1 :
		M_01_t1 = ~|CMPS_FL_C2496_1_DO_t ;	// line#=../rle.cpp:61,62
	1'h0 :
		M_01_t1 = 1'h0 ;	// line#=../rle.cpp:61,62
	default :
		M_01_t1 = 1'hx ;
	endcase
assign	CT_16 = ~|{ RG_i_04 [31:7] , ~RG_i_04 [6] , RG_i_04 [5:0] } ;	// line#=../rle.cpp:66,67
assign	CT_17 = ~|rl_rd00 ;	// line#=../rle.cpp:77,78,83,84
always @ ( CT_17 )	// line#=../rle.cpp:77,78
	case ( CT_17 )
	1'h1 :
		JF_08 = 1'h1 ;
	1'h0 :
		JF_08 = 1'h0 ;
	default :
		JF_08 = 1'hx ;
	endcase
always @ ( CT_17 or RG_15_02 )	// line#=../rle.cpp:83,84
	case ( RG_15_02 )
	1'h1 :
		CT_20 = CT_17 ;	// line#=../rle.cpp:83,84
	1'h0 :
		CT_20 = 1'h0 ;	// line#=../rle.cpp:83,84
	default :
		CT_20 = 1'hx ;
	endcase
assign	FL01_01_Leos_all = ( FL01_01_eos & FL01_02_eos ) ;
assign	FL02_01_Leos_all = ( ( ( ( FL02_01_eos & FL02_02_Leos ) & FL02_04_eos ) & 
	FL02_05_eos ) & FL02_06_eos ) ;
assign	FL02_02_Leos_all = ( FL02_02_eos & FL02_03_eos ) ;
assign	FL02_02_rdy = 1'h1 ;
assign	add3u1i1 = RG_03_02 ;	// line#=../rle.cpp:45
assign	add3u1i2 = RG_y_02 [3] ;	// line#=../rle.cpp:45
assign	sub12s_91i1 = zz_RD1 ;	// line#=../rle.cpp:52,53
assign	sub12s_91i2 = RG_previous_dc ;	// line#=../rle.cpp:52
assign	lop8u_11i1 = RG_k ;	// line#=../rle.cpp:109,110
assign	lop8u_11i2 = 6'h24 ;	// line#=../rle.cpp:109,110
assign	incr3u1i1 = RG_j_x_02 [2:0] ;	// line#=../rle.cpp:42
assign	incr32s3i1 = RG_i_05 ;	// line#=../rle.cpp:74
assign	decr8u_71i1 = RG_len_05 [6:0] ;	// line#=../rle.cpp:77,78
assign	incr8u_71i1 = RG_k_05 [5:0] ;	// line#=../rle.cpp:142
assign	incr8u_61i1 = RG_k ;	// line#=../rle.cpp:111
assign	quantized_block_ad01 = { RG_03_02 , RG_y_02 [2:0] } ;	// line#=../rle.cpp:45
always @ ( jpeg_in_a127 or jpeg_in_a126 or jpeg_in_a125 or jpeg_in_a124 or jpeg_in_a123 or 
	jpeg_in_a122 or jpeg_in_a121 or jpeg_in_a120 or jpeg_in_a119 or jpeg_in_a118 or 
	jpeg_in_a117 or jpeg_in_a116 or jpeg_in_a115 or jpeg_in_a114 or jpeg_in_a113 or 
	jpeg_in_a112 or jpeg_in_a111 or jpeg_in_a110 or jpeg_in_a109 or jpeg_in_a108 or 
	jpeg_in_a107 or jpeg_in_a106 or jpeg_in_a105 or jpeg_in_a104 or jpeg_in_a103 or 
	jpeg_in_a102 or jpeg_in_a101 or jpeg_in_a100 or jpeg_in_a99 or jpeg_in_a98 or 
	jpeg_in_a97 or jpeg_in_a96 or jpeg_in_a95 or jpeg_in_a94 or jpeg_in_a93 or 
	jpeg_in_a92 or jpeg_in_a91 or jpeg_in_a90 or jpeg_in_a89 or jpeg_in_a88 or 
	jpeg_in_a87 or jpeg_in_a86 or jpeg_in_a85 or jpeg_in_a84 or jpeg_in_a83 or 
	jpeg_in_a82 or jpeg_in_a81 or jpeg_in_a80 or jpeg_in_a79 or jpeg_in_a78 or 
	jpeg_in_a77 or jpeg_in_a76 or jpeg_in_a75 or jpeg_in_a74 or jpeg_in_a73 or 
	jpeg_in_a72 or jpeg_in_a71 or jpeg_in_a70 or jpeg_in_a69 or jpeg_in_a68 or 
	jpeg_in_a67 or jpeg_in_a66 or jpeg_in_a65 or jpeg_in_a64 or jpeg_in_a63 or 
	jpeg_in_a62 or jpeg_in_a61 or jpeg_in_a60 or jpeg_in_a59 or jpeg_in_a58 or 
	jpeg_in_a57 or jpeg_in_a56 or jpeg_in_a55 or jpeg_in_a54 or jpeg_in_a53 or 
	jpeg_in_a52 or jpeg_in_a51 or jpeg_in_a50 or jpeg_in_a49 or jpeg_in_a48 or 
	jpeg_in_a47 or jpeg_in_a46 or jpeg_in_a45 or jpeg_in_a44 or jpeg_in_a43 or 
	jpeg_in_a42 or jpeg_in_a41 or jpeg_in_a40 or jpeg_in_a39 or jpeg_in_a38 or 
	jpeg_in_a37 or jpeg_in_a36 or jpeg_in_a35 or jpeg_in_a34 or jpeg_in_a33 or 
	jpeg_in_a32 or jpeg_in_a31 or jpeg_in_a30 or jpeg_in_a29 or jpeg_in_a28 or 
	jpeg_in_a27 or jpeg_in_a26 or jpeg_in_a25 or jpeg_in_a24 or jpeg_in_a23 or 
	jpeg_in_a22 or jpeg_in_a21 or jpeg_in_a20 or jpeg_in_a19 or jpeg_in_a18 or 
	jpeg_in_a17 or jpeg_in_a16 or jpeg_in_a15 or jpeg_in_a14 or jpeg_in_a13 or 
	jpeg_in_a12 or jpeg_in_a11 or jpeg_in_a10 or jpeg_in_a09 or jpeg_in_a08 or 
	jpeg_in_a07 or jpeg_in_a06 or jpeg_in_a05 or jpeg_in_a04 or jpeg_in_a03 or 
	jpeg_in_a02 or jpeg_in_a01 or jpeg_in_a00 or RG_y_02 or add3u1ot )	// line#=../rle.cpp:45
	case ( { add3u1ot , RG_y_02 [2:0] } )
	7'h00 :
		quantized_block_wd01 = jpeg_in_a00 ;	// line#=../rle.cpp:45
	7'h01 :
		quantized_block_wd01 = jpeg_in_a01 ;	// line#=../rle.cpp:45
	7'h02 :
		quantized_block_wd01 = jpeg_in_a02 ;	// line#=../rle.cpp:45
	7'h03 :
		quantized_block_wd01 = jpeg_in_a03 ;	// line#=../rle.cpp:45
	7'h04 :
		quantized_block_wd01 = jpeg_in_a04 ;	// line#=../rle.cpp:45
	7'h05 :
		quantized_block_wd01 = jpeg_in_a05 ;	// line#=../rle.cpp:45
	7'h06 :
		quantized_block_wd01 = jpeg_in_a06 ;	// line#=../rle.cpp:45
	7'h07 :
		quantized_block_wd01 = jpeg_in_a07 ;	// line#=../rle.cpp:45
	7'h08 :
		quantized_block_wd01 = jpeg_in_a08 ;	// line#=../rle.cpp:45
	7'h09 :
		quantized_block_wd01 = jpeg_in_a09 ;	// line#=../rle.cpp:45
	7'h0a :
		quantized_block_wd01 = jpeg_in_a10 ;	// line#=../rle.cpp:45
	7'h0b :
		quantized_block_wd01 = jpeg_in_a11 ;	// line#=../rle.cpp:45
	7'h0c :
		quantized_block_wd01 = jpeg_in_a12 ;	// line#=../rle.cpp:45
	7'h0d :
		quantized_block_wd01 = jpeg_in_a13 ;	// line#=../rle.cpp:45
	7'h0e :
		quantized_block_wd01 = jpeg_in_a14 ;	// line#=../rle.cpp:45
	7'h0f :
		quantized_block_wd01 = jpeg_in_a15 ;	// line#=../rle.cpp:45
	7'h10 :
		quantized_block_wd01 = jpeg_in_a16 ;	// line#=../rle.cpp:45
	7'h11 :
		quantized_block_wd01 = jpeg_in_a17 ;	// line#=../rle.cpp:45
	7'h12 :
		quantized_block_wd01 = jpeg_in_a18 ;	// line#=../rle.cpp:45
	7'h13 :
		quantized_block_wd01 = jpeg_in_a19 ;	// line#=../rle.cpp:45
	7'h14 :
		quantized_block_wd01 = jpeg_in_a20 ;	// line#=../rle.cpp:45
	7'h15 :
		quantized_block_wd01 = jpeg_in_a21 ;	// line#=../rle.cpp:45
	7'h16 :
		quantized_block_wd01 = jpeg_in_a22 ;	// line#=../rle.cpp:45
	7'h17 :
		quantized_block_wd01 = jpeg_in_a23 ;	// line#=../rle.cpp:45
	7'h18 :
		quantized_block_wd01 = jpeg_in_a24 ;	// line#=../rle.cpp:45
	7'h19 :
		quantized_block_wd01 = jpeg_in_a25 ;	// line#=../rle.cpp:45
	7'h1a :
		quantized_block_wd01 = jpeg_in_a26 ;	// line#=../rle.cpp:45
	7'h1b :
		quantized_block_wd01 = jpeg_in_a27 ;	// line#=../rle.cpp:45
	7'h1c :
		quantized_block_wd01 = jpeg_in_a28 ;	// line#=../rle.cpp:45
	7'h1d :
		quantized_block_wd01 = jpeg_in_a29 ;	// line#=../rle.cpp:45
	7'h1e :
		quantized_block_wd01 = jpeg_in_a30 ;	// line#=../rle.cpp:45
	7'h1f :
		quantized_block_wd01 = jpeg_in_a31 ;	// line#=../rle.cpp:45
	7'h20 :
		quantized_block_wd01 = jpeg_in_a32 ;	// line#=../rle.cpp:45
	7'h21 :
		quantized_block_wd01 = jpeg_in_a33 ;	// line#=../rle.cpp:45
	7'h22 :
		quantized_block_wd01 = jpeg_in_a34 ;	// line#=../rle.cpp:45
	7'h23 :
		quantized_block_wd01 = jpeg_in_a35 ;	// line#=../rle.cpp:45
	7'h24 :
		quantized_block_wd01 = jpeg_in_a36 ;	// line#=../rle.cpp:45
	7'h25 :
		quantized_block_wd01 = jpeg_in_a37 ;	// line#=../rle.cpp:45
	7'h26 :
		quantized_block_wd01 = jpeg_in_a38 ;	// line#=../rle.cpp:45
	7'h27 :
		quantized_block_wd01 = jpeg_in_a39 ;	// line#=../rle.cpp:45
	7'h28 :
		quantized_block_wd01 = jpeg_in_a40 ;	// line#=../rle.cpp:45
	7'h29 :
		quantized_block_wd01 = jpeg_in_a41 ;	// line#=../rle.cpp:45
	7'h2a :
		quantized_block_wd01 = jpeg_in_a42 ;	// line#=../rle.cpp:45
	7'h2b :
		quantized_block_wd01 = jpeg_in_a43 ;	// line#=../rle.cpp:45
	7'h2c :
		quantized_block_wd01 = jpeg_in_a44 ;	// line#=../rle.cpp:45
	7'h2d :
		quantized_block_wd01 = jpeg_in_a45 ;	// line#=../rle.cpp:45
	7'h2e :
		quantized_block_wd01 = jpeg_in_a46 ;	// line#=../rle.cpp:45
	7'h2f :
		quantized_block_wd01 = jpeg_in_a47 ;	// line#=../rle.cpp:45
	7'h30 :
		quantized_block_wd01 = jpeg_in_a48 ;	// line#=../rle.cpp:45
	7'h31 :
		quantized_block_wd01 = jpeg_in_a49 ;	// line#=../rle.cpp:45
	7'h32 :
		quantized_block_wd01 = jpeg_in_a50 ;	// line#=../rle.cpp:45
	7'h33 :
		quantized_block_wd01 = jpeg_in_a51 ;	// line#=../rle.cpp:45
	7'h34 :
		quantized_block_wd01 = jpeg_in_a52 ;	// line#=../rle.cpp:45
	7'h35 :
		quantized_block_wd01 = jpeg_in_a53 ;	// line#=../rle.cpp:45
	7'h36 :
		quantized_block_wd01 = jpeg_in_a54 ;	// line#=../rle.cpp:45
	7'h37 :
		quantized_block_wd01 = jpeg_in_a55 ;	// line#=../rle.cpp:45
	7'h38 :
		quantized_block_wd01 = jpeg_in_a56 ;	// line#=../rle.cpp:45
	7'h39 :
		quantized_block_wd01 = jpeg_in_a57 ;	// line#=../rle.cpp:45
	7'h3a :
		quantized_block_wd01 = jpeg_in_a58 ;	// line#=../rle.cpp:45
	7'h3b :
		quantized_block_wd01 = jpeg_in_a59 ;	// line#=../rle.cpp:45
	7'h3c :
		quantized_block_wd01 = jpeg_in_a60 ;	// line#=../rle.cpp:45
	7'h3d :
		quantized_block_wd01 = jpeg_in_a61 ;	// line#=../rle.cpp:45
	7'h3e :
		quantized_block_wd01 = jpeg_in_a62 ;	// line#=../rle.cpp:45
	7'h3f :
		quantized_block_wd01 = jpeg_in_a63 ;	// line#=../rle.cpp:45
	7'h40 :
		quantized_block_wd01 = jpeg_in_a64 ;	// line#=../rle.cpp:45
	7'h41 :
		quantized_block_wd01 = jpeg_in_a65 ;	// line#=../rle.cpp:45
	7'h42 :
		quantized_block_wd01 = jpeg_in_a66 ;	// line#=../rle.cpp:45
	7'h43 :
		quantized_block_wd01 = jpeg_in_a67 ;	// line#=../rle.cpp:45
	7'h44 :
		quantized_block_wd01 = jpeg_in_a68 ;	// line#=../rle.cpp:45
	7'h45 :
		quantized_block_wd01 = jpeg_in_a69 ;	// line#=../rle.cpp:45
	7'h46 :
		quantized_block_wd01 = jpeg_in_a70 ;	// line#=../rle.cpp:45
	7'h47 :
		quantized_block_wd01 = jpeg_in_a71 ;	// line#=../rle.cpp:45
	7'h48 :
		quantized_block_wd01 = jpeg_in_a72 ;	// line#=../rle.cpp:45
	7'h49 :
		quantized_block_wd01 = jpeg_in_a73 ;	// line#=../rle.cpp:45
	7'h4a :
		quantized_block_wd01 = jpeg_in_a74 ;	// line#=../rle.cpp:45
	7'h4b :
		quantized_block_wd01 = jpeg_in_a75 ;	// line#=../rle.cpp:45
	7'h4c :
		quantized_block_wd01 = jpeg_in_a76 ;	// line#=../rle.cpp:45
	7'h4d :
		quantized_block_wd01 = jpeg_in_a77 ;	// line#=../rle.cpp:45
	7'h4e :
		quantized_block_wd01 = jpeg_in_a78 ;	// line#=../rle.cpp:45
	7'h4f :
		quantized_block_wd01 = jpeg_in_a79 ;	// line#=../rle.cpp:45
	7'h50 :
		quantized_block_wd01 = jpeg_in_a80 ;	// line#=../rle.cpp:45
	7'h51 :
		quantized_block_wd01 = jpeg_in_a81 ;	// line#=../rle.cpp:45
	7'h52 :
		quantized_block_wd01 = jpeg_in_a82 ;	// line#=../rle.cpp:45
	7'h53 :
		quantized_block_wd01 = jpeg_in_a83 ;	// line#=../rle.cpp:45
	7'h54 :
		quantized_block_wd01 = jpeg_in_a84 ;	// line#=../rle.cpp:45
	7'h55 :
		quantized_block_wd01 = jpeg_in_a85 ;	// line#=../rle.cpp:45
	7'h56 :
		quantized_block_wd01 = jpeg_in_a86 ;	// line#=../rle.cpp:45
	7'h57 :
		quantized_block_wd01 = jpeg_in_a87 ;	// line#=../rle.cpp:45
	7'h58 :
		quantized_block_wd01 = jpeg_in_a88 ;	// line#=../rle.cpp:45
	7'h59 :
		quantized_block_wd01 = jpeg_in_a89 ;	// line#=../rle.cpp:45
	7'h5a :
		quantized_block_wd01 = jpeg_in_a90 ;	// line#=../rle.cpp:45
	7'h5b :
		quantized_block_wd01 = jpeg_in_a91 ;	// line#=../rle.cpp:45
	7'h5c :
		quantized_block_wd01 = jpeg_in_a92 ;	// line#=../rle.cpp:45
	7'h5d :
		quantized_block_wd01 = jpeg_in_a93 ;	// line#=../rle.cpp:45
	7'h5e :
		quantized_block_wd01 = jpeg_in_a94 ;	// line#=../rle.cpp:45
	7'h5f :
		quantized_block_wd01 = jpeg_in_a95 ;	// line#=../rle.cpp:45
	7'h60 :
		quantized_block_wd01 = jpeg_in_a96 ;	// line#=../rle.cpp:45
	7'h61 :
		quantized_block_wd01 = jpeg_in_a97 ;	// line#=../rle.cpp:45
	7'h62 :
		quantized_block_wd01 = jpeg_in_a98 ;	// line#=../rle.cpp:45
	7'h63 :
		quantized_block_wd01 = jpeg_in_a99 ;	// line#=../rle.cpp:45
	7'h64 :
		quantized_block_wd01 = jpeg_in_a100 ;	// line#=../rle.cpp:45
	7'h65 :
		quantized_block_wd01 = jpeg_in_a101 ;	// line#=../rle.cpp:45
	7'h66 :
		quantized_block_wd01 = jpeg_in_a102 ;	// line#=../rle.cpp:45
	7'h67 :
		quantized_block_wd01 = jpeg_in_a103 ;	// line#=../rle.cpp:45
	7'h68 :
		quantized_block_wd01 = jpeg_in_a104 ;	// line#=../rle.cpp:45
	7'h69 :
		quantized_block_wd01 = jpeg_in_a105 ;	// line#=../rle.cpp:45
	7'h6a :
		quantized_block_wd01 = jpeg_in_a106 ;	// line#=../rle.cpp:45
	7'h6b :
		quantized_block_wd01 = jpeg_in_a107 ;	// line#=../rle.cpp:45
	7'h6c :
		quantized_block_wd01 = jpeg_in_a108 ;	// line#=../rle.cpp:45
	7'h6d :
		quantized_block_wd01 = jpeg_in_a109 ;	// line#=../rle.cpp:45
	7'h6e :
		quantized_block_wd01 = jpeg_in_a110 ;	// line#=../rle.cpp:45
	7'h6f :
		quantized_block_wd01 = jpeg_in_a111 ;	// line#=../rle.cpp:45
	7'h70 :
		quantized_block_wd01 = jpeg_in_a112 ;	// line#=../rle.cpp:45
	7'h71 :
		quantized_block_wd01 = jpeg_in_a113 ;	// line#=../rle.cpp:45
	7'h72 :
		quantized_block_wd01 = jpeg_in_a114 ;	// line#=../rle.cpp:45
	7'h73 :
		quantized_block_wd01 = jpeg_in_a115 ;	// line#=../rle.cpp:45
	7'h74 :
		quantized_block_wd01 = jpeg_in_a116 ;	// line#=../rle.cpp:45
	7'h75 :
		quantized_block_wd01 = jpeg_in_a117 ;	// line#=../rle.cpp:45
	7'h76 :
		quantized_block_wd01 = jpeg_in_a118 ;	// line#=../rle.cpp:45
	7'h77 :
		quantized_block_wd01 = jpeg_in_a119 ;	// line#=../rle.cpp:45
	7'h78 :
		quantized_block_wd01 = jpeg_in_a120 ;	// line#=../rle.cpp:45
	7'h79 :
		quantized_block_wd01 = jpeg_in_a121 ;	// line#=../rle.cpp:45
	7'h7a :
		quantized_block_wd01 = jpeg_in_a122 ;	// line#=../rle.cpp:45
	7'h7b :
		quantized_block_wd01 = jpeg_in_a123 ;	// line#=../rle.cpp:45
	7'h7c :
		quantized_block_wd01 = jpeg_in_a124 ;	// line#=../rle.cpp:45
	7'h7d :
		quantized_block_wd01 = jpeg_in_a125 ;	// line#=../rle.cpp:45
	7'h7e :
		quantized_block_wd01 = jpeg_in_a126 ;	// line#=../rle.cpp:45
	7'h7f :
		quantized_block_wd01 = jpeg_in_a127 ;	// line#=../rle.cpp:45
	default :
		quantized_block_wd01 = 9'hx ;
	endcase
assign	C_01 = ~|{ ~incr4s1ot [3] , incr4s1ot [2:0] } ;	// line#=../rle.cpp:34,35
assign	U_04 = ( ST1_02d & ( ~JF_01 ) ) ;
assign	U_05 = ( ST1_03d & FL01_01_01a ) ;
assign	U_06 = ( U_05 & ( ~RG_j_x_02 [3] ) ) ;	// line#=../rle.cpp:42
assign	U_10 = ( ST1_03d & FL01_02_01a ) ;
assign	U_15 = ( ST1_03d & FL01_01_streg ) ;
assign	U_17 = ( U_15 & ( ~FL01_02_01_stall ) ) ;
assign	U_19 = ( U_17 & ( ~FJ_03_05 ) ) ;
assign	U_20 = ( ST1_03d & ( ~FL01_02_streg ) ) ;
assign	U_21 = ( ST1_03d & FL01_02_streg ) ;
assign	U_24 = ( U_21 & FJ_04_04 ) ;
assign	U_25 = ( U_21 & ( ~FJ_04_04 ) ) ;
assign	U_28 = ( ST1_03d & FL01_01_break ) ;
assign	U_34 = ( ST1_05d & lop8u_11ot ) ;	// line#=../rle.cpp:109,110
assign	U_35 = ( ST1_05d & ( ~lop8u_11ot ) ) ;	// line#=../rle.cpp:109,110
assign	C_04 = ( ( ~|RG_i ) & M_442 ) ;	// line#=../rle.cpp:112,113
assign	U_36 = ( U_34 & C_04 ) ;	// line#=../rle.cpp:112,113
assign	U_37 = ( U_34 & ( ~C_04 ) ) ;	// line#=../rle.cpp:112,113
assign	U_38 = ( U_37 & CT_06 ) ;	// line#=../rle.cpp:117,118
assign	U_39 = ( U_37 & ( ~CT_06 ) ) ;	// line#=../rle.cpp:117,118
assign	U_40 = ( U_39 & ( ~FF_d_05 ) ) ;	// line#=../rle.cpp:122,123
assign	U_41 = ( U_39 & FF_d_05 ) ;	// line#=../rle.cpp:122,123
assign	U_44 = ( ST1_06d & ( ~RG_k_05 [6] ) ) ;	// line#=../rle.cpp:140,141
assign	M_442 = ~|{ ( RG_j_k [31] & RG_j_k [0] ) , RG_j_k [0] } ;	// line#=../rle.cpp:112,113,143,144
assign	C_06 = ( ( ~|{ RG_i [31:3] , ~RG_i [2:0] } ) & M_442 ) ;	// line#=../rle.cpp:143,144
assign	U_46 = ( U_44 & C_06 ) ;	// line#=../rle.cpp:143,144
assign	U_47 = ( U_44 & ( ~C_06 ) ) ;	// line#=../rle.cpp:143,144
assign	U_48 = ( U_47 & CT_11 ) ;	// line#=../rle.cpp:148,149
assign	U_49 = ( U_47 & ( ~CT_11 ) ) ;	// line#=../rle.cpp:148,149
assign	U_50 = ( U_49 & ( ~FF_d_05 ) ) ;	// line#=../rle.cpp:153,154
assign	U_51 = ( U_49 & FF_d_05 ) ;	// line#=../rle.cpp:153,154
assign	U_54 = ( ST1_08d & FL02_01_01a ) ;
assign	C_08 = ( RG_i_06 [31] | ( ~|RG_i_06 [30:6] ) ) ;	// line#=../rle.cpp:57,58
assign	U_55 = ( U_54 & C_08 ) ;	// line#=../rle.cpp:57,58
assign	U_58 = ( ST1_08d & FL02_02_01a ) ;
assign	U_59 = ( U_58 & CT_14 ) ;	// line#=../rle.cpp:61,62
assign	U_61 = ( ST1_08d & FL02_03_01a ) ;
assign	U_67 = ( ST1_08d & FL02_04_01a ) ;
assign	U_68 = ( ST1_08d & FL02_05_01a ) ;
assign	U_69 = ( U_68 & CT_16 ) ;	// line#=../rle.cpp:66,67
assign	U_70 = ( U_68 & ( ~CT_16 ) ) ;	// line#=../rle.cpp:66,67
assign	U_72 = ( ST1_08d & FL02_06_01a ) ;
assign	U_73 = ( U_72 & FF_d_05 ) ;	// line#=../rle.cpp:66,67
assign	U_74 = ( U_72 & ( ~FF_d_05 ) ) ;	// line#=../rle.cpp:66,67
assign	U_75 = ( ST1_08d & ( ~|( FL02_01_streg ^ 2'h2 ) ) ) ;
assign	U_77 = ( ST1_08d & M_435 ) ;
assign	U_79 = ( U_75 & ( ~FL02_02_Lrdy ) ) ;
assign	C_12 = ( flag_r1 & flag_r2 ) ;
assign	U_82 = ( U_77 & C_12 ) ;
assign	U_85 = ( U_82 & ( ~FJ_09_15 ) ) ;
assign	U_87 = ( U_85 & ( ~FL02_02_Lrdy ) ) ;
assign	U_91 = ( ST1_08d & ( ~|( FL02_02_streg ^ 2'h1 ) ) ) ;
assign	U_92 = ( ST1_08d & ( ~|( FL02_02_streg ^ 2'h2 ) ) ) ;
assign	U_93 = ( ST1_08d & ( ~|( FL02_02_streg ^ 2'h3 ) ) ) ;
assign	U_94 = ( ( ST1_08d & ( ~|FL02_02_streg ) ) & flag_r3 ) ;
assign	U_95 = ( U_94 & FL02_01_ndat ) ;
assign	U_96 = ( U_94 & ( ~FL02_01_ndat ) ) ;
assign	U_99 = ( U_92 & FL02_02_Leos_all ) ;
assign	U_102 = ( U_99 & ( ~FL02_04_rdy ) ) ;
assign	U_103 = ( U_93 & ( ~U_112 ) ) ;
assign	U_105 = ( U_103 & FA02_02_gnt ) ;
assign	U_107 = ( ST1_08d & ( ~FL02_03_streg ) ) ;
assign	U_108 = ( ST1_08d & FL02_03_streg ) ;
assign	U_111 = ( U_108 & FA02_03_gnt ) ;
assign	U_112 = ( U_108 & ( ~FA02_03_gnt ) ) ;
assign	U_114 = ( U_111 & ( ~FJ_11_12 ) ) ;
assign	U_117 = ( ST1_08d & ( ~FL02_04_streg ) ) ;
assign	U_118 = ( ST1_08d & FL02_04_streg ) ;
assign	U_121 = ( U_118 & ( ~FL02_05_ngo ) ) ;
assign	U_123 = ( U_121 & FL02_02_Lndat ) ;
assign	U_125 = ( ST1_08d & ( ~FL02_05_streg ) ) ;
assign	U_126 = ( ST1_08d & FL02_05_streg ) ;
assign	U_129 = ( U_126 & ( ~U_140 ) ) ;
assign	U_130 = ( U_126 & U_140 ) ;
assign	U_131 = ( U_129 & U_129 ) ;
assign	U_132 = ( U_129 & ( ~U_129 ) ) ;
assign	U_135 = ( ST1_08d & ( ~FL02_06_streg ) ) ;
assign	U_136 = ( ST1_08d & FL02_06_streg ) ;
assign	U_139 = ( U_136 & U_136 ) ;
assign	U_140 = ( U_136 & ( ~U_136 ) ) ;
assign	U_143 = ( ST1_08d & FL02_01_break ) ;
assign	U_147 = ( ST1_08d & FL02_03_break ) ;
assign	U_159 = ( ST1_11d & ( ~FF_d_05 ) ) ;	// line#=../rle.cpp:77,78
assign	U_164 = ( ST1_14d & ( ~CT_20 ) ) ;	// line#=../rle.cpp:83,84
assign	U_165 = ( ST1_14d & RG_15_02 ) ;	// line#=../rle.cpp:61,62,83,84
assign	RG_previous_dc_en = ST1_07d ;
always @ ( posedge clk )	// line#=../rle.cpp:52,53
	if ( !rst )
		RG_previous_dc <= 9'h000 ;
	else if ( RG_previous_dc_en )
		RG_previous_dc <= zz_RD1 ;
always @ ( incr4s1ot or U_10 or FL01_02_01_stall or U_06 )	// line#=../rle.cpp:44
	begin
	RG_y_02_t_c1 = ( U_06 & ( ~FL01_02_01_stall ) ) ;	// line#=../rle.cpp:44
	RG_y_02_t_c2 = ( U_10 & ( ~incr4s1ot [3] ) ) ;	// line#=../rle.cpp:44
	RG_y_02_t = ( { 4{ RG_y_02_t_c2 } } & incr4s1ot )	// line#=../rle.cpp:44
		 ;	// line#=../rle.cpp:44
	end
assign	RG_y_02_en = ( RG_y_02_t_c1 | RG_y_02_t_c2 ) ;	// line#=../rle.cpp:44
always @ ( posedge clk )	// line#=../rle.cpp:44
	if ( RG_y_02_en )
		RG_y_02 <= RG_y_02_t ;	// line#=../rle.cpp:44
always @ ( incr3u1ot or U_06 or incr4s1ot or FF_j or ST1_14d or C_01 or ST1_02d or 
	ST1_01d )	// line#=../rle.cpp:35
	begin
	RG_j_x_02_t_c1 = ( ( ST1_02d & C_01 ) | ST1_14d ) ;	// line#=../rle.cpp:42
	RG_j_x_02_t_c2 = ( ST1_02d & ( ~C_01 ) ) ;	// line#=../rle.cpp:34
	RG_j_x_02_t = ( ( { 4{ ST1_01d } } & 4'hf /*-4'h1*/ )			// line#=../rle.cpp:34
		| ( { 4{ RG_j_x_02_t_c1 } } & { 3'h0 , ( ST1_14d & FF_j ) } )	// line#=../rle.cpp:42
		| ( { 4{ RG_j_x_02_t_c2 } } & incr4s1ot )			// line#=../rle.cpp:34
		| ( { 4{ U_06 } } & incr3u1ot )					// line#=../rle.cpp:42
		) ;
	end
assign	RG_j_x_02_en = ( ST1_01d | RG_j_x_02_t_c1 | RG_j_x_02_t_c2 | U_06 ) ;	// line#=../rle.cpp:35
always @ ( posedge clk )	// line#=../rle.cpp:35
	if ( ( RG_j_x_02_en & ( !FL01_02_01_stall ) ) )
		RG_j_x_02 <= RG_j_x_02_t ;	// line#=../rle.cpp:34,35,42
assign	RG_03_02_en = U_06 ;
always @ ( posedge clk )	// line#=../rle.cpp:42
	if ( ( RG_03_02_en & ( !FL01_02_01_stall ) ) )
		RG_03_02 <= RG_j_x_02 [2:0] ;
always @ ( RG_i_05 or U_73 or incr32s3ot or U_74 or U_72 or ST1_02d )
	begin
	RG_i_06_t_c1 = ( U_72 & U_74 ) ;	// line#=../rle.cpp:74
	RG_i_06_t_c2 = ( U_72 & U_73 ) ;
	RG_i_06_t = ( ( { 32{ ST1_02d } } & 32'h00000001 )	// line#=../rle.cpp:37
		| ( { 32{ RG_i_06_t_c1 } } & incr32s3ot )	// line#=../rle.cpp:74
		| ( { 32{ RG_i_06_t_c2 } } & RG_i_05 ) ) ;
	end
assign	RG_i_06_en = ( ST1_02d | RG_i_06_t_c1 | RG_i_06_t_c2 ) ;
always @ ( posedge clk )
	if ( RG_i_06_en )
		RG_i_06 <= RG_i_06_t ;	// line#=../rle.cpp:37,74
always @ ( sub8u1ot or ST1_15d or incr8u1ot or ST1_12d or U_159 or incr8u2ot or 
	U_68 or ST1_02d )
	begin
	RG_len_05_t_c1 = ( U_159 | ST1_12d ) ;	// line#=../rle.cpp:79,80
	RG_len_05_t = ( ( { 8{ ST1_02d } } & 8'h01 )		// line#=../rle.cpp:39
		| ( { 8{ U_68 } } & incr8u2ot )			// line#=../rle.cpp:66,67,69,74
		| ( { 8{ RG_len_05_t_c1 } } & incr8u1ot )	// line#=../rle.cpp:79,80
		| ( { 8{ ST1_15d } } & sub8u1ot )		// line#=../rle.cpp:86
		) ;
	end
assign	RG_len_05_en = ( ST1_02d | U_68 | RG_len_05_t_c1 | ST1_15d ) ;
always @ ( posedge clk )
	if ( RG_len_05_en )
		RG_len_05 <= RG_len_05_t ;	// line#=../rle.cpp:39,66,67,69,74,79,80
						// ,86
assign	FF_j_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:36
	if ( FF_j_en )
		FF_j <= 1'h0 ;
assign	RG_i_03_en = U_61 ;
always @ ( posedge clk )
	if ( RG_i_03_en )
		RG_i_03 <= RG_i_02 ;
assign	RG_k_03_en = U_61 ;
always @ ( posedge clk )
	if ( RG_k_03_en )
		RG_k_03 <= RG_k_02 [8:0] ;
always @ ( U_35 )
	TR_02 = ( { 3{ U_35 } } & 3'h7 )	// line#=../rle.cpp:134
		 ;	// line#=../rle.cpp:105
always @ ( RG_i_06 or U_55 or decr32s1ot or U_50 or U_40 or incr32s2ot or U_58 or 
	U_51 or U_48 or U_41 or U_38 or TR_02 or M_447 )
	begin
	RG_i_t_c1 = ( ( ( ( U_38 | U_41 ) | U_48 ) | U_51 ) | U_58 ) ;	// line#=../rle.cpp:61,62,63,119,129,150
									// ,160
	RG_i_t_c2 = ( U_40 | U_50 ) ;	// line#=../rle.cpp:124,155
	RG_i_t = ( ( { 32{ M_447 } } & { 29'h00000000 , TR_02 } )	// line#=../rle.cpp:105,134
		| ( { 32{ RG_i_t_c1 } } & incr32s2ot )			// line#=../rle.cpp:61,62,63,119,129,150
									// ,160
		| ( { 32{ RG_i_t_c2 } } & decr32s1ot )			// line#=../rle.cpp:124,155
		| ( { 32{ U_55 } } & RG_i_06 ) ) ;
	end
assign	RG_i_en = ( M_447 | RG_i_t_c1 | RG_i_t_c2 | U_55 ) ;
always @ ( posedge clk )
	if ( RG_i_en )
		RG_i <= RG_i_t ;	// line#=../rle.cpp:61,62,63,105,119,124
					// ,129,134,150,155,160
always @ ( decr32s2ot or U_51 or U_41 or incr32s1ot or U_58 or U_50 or U_46 or U_40 or 
	U_36 or U_35 or U_55 or ST1_04d )
	begin
	RG_j_k_t_c1 = ( ( ST1_04d | U_55 ) | U_35 ) ;	// line#=../rle.cpp:59,105,135
	RG_j_k_t_c2 = ( ( ( ( U_36 | U_40 ) | U_46 ) | U_50 ) | U_58 ) ;	// line#=../rle.cpp:64,114,125,145,156
	RG_j_k_t_c3 = ( U_41 | U_51 ) ;	// line#=../rle.cpp:130,161
	RG_j_k_t = ( ( { 32{ RG_j_k_t_c1 } } & { 31'h00000000 , U_35 } )	// line#=../rle.cpp:59,105,135
		| ( { 32{ RG_j_k_t_c2 } } & incr32s1ot )			// line#=../rle.cpp:64,114,125,145,156
		| ( { 32{ RG_j_k_t_c3 } } & decr32s2ot )			// line#=../rle.cpp:130,161
		) ;
	end
assign	RG_j_k_en = ( RG_j_k_t_c1 | RG_j_k_t_c2 | RG_j_k_t_c3 ) ;
always @ ( posedge clk )
	if ( RG_j_k_en )
		RG_j_k <= RG_j_k_t ;	// line#=../rle.cpp:59,64,105,114,125,130
					// ,135,145,156,161
always @ ( incr8u_61ot or ST1_05d )
	RG_k_t = ( { 6{ ST1_05d } } & incr8u_61ot )	// line#=../rle.cpp:111
		 ;	// line#=../rle.cpp:105
always @ ( posedge clk )
	RG_k <= RG_k_t ;	// line#=../rle.cpp:105,111
assign	M_447 = ( ST1_04d | U_35 ) ;
always @ ( CT_17 or ST1_10d or CT_16 or U_68 or U_48 or U_36 or ST1_09d or U_46 or 
	U_38 or M_447 )
	begin
	FF_d_05_t_c1 = ( ( ( M_447 | U_38 ) | U_46 ) | ST1_09d ) ;	// line#=../rle.cpp:77,78,105,120,136,146
	FF_d_05_t_c2 = ( U_36 | U_48 ) ;	// line#=../rle.cpp:115,151
	FF_d_05_t = ( ( { 1{ FF_d_05_t_c2 } } & 1'h1 )	// line#=../rle.cpp:115,151
		| ( { 1{ U_68 } } & CT_16 )		// line#=../rle.cpp:66,67
		| ( { 1{ ST1_10d } } & CT_17 )		// line#=../rle.cpp:77,78
		) ;	// line#=../rle.cpp:77,78,105,120,136,146
	end
assign	FF_d_05_en = ( FF_d_05_t_c1 | FF_d_05_t_c2 | U_68 | ST1_10d ) ;
always @ ( posedge clk )
	if ( FF_d_05_en )
		FF_d_05 <= FF_d_05_t ;	// line#=../rle.cpp:66,67,77,78,105,115
					// ,120,136,146,151
assign	RG_i_02_en = U_58 ;
always @ ( posedge clk )
	if ( RG_i_02_en )
		RG_i_02 <= RG_i ;
assign	RG_k_02_en = U_58 ;
always @ ( posedge clk )	// line#=../rle.cpp:61,62
	if ( RG_k_02_en )
		RG_k_02 <= RG_j_k ;
always @ ( CT_20 or ST1_14d or rl_rd00 or ST1_13d or FF_d_05 or ST1_11d or CT_17 or 
	ST1_09d or CT_14 or U_58 or RG_k_05 or ST1_06d )
	RG_15_02_t = ( ( { 1{ ST1_06d } } & ( ~RG_k_05 [6] ) )				// line#=../rle.cpp:140,141
		| ( { 1{ U_58 } } & CT_14 )						// line#=../rle.cpp:61,62
		| ( { 1{ ST1_09d } } & CT_17 )						// line#=../rle.cpp:77,78
		| ( { 1{ ST1_11d } } & ( ~FF_d_05 ) )					// line#=../rle.cpp:77,78
		| ( { 1{ ST1_13d } } & ( ~|{ rl_rd00 [8:4] , ~rl_rd00 [3:0] } ) )	// line#=../rle.cpp:83,84
		| ( { 1{ ST1_14d } } & CT_20 )						// line#=../rle.cpp:83,84
		) ;
assign	RG_15_02_en = ( ST1_06d | U_58 | ST1_09d | ST1_11d | ST1_13d | ST1_14d ) ;
always @ ( posedge clk )
	if ( RG_15_02_en )
		RG_15_02 <= RG_15_02_t ;	// line#=../rle.cpp:61,62,77,78,83,84,140
						// ,141
always @ ( sub8u1ot or ST1_13d or incr8u1ot or M_454 or incr8u_71ot or ST1_06d or 
	RG_k or ST1_05d )
	RG_k_05_t = ( ( { 7{ ST1_05d } } & { 1'h0 , RG_k } )
		| ( { 7{ ST1_06d } } & incr8u_71ot )	// line#=../rle.cpp:142
		| ( { 7{ M_454 } } & incr8u1ot [6:0] )	// line#=../rle.cpp:68,69,73,74
		| ( { 7{ ST1_13d } } & sub8u1ot [6:0] )	// line#=../rle.cpp:83,84
		) ;
assign	RG_k_05_en = ( ST1_05d | ST1_06d | M_454 | ST1_13d ) ;
always @ ( posedge clk )
	if ( RG_k_05_en )
		RG_k_05 <= RG_k_05_t ;	// line#=../rle.cpp:68,69,73,74,83,84,142
assign	RG_i_04_en = U_67 ;
always @ ( posedge clk )
	if ( RG_i_04_en )
		RG_i_04 <= RG_i_03 ;
assign	RG_k_04_en = U_67 ;
always @ ( posedge clk )
	if ( RG_k_04_en )
		RG_k_04 <= RG_k_03 ;
assign	RG_i_05_en = U_68 ;
always @ ( posedge clk )
	if ( RG_i_05_en )
		RG_i_05 <= RG_i_04 ;
assign	JF_01 = ~C_01 ;
assign	JF_01_port = JF_01 ;
assign	JF_05 = ~RG_k_05 [6] ;
assign	JF_09 = ~FF_d_05 ;	// line#=../rle.cpp:77,78
assign	JF_10 = ~CT_20 ;	// line#=../rle.cpp:83,84
assign	FL01_01_break = ( FL01_01_streg & FJ_03_05 ) ;
assign	FL01_01_01a = U_15 ;
assign	FL01_02_01a = U_21 ;
assign	FJ_03_05 = ( ( ~FL01_02_01_stall ) & ( U_05 & ( ~( ~RG_j_x_02 [3] ) ) ) ) ;	// line#=../rle.cpp:42
assign	FJ_04_04 = ( U_10 & ( ~incr4s1ot [3] ) ) ;	// line#=../rle.cpp:44
assign	FL01_01_eos = ( M_452 | U_28 ) ;
assign	FL01_02_eos = M_453 ;
assign	M_445 = ( ST1_03d & ( ~FL01_01_break ) ) ;
assign	M_452 = ( ( U_17 & FJ_03_05 ) | ( ST1_03d & ( ~FL01_01_streg ) ) ) ;
always @ ( U_04 or U_19 or FL01_02_01_stall or U_15 or M_452 or M_445 or U_28 )
	begin
	FL01_01_streg_t_c1 = ( U_28 | ( M_445 & M_452 ) ) ;
	FL01_01_streg_t_c2 = ( ( M_445 & ( ( U_15 & FL01_02_01_stall ) | U_19 ) ) | 
		U_04 ) ;
	FL01_01_streg_t = ( { 1{ FL01_01_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_01_streg_en = ( FL01_01_streg_t_c1 | FL01_01_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_01_streg_en )
		FL01_01_streg <= FL01_01_streg_t ;
assign	M_453 = ( ( U_25 & ( ~FL01_01_ndat ) ) | ( U_20 & ( ~FL01_01_ndat ) ) ) ;
always @ ( U_20 or FL01_01_ndat or U_25 or U_24 or M_453 or ST1_03d or U_04 )
	begin
	FL01_02_streg_t_c1 = ( U_04 | ( ST1_03d & M_453 ) ) ;
	FL01_02_streg_t_c2 = ( ST1_03d & ( ( U_24 | ( U_25 & FL01_01_ndat ) ) | ( 
		U_20 & FL01_01_ndat ) ) ) ;
	FL01_02_streg_t = ( { 1{ FL01_02_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL01_02_streg_en = ( FL01_02_streg_t_c1 | FL01_02_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL01_02_streg_en )
		FL01_02_streg <= FL01_02_streg_t ;
assign	FL01_02_01_stall = U_24 ;
assign	FL01_02_01_stall_port = FL01_02_01_stall ;
assign	FL01_01_ndat = U_19 ;
assign	M_435 = ~|( FL02_01_streg ^ 2'h1 ) ;
assign	FL02_01_break = ( M_435 & FJ_09_15 ) ;
assign	FL02_02_break = ( ( U_93 | U_92 ) & FJ_11_12 ) ;
assign	FL02_03_break = ( FL02_03_streg & FJ_11_12 ) ;
always @ ( ST1_07d or U_139 )
	begin
	flag_r1_t_c1 = ( U_139 | ST1_07d ) ;
	flag_r1_t = ( { 1{ flag_r1_t_c1 } } & 1'h1 )
		 ;
	end
assign	flag_r1_en = ( flag_r1_t_c1 | U_85 ) ;
always @ ( posedge clk )
	if ( flag_r1_en )
		flag_r1 <= flag_r1_t ;
always @ ( ST1_07d or U_99 )
	begin
	flag_r2_t_c1 = ( U_99 | ST1_07d ) ;
	flag_r2_t = ( { 1{ flag_r2_t_c1 } } & 1'h1 )
		 ;
	end
assign	flag_r2_en = ( U_85 | flag_r2_t_c1 ) ;
always @ ( posedge clk )
	if ( flag_r2_en )
		flag_r2 <= flag_r2_t ;
always @ ( ST1_07d or U_121 )
	begin
	flag_r3_t_c1 = ( U_121 | ST1_07d ) ;
	flag_r3_t = ( { 1{ flag_r3_t_c1 } } & 1'h1 )
		 ;
	end
assign	flag_r3_en = ( flag_r3_t_c1 | U_95 ) ;
always @ ( posedge clk )
	if ( flag_r3_en )
		flag_r3 <= flag_r3_t ;
assign	FL02_01_01a = U_82 ;
assign	FL02_02_01a = U_105 ;
assign	FL02_03_01a = U_111 ;
assign	FL02_04_01a = U_121 ;
assign	FL02_05_01a = U_131 ;
assign	FL02_06_01a = U_139 ;
assign	FJ_09_15 = ( U_54 & ( ~C_08 ) ) ;	// line#=../rle.cpp:57,58
assign	FJ_11_12 = ( U_61 & ( ~( M_01_t1 & ( RG_k_02 [31] | ( ( ~|RG_k_02 [30:4] ) & ( 
	~&RG_k_02 [3:0] ) ) ) ) ) ) ;	// line#=../rle.cpp:61,62
assign	FL02_02_Leos = U_96 ;
assign	FL02_01_eos = ( M_455 | U_143 ) ;
assign	FL02_02_eos = ( U_96 | U_92 ) ;
assign	FL02_03_eos = ( M_456 | U_147 ) ;
assign	FL02_04_eos = M_457 ;
assign	FL02_05_eos = M_458 ;
assign	FL02_06_eos = M_459 ;
assign	M_444 = ( ( M_449 & ( ( ( U_77 & ( ~C_12 ) ) | ( U_85 & FL02_02_Lrdy ) ) | 
	( U_75 & FL02_02_Lrdy ) ) ) | ST1_07d ) ;
assign	M_449 = ( ST1_08d & ( ~FL02_01_break ) ) ;
assign	M_455 = ( ( ( ( U_82 & FJ_09_15 ) | ( U_87 & FL02_02_Lrdy ) ) | ( U_79 & 
	FL02_02_Lrdy ) ) | ( ST1_08d & ( ~|FL02_01_streg ) ) ) ;
always @ ( U_79 or FL02_02_Lrdy or U_87 or M_444 or M_455 or M_449 or U_143 )
	begin
	FL02_01_streg_t_c1 = ( ( U_143 | ( M_449 & M_455 ) ) | M_444 ) ;
	FL02_01_streg_t_c2 = ( M_449 & ( ( U_87 & ( ~FL02_02_Lrdy ) ) | ( U_79 & ( 
		~FL02_02_Lrdy ) ) ) ) ;
	FL02_01_streg_t = ( ( { 2{ FL02_01_streg_t_c1 } } & { 1'h0 , M_444 } )
		| ( { 2{ FL02_01_streg_t_c2 } } & 2'h2 ) ) ;
	end
assign	FL02_01_streg_en = ( FL02_01_streg_t_c1 | FL02_01_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL02_01_streg_en )
		FL02_01_streg <= FL02_01_streg_t ;
assign	M_443 = ( ST1_08d & FL02_02_break ) ;
always @ ( FL02_02_Leos_all or U_92 or U_102 or FL02_04_rdy or U_91 or U_95 or U_93 )
	begin
	FL02_02_streg_t1_c1 = ( U_93 | U_95 ) ;
	FL02_02_streg_t1_c2 = ( ( U_91 & ( ~FL02_04_rdy ) ) | U_102 ) ;
	FL02_02_streg_t1_c3 = ( U_92 & ( ~FL02_02_Leos_all ) ) ;
	FL02_02_streg_t1 = ( ( { 2{ FL02_02_streg_t1_c1 } } & 2'h3 )
		| ( { 2{ FL02_02_streg_t1_c2 } } & 2'h1 )
		| ( { 2{ FL02_02_streg_t1_c3 } } & 2'h2 ) ) ;
	end
always @ ( FL02_02_streg_t1 or FL02_02_break or ST1_08d or ST1_07d or M_443 )
	begin
	FL02_02_streg_t_c1 = ( M_443 | ST1_07d ) ;
	FL02_02_streg_t_c2 = ( ST1_08d & ( ~FL02_02_break ) ) ;
	FL02_02_streg_t = ( ( { 2{ FL02_02_streg_t_c1 } } & { M_443 , 1'h0 } )
		| ( { 2{ FL02_02_streg_t_c2 } } & FL02_02_streg_t1 ) ) ;
	end
assign	FL02_02_streg_en = ( FL02_02_streg_t_c1 | FL02_02_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL02_02_streg_en )
		FL02_02_streg <= FL02_02_streg_t ;
assign	M_450 = ( ST1_08d & ( ~FL02_03_break ) ) ;
assign	M_456 = ( ( ( U_111 & FJ_11_12 ) | ( U_114 & ( ~FL02_02_ndat ) ) ) | ( U_107 & ( 
	~FL02_02_ndat ) ) ) ;
always @ ( U_107 or FL02_02_ndat or U_114 or U_112 or M_456 or M_450 or ST1_07d or 
	U_147 )
	begin
	FL02_03_streg_t_c1 = ( ( U_147 | ST1_07d ) | ( M_450 & M_456 ) ) ;
	FL02_03_streg_t_c2 = ( M_450 & ( ( U_112 | ( U_114 & FL02_02_ndat ) ) | ( 
		U_107 & FL02_02_ndat ) ) ) ;
	FL02_03_streg_t = ( { 1{ FL02_03_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL02_03_streg_en = ( FL02_03_streg_t_c1 | FL02_03_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL02_03_streg_en )
		FL02_03_streg <= FL02_03_streg_t ;
assign	M_457 = ( ( U_121 & ( ~FL02_02_Lndat ) ) | ( U_117 & ( ~FL02_02_Lndat ) ) ) ;
always @ ( FL02_02_Lndat or U_117 or U_123 or FL02_05_ngo or U_118 or M_457 or ST1_08d or 
	ST1_07d )
	begin
	FL02_04_streg_t_c1 = ( ST1_07d | ( ST1_08d & M_457 ) ) ;
	FL02_04_streg_t_c2 = ( ST1_08d & ( ( ( U_118 & FL02_05_ngo ) | U_123 ) | 
		( U_117 & FL02_02_Lndat ) ) ) ;
	FL02_04_streg_t = ( { 1{ FL02_04_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL02_04_streg_en = ( FL02_04_streg_t_c1 | FL02_04_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL02_04_streg_en )
		FL02_04_streg <= FL02_04_streg_t ;
assign	M_458 = ( ( U_131 & ( ~FL02_04_ndat ) ) | ( U_125 & ( ~FL02_04_ndat ) ) ) ;
always @ ( U_125 or FL02_04_ndat or U_131 or U_130 or U_132 or M_458 or ST1_08d or 
	ST1_07d )
	begin
	FL02_05_streg_t_c1 = ( ST1_07d | ( ST1_08d & M_458 ) ) ;
	FL02_05_streg_t_c2 = ( ST1_08d & ( ( ( U_132 | U_130 ) | ( U_131 & FL02_04_ndat ) ) | 
		( U_125 & FL02_04_ndat ) ) ) ;
	FL02_05_streg_t = ( { 1{ FL02_05_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL02_05_streg_en = ( FL02_05_streg_t_c1 | FL02_05_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL02_05_streg_en )
		FL02_05_streg <= FL02_05_streg_t ;
assign	M_459 = ( ( U_139 & ( ~FL02_05_ndat ) ) | ( U_135 & ( ~FL02_05_ndat ) ) ) ;
always @ ( U_135 or FL02_05_ndat or U_139 or U_140 or M_459 or ST1_08d or ST1_07d )
	begin
	FL02_06_streg_t_c1 = ( ST1_07d | ( ST1_08d & M_459 ) ) ;
	FL02_06_streg_t_c2 = ( ST1_08d & ( ( U_140 | ( U_139 & FL02_05_ndat ) ) | 
		( U_135 & FL02_05_ndat ) ) ) ;
	FL02_06_streg_t = ( { 1{ FL02_06_streg_t_c2 } } & 1'h1 )
		 ;
	end
assign	FL02_06_streg_en = ( FL02_06_streg_t_c1 | FL02_06_streg_t_c2 ) ;
always @ ( posedge clk )
	if ( FL02_06_streg_en )
		FL02_06_streg <= FL02_06_streg_t ;
assign	FL02_05_ngo = ( U_130 | U_132 ) ;
assign	FL02_01_ndat = ( U_85 | U_75 ) ;
assign	FL02_02_ndat = U_105 ;
assign	FL02_02_Lrdy = U_94 ;
assign	FL02_02_Lndat = ( U_91 | U_99 ) ;
assign	FL02_04_rdy = ( U_123 | U_117 ) ;
assign	FL02_04_ndat = U_121 ;
assign	FL02_05_ndat = U_131 ;
assign	CMPS_FL_C2496_1_DO_v = ( U_61 & RG_15_02 ) ;
assign	jpeg_out_a00_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a00_r_en )
		jpeg_out_a00_r <= rl_rg00 ;
assign	jpeg_out_a01_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a01_r_en )
		jpeg_out_a01_r <= rl_rg01 ;
assign	jpeg_out_a02_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a02_r_en )
		jpeg_out_a02_r <= rl_rg02 ;
assign	jpeg_out_a03_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a03_r_en )
		jpeg_out_a03_r <= rl_rg03 ;
assign	jpeg_out_a04_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a04_r_en )
		jpeg_out_a04_r <= rl_rg04 ;
assign	jpeg_out_a05_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a05_r_en )
		jpeg_out_a05_r <= rl_rg05 ;
assign	jpeg_out_a06_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a06_r_en )
		jpeg_out_a06_r <= rl_rg06 ;
assign	jpeg_out_a07_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a07_r_en )
		jpeg_out_a07_r <= rl_rg07 ;
assign	jpeg_out_a08_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a08_r_en )
		jpeg_out_a08_r <= rl_rg08 ;
assign	jpeg_out_a09_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a09_r_en )
		jpeg_out_a09_r <= rl_rg09 ;
assign	jpeg_out_a10_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a10_r_en )
		jpeg_out_a10_r <= rl_rg10 ;
assign	jpeg_out_a11_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a11_r_en )
		jpeg_out_a11_r <= rl_rg11 ;
assign	jpeg_out_a12_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a12_r_en )
		jpeg_out_a12_r <= rl_rg12 ;
assign	jpeg_out_a13_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a13_r_en )
		jpeg_out_a13_r <= rl_rg13 ;
assign	jpeg_out_a14_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a14_r_en )
		jpeg_out_a14_r <= rl_rg14 ;
assign	jpeg_out_a15_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a15_r_en )
		jpeg_out_a15_r <= rl_rg15 ;
assign	jpeg_out_a16_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a16_r_en )
		jpeg_out_a16_r <= rl_rg16 ;
assign	jpeg_out_a17_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a17_r_en )
		jpeg_out_a17_r <= rl_rg17 ;
assign	jpeg_out_a18_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a18_r_en )
		jpeg_out_a18_r <= rl_rg18 ;
assign	jpeg_out_a19_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a19_r_en )
		jpeg_out_a19_r <= rl_rg19 ;
assign	jpeg_out_a20_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a20_r_en )
		jpeg_out_a20_r <= rl_rg20 ;
assign	jpeg_out_a21_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a21_r_en )
		jpeg_out_a21_r <= rl_rg21 ;
assign	jpeg_out_a22_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a22_r_en )
		jpeg_out_a22_r <= rl_rg22 ;
assign	jpeg_out_a23_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a23_r_en )
		jpeg_out_a23_r <= rl_rg23 ;
assign	jpeg_out_a24_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a24_r_en )
		jpeg_out_a24_r <= rl_rg24 ;
assign	jpeg_out_a25_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a25_r_en )
		jpeg_out_a25_r <= rl_rg25 ;
assign	jpeg_out_a26_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a26_r_en )
		jpeg_out_a26_r <= rl_rg26 ;
assign	jpeg_out_a27_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a27_r_en )
		jpeg_out_a27_r <= rl_rg27 ;
assign	jpeg_out_a28_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a28_r_en )
		jpeg_out_a28_r <= rl_rg28 ;
assign	jpeg_out_a29_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a29_r_en )
		jpeg_out_a29_r <= rl_rg29 ;
assign	jpeg_out_a30_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a30_r_en )
		jpeg_out_a30_r <= rl_rg30 ;
assign	jpeg_out_a31_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a31_r_en )
		jpeg_out_a31_r <= rl_rg31 ;
assign	jpeg_out_a32_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a32_r_en )
		jpeg_out_a32_r <= rl_rg32 ;
assign	jpeg_out_a33_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a33_r_en )
		jpeg_out_a33_r <= rl_rg33 ;
assign	jpeg_out_a34_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a34_r_en )
		jpeg_out_a34_r <= rl_rg34 ;
assign	jpeg_out_a35_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a35_r_en )
		jpeg_out_a35_r <= rl_rg35 ;
assign	jpeg_out_a36_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a36_r_en )
		jpeg_out_a36_r <= rl_rg36 ;
assign	jpeg_out_a37_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a37_r_en )
		jpeg_out_a37_r <= rl_rg37 ;
assign	jpeg_out_a38_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a38_r_en )
		jpeg_out_a38_r <= rl_rg38 ;
assign	jpeg_out_a39_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a39_r_en )
		jpeg_out_a39_r <= rl_rg39 ;
assign	jpeg_out_a40_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a40_r_en )
		jpeg_out_a40_r <= rl_rg40 ;
assign	jpeg_out_a41_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a41_r_en )
		jpeg_out_a41_r <= rl_rg41 ;
assign	jpeg_out_a42_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a42_r_en )
		jpeg_out_a42_r <= rl_rg42 ;
assign	jpeg_out_a43_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a43_r_en )
		jpeg_out_a43_r <= rl_rg43 ;
assign	jpeg_out_a44_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a44_r_en )
		jpeg_out_a44_r <= rl_rg44 ;
assign	jpeg_out_a45_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a45_r_en )
		jpeg_out_a45_r <= rl_rg45 ;
assign	jpeg_out_a46_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a46_r_en )
		jpeg_out_a46_r <= rl_rg46 ;
assign	jpeg_out_a47_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a47_r_en )
		jpeg_out_a47_r <= rl_rg47 ;
assign	jpeg_out_a48_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a48_r_en )
		jpeg_out_a48_r <= rl_rg48 ;
assign	jpeg_out_a49_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a49_r_en )
		jpeg_out_a49_r <= rl_rg49 ;
assign	jpeg_out_a50_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a50_r_en )
		jpeg_out_a50_r <= rl_rg50 ;
assign	jpeg_out_a51_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a51_r_en )
		jpeg_out_a51_r <= rl_rg51 ;
assign	jpeg_out_a52_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a52_r_en )
		jpeg_out_a52_r <= rl_rg52 ;
assign	jpeg_out_a53_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a53_r_en )
		jpeg_out_a53_r <= rl_rg53 ;
assign	jpeg_out_a54_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a54_r_en )
		jpeg_out_a54_r <= rl_rg54 ;
assign	jpeg_out_a55_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a55_r_en )
		jpeg_out_a55_r <= rl_rg55 ;
assign	jpeg_out_a56_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a56_r_en )
		jpeg_out_a56_r <= rl_rg56 ;
assign	jpeg_out_a57_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a57_r_en )
		jpeg_out_a57_r <= rl_rg57 ;
assign	jpeg_out_a58_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a58_r_en )
		jpeg_out_a58_r <= rl_rg58 ;
assign	jpeg_out_a59_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a59_r_en )
		jpeg_out_a59_r <= rl_rg59 ;
assign	jpeg_out_a60_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a60_r_en )
		jpeg_out_a60_r <= rl_rg60 ;
assign	jpeg_out_a61_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a61_r_en )
		jpeg_out_a61_r <= rl_rg61 ;
assign	jpeg_out_a62_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a62_r_en )
		jpeg_out_a62_r <= rl_rg62 ;
assign	jpeg_out_a63_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a63_r_en )
		jpeg_out_a63_r <= rl_rg63 ;
assign	jpeg_out_a64_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a64_r_en )
		jpeg_out_a64_r <= rl_rg64 ;
assign	jpeg_out_a65_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a65_r_en )
		jpeg_out_a65_r <= rl_rg65 ;
assign	jpeg_out_a66_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a66_r_en )
		jpeg_out_a66_r <= rl_rg66 ;
assign	jpeg_out_a67_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a67_r_en )
		jpeg_out_a67_r <= rl_rg67 ;
assign	jpeg_out_a68_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a68_r_en )
		jpeg_out_a68_r <= rl_rg68 ;
assign	jpeg_out_a69_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a69_r_en )
		jpeg_out_a69_r <= rl_rg69 ;
assign	jpeg_out_a70_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a70_r_en )
		jpeg_out_a70_r <= rl_rg70 ;
assign	jpeg_out_a71_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a71_r_en )
		jpeg_out_a71_r <= rl_rg71 ;
assign	jpeg_out_a72_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a72_r_en )
		jpeg_out_a72_r <= rl_rg72 ;
assign	jpeg_out_a73_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a73_r_en )
		jpeg_out_a73_r <= rl_rg73 ;
assign	jpeg_out_a74_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a74_r_en )
		jpeg_out_a74_r <= rl_rg74 ;
assign	jpeg_out_a75_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a75_r_en )
		jpeg_out_a75_r <= rl_rg75 ;
assign	jpeg_out_a76_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a76_r_en )
		jpeg_out_a76_r <= rl_rg76 ;
assign	jpeg_out_a77_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a77_r_en )
		jpeg_out_a77_r <= rl_rg77 ;
assign	jpeg_out_a78_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a78_r_en )
		jpeg_out_a78_r <= rl_rg78 ;
assign	jpeg_out_a79_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a79_r_en )
		jpeg_out_a79_r <= rl_rg79 ;
assign	jpeg_out_a80_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a80_r_en )
		jpeg_out_a80_r <= rl_rg80 ;
assign	jpeg_out_a81_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a81_r_en )
		jpeg_out_a81_r <= rl_rg81 ;
assign	jpeg_out_a82_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a82_r_en )
		jpeg_out_a82_r <= rl_rg82 ;
assign	jpeg_out_a83_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a83_r_en )
		jpeg_out_a83_r <= rl_rg83 ;
assign	jpeg_out_a84_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a84_r_en )
		jpeg_out_a84_r <= rl_rg84 ;
assign	jpeg_out_a85_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a85_r_en )
		jpeg_out_a85_r <= rl_rg85 ;
assign	jpeg_out_a86_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a86_r_en )
		jpeg_out_a86_r <= rl_rg86 ;
assign	jpeg_out_a87_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a87_r_en )
		jpeg_out_a87_r <= rl_rg87 ;
assign	jpeg_out_a88_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a88_r_en )
		jpeg_out_a88_r <= rl_rg88 ;
assign	jpeg_out_a89_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a89_r_en )
		jpeg_out_a89_r <= rl_rg89 ;
assign	jpeg_out_a90_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a90_r_en )
		jpeg_out_a90_r <= rl_rg90 ;
assign	jpeg_out_a91_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a91_r_en )
		jpeg_out_a91_r <= rl_rg91 ;
assign	jpeg_out_a92_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a92_r_en )
		jpeg_out_a92_r <= rl_rg92 ;
assign	jpeg_out_a93_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a93_r_en )
		jpeg_out_a93_r <= rl_rg93 ;
assign	jpeg_out_a94_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a94_r_en )
		jpeg_out_a94_r <= rl_rg94 ;
assign	jpeg_out_a95_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a95_r_en )
		jpeg_out_a95_r <= rl_rg95 ;
assign	jpeg_out_a96_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a96_r_en )
		jpeg_out_a96_r <= rl_rg96 ;
assign	jpeg_out_a97_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a97_r_en )
		jpeg_out_a97_r <= rl_rg97 ;
assign	jpeg_out_a98_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a98_r_en )
		jpeg_out_a98_r <= rl_rg98 ;
assign	jpeg_out_a99_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a99_r_en )
		jpeg_out_a99_r <= rl_rg99 ;
assign	jpeg_out_a100_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a100_r_en )
		jpeg_out_a100_r <= rl_rg100 ;
assign	jpeg_out_a101_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a101_r_en )
		jpeg_out_a101_r <= rl_rg101 ;
assign	jpeg_out_a102_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a102_r_en )
		jpeg_out_a102_r <= rl_rg102 ;
assign	jpeg_out_a103_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a103_r_en )
		jpeg_out_a103_r <= rl_rg103 ;
assign	jpeg_out_a104_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a104_r_en )
		jpeg_out_a104_r <= rl_rg104 ;
assign	jpeg_out_a105_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a105_r_en )
		jpeg_out_a105_r <= rl_rg105 ;
assign	jpeg_out_a106_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a106_r_en )
		jpeg_out_a106_r <= rl_rg106 ;
assign	jpeg_out_a107_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a107_r_en )
		jpeg_out_a107_r <= rl_rg107 ;
assign	jpeg_out_a108_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a108_r_en )
		jpeg_out_a108_r <= rl_rg108 ;
assign	jpeg_out_a109_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a109_r_en )
		jpeg_out_a109_r <= rl_rg109 ;
assign	jpeg_out_a110_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a110_r_en )
		jpeg_out_a110_r <= rl_rg110 ;
assign	jpeg_out_a111_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a111_r_en )
		jpeg_out_a111_r <= rl_rg111 ;
assign	jpeg_out_a112_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a112_r_en )
		jpeg_out_a112_r <= rl_rg112 ;
assign	jpeg_out_a113_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a113_r_en )
		jpeg_out_a113_r <= rl_rg113 ;
assign	jpeg_out_a114_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a114_r_en )
		jpeg_out_a114_r <= rl_rg114 ;
assign	jpeg_out_a115_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a115_r_en )
		jpeg_out_a115_r <= rl_rg115 ;
assign	jpeg_out_a116_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a116_r_en )
		jpeg_out_a116_r <= rl_rg116 ;
assign	jpeg_out_a117_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a117_r_en )
		jpeg_out_a117_r <= rl_rg117 ;
assign	jpeg_out_a118_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a118_r_en )
		jpeg_out_a118_r <= rl_rg118 ;
assign	jpeg_out_a119_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a119_r_en )
		jpeg_out_a119_r <= rl_rg119 ;
assign	jpeg_out_a120_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a120_r_en )
		jpeg_out_a120_r <= rl_rg120 ;
assign	jpeg_out_a121_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a121_r_en )
		jpeg_out_a121_r <= rl_rg121 ;
assign	jpeg_out_a122_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a122_r_en )
		jpeg_out_a122_r <= rl_rg122 ;
assign	jpeg_out_a123_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a123_r_en )
		jpeg_out_a123_r <= rl_rg123 ;
assign	jpeg_out_a124_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a124_r_en )
		jpeg_out_a124_r <= rl_rg124 ;
assign	jpeg_out_a125_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a125_r_en )
		jpeg_out_a125_r <= rl_rg125 ;
assign	jpeg_out_a126_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a126_r_en )
		jpeg_out_a126_r <= rl_rg126 ;
assign	jpeg_out_a127_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a127_r_en )
		jpeg_out_a127_r <= rl_rg127 ;
assign	jpeg_len_out_r_en = U_164 ;
always @ ( posedge clk )	// line#=../rle.cpp:93
	if ( jpeg_len_out_r_en )
		jpeg_len_out_r <= { 4'h0 , RG_len_05 } ;
always @ ( U_164 )
	valid_r_t = ( { 1{ U_164 } } & 1'h1 )	// line#=../rle.cpp:95
		 ;	// line#=../rle.cpp:30
assign	valid_r_en = ( ST1_01d | U_164 ) ;
always @ ( posedge clk )
	if ( valid_r_en )
		valid_r <= valid_r_t ;	// line#=../rle.cpp:30,95
assign	sub8u1i1 = { ( ST1_15d & RG_len_05 [7] ) , RG_len_05 [6:0] } ;	// line#=../rle.cpp:77,78,83,84,86
always @ ( U_165 or ST1_13d or ST1_15d or ST1_10d )
	begin
	sub8u1i2_c1 = ( ST1_10d | ST1_15d ) ;	// line#=../rle.cpp:77,78,86
	sub8u1i2 = ( ( { 3{ sub8u1i2_c1 } } & 3'h2 )	// line#=../rle.cpp:77,78,86
		| ( { 3{ ST1_13d } } & 3'h4 )		// line#=../rle.cpp:83,84
		| ( { 3{ U_165 } } & 3'h3 )		// line#=../rle.cpp:83,84
		) ;
	end
always @ ( RG_y_02 or U_10 or RG_j_x_02 or ST1_02d )
	incr4s1i1 = ( ( { 4{ ST1_02d } } & RG_j_x_02 )	// line#=../rle.cpp:34
		| ( { 4{ U_10 } } & RG_y_02 )		// line#=../rle.cpp:44
		) ;
assign	incr8u1i1 = RG_len_05 ;	// line#=../rle.cpp:68,73,79,80
assign	incr8u2i1 = incr8u1ot ;	// line#=../rle.cpp:68,69,73,74
assign	incr32s1i1 = RG_j_k ;	// line#=../rle.cpp:61,62,64,114,125,145
				// ,156
assign	incr32s2i1 = RG_i ;	// line#=../rle.cpp:61,62,63,119,129,150
				// ,160
assign	decr32s1i1 = RG_i ;	// line#=../rle.cpp:124,155
assign	decr32s2i1 = RG_j_k ;	// line#=../rle.cpp:130,161
always @ ( RG_i or U_59 or RG_i_04 or U_70 )	// line#=../rle.cpp:140,141
	zz_RA1 = ( ( { 6{ U_70 } } & RG_i_04 [5:0] )	// line#=../rle.cpp:74
		| ( { 6{ U_59 } } & RG_i [5:0] )	// line#=../rle.cpp:61,62
		) ;	// line#=../rle.cpp:52,53
always @ ( RG_k_05 or U_44 or RG_k or U_34 )
	zz_WA2 = ( ( { 6{ U_34 } } & RG_k )		// line#=../rle.cpp:111
		| ( { 6{ U_44 } } & RG_k_05 [5:0] )	// line#=../rle.cpp:142
		) ;
assign	zz_WE2 = ( U_34 | U_44 ) ;
always @ ( sub8u1ot or ST1_13d or U_165 or ST1_10d or decr8u_71ot or ST1_09d )
	begin
	rl_ad00_c1 = ( ( ST1_10d | U_165 ) | ST1_13d ) ;	// line#=../rle.cpp:77,78,83,84
	rl_ad00 = ( ( { 7{ ST1_09d } } & decr8u_71ot )		// line#=../rle.cpp:77,78
		| ( { 7{ rl_ad00_c1 } } & sub8u1ot [6:0] )	// line#=../rle.cpp:77,78,83,84
		) ;
	end
assign	rl_ad01 = RG_k_05 ;	// line#=../rle.cpp:69,74,85
assign	rl_ad02 = RG_len_05 [6:0] ;	// line#=../rle.cpp:68,73,79,80
jpeg_CMPS_FL_C2603 #(9) CMPS_FL_C2603_1 ( .CLOCK(clk) ,.RESET(rst) ,.DO(zz_RD1) ,
	.DO_v(U_74) ,.AD_v(U_70) ,.FL_RESET(ST1_07d) ,.DO_t(CMPS_FL_C2603_1_DO_t) );
always @ ( CMPS_FL_C2603_1_DO_t or U_74 )
	rl_wd01 = ( { 9{ U_74 } } & CMPS_FL_C2603_1_DO_t )	// line#=../rle.cpp:74
		 ;	// line#=../rle.cpp:69,85
always @ ( RG_k_04 or U_70 )
	rl_wd02 = ( { 9{ U_70 } } & RG_k_04 )	// line#=../rle.cpp:73
		 ;	// line#=../rle.cpp:68,79,80
assign	rl_we01 = ( U_72 | ST1_15d ) ;	// line#=../rle.cpp:69,74,85
assign	M_454 = U_68 ;
assign	rl_we02 = ( ( M_454 | U_159 ) | ST1_12d ) ;	// line#=../rle.cpp:68,73,79,80

endmodule

module jpeg_incr8u_6 ( i1 ,o1 );
input	[5:0]	i1 ;
output	[5:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr8u_7 ( i1 ,o1 );
input	[5:0]	i1 ;
output	[6:0]	o1 ;

assign	o1 = ( { 1'h0 , i1 } + 1'h1 ) ;

endmodule

module jpeg_decr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_decr8u_7 ( i1 ,o1 );
input	[6:0]	i1 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_incr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr8u ( i1 ,o1 );
input	[7:0]	i1 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr4s ( i1 ,o1 );
input	[3:0]	i1 ;
output	[3:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr3u ( i1 ,o1 );
input	[2:0]	i1 ;
output	[3:0]	o1 ;

assign	o1 = ( { 1'h0 , i1 } + 1'h1 ) ;

endmodule

module jpeg_lop8u_1 ( i1 ,i2 ,o1 );
input	[5:0]	i1 ;
input	[5:0]	i2 ;
output		o1 ;
wire		M_01 ;

assign	M_01 = ( i1 < i2 ) ;
assign	o1 = M_01 ;

endmodule

module jpeg_sub12s_9 ( i1 ,i2 ,o1 );
input	[8:0]	i1 ;
input	[8:0]	i2 ;
output	[8:0]	o1 ;

assign	o1 = ( i1 - i2 ) ;

endmodule

module jpeg_sub8u ( i1 ,i2 ,o1 );
input	[7:0]	i1 ;
input	[2:0]	i2 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 - { 5'h00 , i2 } ) ;

endmodule

module jpeg_add3u ( i1 ,i2 ,o1 );
input	[2:0]	i1 ;
input		i2 ;
output	[3:0]	o1 ;

assign	o1 = ( { 1'h0 , i1 } + { 3'h0 , i2 } ) ;

endmodule

module jpeg_decoder_6to64 ( DECODER_in ,DECODER_out );
input	[5:0]	DECODER_in ;
output	[63:0]	DECODER_out ;
reg	[63:0]	DECODER_out ;

always @ ( DECODER_in )
	begin
	DECODER_out = 64'h0000000000000000 ;
	DECODER_out [63 - DECODER_in] = 1'h1 ;
	end

endmodule

module jpeg_decoder_7to128 ( DECODER_in ,DECODER_out );
input	[6:0]	DECODER_in ;
output	[127:0]	DECODER_out ;
reg	[127:0]	DECODER_out ;

always @ ( DECODER_in )
	begin
	DECODER_out = 128'h00000000000000000000000000000000 ;
	DECODER_out [127 - DECODER_in] = 1'h1 ;
	end

endmodule

module jpeg_CMPS_FL_C2496 #(parameter DATA_BITW = 8)
   ( CLOCK ,
     RESET ,
     DO ,DO_v ,AD_v ,FL_RESET ,DO_t );
   input  CLOCK ;
   input  RESET ;
   input [DATA_BITW-1:0] DO ;
   input                 DO_v ;
   input                 AD_v ;
   input                 FL_RESET ;
   output [DATA_BITW-1:0] DO_t ;

   jpeg_CMPS_FL_C2496_sub #(DATA_BITW)
   jpeg_CMPS_FL_C2496_sub_1 ( .CLOCK(CLOCK) ,
        .RESET(RESET) ,
        .DO(DO) ,.DO_v(DO_v) , .AD_v(AD_v) ,.STALL(1'b0) ,
        .FL_RESET(FL_RESET) ,.DO_t(DO_t) );

endmodule

module jpeg_CMPS_FL_C2496_sub #(parameter DATA_BITW = 8)
   ( CLOCK ,
     RESET ,
     DO ,DO_v ,AD_v ,STALL ,FL_RESET ,DO_t );
   input  CLOCK ;
   input  RESET ;
   input [DATA_BITW-1:0] DO ;
   input                 DO_v ;
   input                 AD_v ;
   input                 STALL ;
   input                 FL_RESET ;
   output [DATA_BITW-1:0] DO_t ;

   wire                   enq ;
   wire                   deq ;
   wire                   queue_v ;
   reg [DATA_BITW-1:0]    q_s;
   wire [DATA_BITW-1:0]   q_s_t;
   reg                    q_s_f ;
   wire                   q_s_f_t ;
   reg                    rg_s ;
   reg [DATA_BITW-1:0]    DO_t ;
   assign enq = ( ( ( ~queue_v ) | q_s_f ) & ( rg_s ) ) ;
   assign deq = ( queue_v & q_s_f ) ;
   assign q_s_f_t = q_s_f;
   assign q_s_t = q_s;

   always @ ( posedge CLOCK )
     if ( !RESET )
       q_s <= {DATA_BITW {1'b0}} ;
     else begin
       case ( { ( ( deq & ( ~enq ) ) | FL_RESET )  ,
                ( enq & ( ~q_s_f ) )  } )
         2'b10 :
           q_s <= {DATA_BITW {1'b0}} ;
         2'b01 :
           q_s <= DO ;
         default :
           q_s <= q_s_t ;
       endcase
     end

   always @ ( posedge CLOCK )
     if ( !RESET )
       q_s_f <= 1'h0 ;
     else  begin
       case ( { ( ( deq & ( ~enq ) ) | FL_RESET ) ,
                ( enq & ( ~q_s_f ) )  } )
         2'b10 :
           q_s_f <= 1'h0 ;
         2'b01 :
           q_s_f <= 1'h1 ;
         default :
           q_s_f <= q_s_f_t ;
       endcase
     end

   assign queue_v = ( DO_v & ( ~STALL ) ) ;

   always @ ( posedge CLOCK ) begin
      if ( !RESET )
        rg_s <= 1'h0 ;
      else
        rg_s <= ( ~( ( ( ~AD_v ) | STALL ) | FL_RESET ) ) ;
   end

   always @ ( q_s or q_s_f or DO )
     begin
       case ( {~q_s_f} )
         1'b1 :
           DO_t = DO ;
         1'b0 :
           DO_t = q_s ;
         default :
           DO_t = {DATA_BITW {1'bx}} ;
       endcase
     end

endmodule

module jpeg_CMPS_FL_C2603 #(parameter DATA_BITW = 8)
   ( CLOCK ,
     RESET ,
     DO ,DO_v ,AD_v ,FL_RESET ,DO_t );
   input  CLOCK ;
   input  RESET ;
   input [DATA_BITW-1:0] DO ;
   input                 DO_v ;
   input                 AD_v ;
   input                 FL_RESET ;
   output [DATA_BITW-1:0] DO_t ;

   jpeg_CMPS_FL_C2603_sub #(DATA_BITW)
   jpeg_CMPS_FL_C2603_sub_1 ( .CLOCK(CLOCK) ,
        .RESET(RESET) ,
        .DO(DO) ,.DO_v(DO_v) , .AD_v(AD_v) ,.STALL(1'b0) ,
        .FL_RESET(FL_RESET) ,.DO_t(DO_t) );

endmodule

module jpeg_CMPS_FL_C2603_sub #(parameter DATA_BITW = 8)
   ( CLOCK ,
     RESET ,
     DO ,DO_v ,AD_v ,STALL ,FL_RESET ,DO_t );
   input  CLOCK ;
   input  RESET ;
   input [DATA_BITW-1:0] DO ;
   input                 DO_v ;
   input                 AD_v ;
   input                 STALL ;
   input                 FL_RESET ;
   output [DATA_BITW-1:0] DO_t ;

   wire                   enq ;
   wire                   deq ;
   wire                   queue_v ;
   reg [DATA_BITW-1:0]    q_s;
   wire [DATA_BITW-1:0]   q_s_t;
   reg                    q_s_f ;
   wire                   q_s_f_t ;
   reg                    rg_s ;
   reg [DATA_BITW-1:0]    DO_t ;
   assign enq = ( ( ( ~queue_v ) | q_s_f ) & ( rg_s ) ) ;
   assign deq = ( queue_v & q_s_f ) ;
   assign q_s_f_t = q_s_f;
   assign q_s_t = q_s;

   always @ ( posedge CLOCK )
     if ( !RESET )
       q_s <= {DATA_BITW {1'b0}} ;
     else begin
       case ( { ( ( deq & ( ~enq ) ) | FL_RESET )  ,
                ( enq & ( ~q_s_f ) )  } )
         2'b10 :
           q_s <= {DATA_BITW {1'b0}} ;
         2'b01 :
           q_s <= DO ;
         default :
           q_s <= q_s_t ;
       endcase
     end

   always @ ( posedge CLOCK )
     if ( !RESET )
       q_s_f <= 1'h0 ;
     else  begin
       case ( { ( ( deq & ( ~enq ) ) | FL_RESET ) ,
                ( enq & ( ~q_s_f ) )  } )
         2'b10 :
           q_s_f <= 1'h0 ;
         2'b01 :
           q_s_f <= 1'h1 ;
         default :
           q_s_f <= q_s_f_t ;
       endcase
     end

   assign queue_v = ( DO_v & ( ~STALL ) ) ;

   always @ ( posedge CLOCK ) begin
      if ( !RESET )
        rg_s <= 1'h0 ;
      else
        rg_s <= ( ~( ( ( ~AD_v ) | STALL ) | FL_RESET ) ) ;
   end

   always @ ( q_s or q_s_f or DO )
     begin
       case ( {~q_s_f} )
         1'b1 :
           DO_t = DO ;
         1'b0 :
           DO_t = q_s ;
         default :
           DO_t = {DATA_BITW {1'bx}} ;
       endcase
     end

endmodule

module jpeg_MEMB9W64 ( RA1 ,RD1 ,RCLK1 ,WA2 ,WD2 ,WE2 ,WCLK2 );
input	[5:0]	RA1 ;
output	[8:0]	RD1 ;
input		RCLK1 ;
input	[5:0]	WA2 ;
input	[8:0]	WD2 ;
input		WE2 ;
input		WCLK2 ;

jpeg_MEMB9W64_sub INST_MEMB9W64_sub_1 ( .RD1(RD1) ,.WE2(WE2) ,.WD2(WD2) ,.RA1(RA1) ,
	.WA2(WA2) ,.RCLK1(RCLK1) ,.WCLK2(WCLK2) );

endmodule

(* ram_extract = "yes" *)
module jpeg_MEMB9W64_sub ( RD1 ,WE2 ,WD2 ,RA1 ,WA2 ,RCLK1 ,WCLK2 );
output	[8:0]	RD1 ;
input		WE2 ;
input	[8:0]	WD2 ;
input	[5:0]	RA1 ;
input	[5:0]	WA2 ;
input		RCLK1 ;
input		WCLK2 ;
wire		Wen1_wire ;
reg	[8:0]	Rd1_sr	[0:0] ;
(* ram_style = "block" *)reg	[8:0]	MEMB9W64_r	[0:63] ;

assign	RD1 = Rd1_sr[0] ;
assign	Wen1_wire = WE2 ;

always @ ( posedge RCLK1 )
	begin
	Rd1_sr [0] <= MEMB9W64_r[RA1] ;
	end

always @ ( posedge WCLK2 )
	begin
	if ( Wen1_wire )
		begin
		MEMB9W64_r [WA2] <= WD2 ;
		end
	end

endmodule
