// verilog_out version 6.79.2
// options:  veriloggen jpeg_E.IFF
// bdlpars options:  -DDSE ../rle.cpp
// bdltran options:  -c1000 -s -Zresource_fcnt=GENERATE -Zresource_mcnt=GENERATE -lb /home/shuangnan/share/packages/zynq-1.BLIB -lfl /home/shuangnan/share/packages/zynq-1.FLIB jpeg.IFF -OX -a8196 -Zfu_cnt_incr_rate=0 -tcio 
// timestamp_0: 20180213182241_17595_01259
// timestamp_5: 20180213182246_18930_09871
// timestamp_9: 20180213182506_18930_37026
// timestamp_C: 20180213182501_18930_01793
// timestamp_E: 20180213182512_18930_82825
// timestamp_V: 20180213182533_19076_78847

module jpeg ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,jpeg_in_a04 ,
	jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,jpeg_in_a10 ,
	jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,jpeg_in_a16 ,
	jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,jpeg_in_a22 ,
	jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,jpeg_in_a28 ,
	jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,jpeg_in_a34 ,
	jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,jpeg_in_a40 ,
	jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,jpeg_in_a46 ,
	jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,jpeg_in_a52 ,
	jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,jpeg_in_a58 ,
	jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,jpeg_in_a64 ,
	jpeg_in_a65 ,jpeg_in_a66 ,jpeg_in_a67 ,jpeg_in_a68 ,jpeg_in_a69 ,jpeg_in_a70 ,
	jpeg_in_a71 ,jpeg_in_a72 ,jpeg_in_a73 ,jpeg_in_a74 ,jpeg_in_a75 ,jpeg_in_a76 ,
	jpeg_in_a77 ,jpeg_in_a78 ,jpeg_in_a79 ,jpeg_in_a80 ,jpeg_in_a81 ,jpeg_in_a82 ,
	jpeg_in_a83 ,jpeg_in_a84 ,jpeg_in_a85 ,jpeg_in_a86 ,jpeg_in_a87 ,jpeg_in_a88 ,
	jpeg_in_a89 ,jpeg_in_a90 ,jpeg_in_a91 ,jpeg_in_a92 ,jpeg_in_a93 ,jpeg_in_a94 ,
	jpeg_in_a95 ,jpeg_in_a96 ,jpeg_in_a97 ,jpeg_in_a98 ,jpeg_in_a99 ,jpeg_in_a100 ,
	jpeg_in_a101 ,jpeg_in_a102 ,jpeg_in_a103 ,jpeg_in_a104 ,jpeg_in_a105 ,jpeg_in_a106 ,
	jpeg_in_a107 ,jpeg_in_a108 ,jpeg_in_a109 ,jpeg_in_a110 ,jpeg_in_a111 ,jpeg_in_a112 ,
	jpeg_in_a113 ,jpeg_in_a114 ,jpeg_in_a115 ,jpeg_in_a116 ,jpeg_in_a117 ,jpeg_in_a118 ,
	jpeg_in_a119 ,jpeg_in_a120 ,jpeg_in_a121 ,jpeg_in_a122 ,jpeg_in_a123 ,jpeg_in_a124 ,
	jpeg_in_a125 ,jpeg_in_a126 ,jpeg_in_a127 ,jpeg_len_in ,jpeg_out_a00 ,jpeg_out_a01 ,
	jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,jpeg_out_a06 ,jpeg_out_a07 ,
	jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,jpeg_out_a12 ,jpeg_out_a13 ,
	jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,jpeg_out_a18 ,jpeg_out_a19 ,
	jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,jpeg_out_a24 ,jpeg_out_a25 ,
	jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,jpeg_out_a30 ,jpeg_out_a31 ,
	jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,jpeg_out_a36 ,jpeg_out_a37 ,
	jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,jpeg_out_a42 ,jpeg_out_a43 ,
	jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,jpeg_out_a48 ,jpeg_out_a49 ,
	jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,jpeg_out_a54 ,jpeg_out_a55 ,
	jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,jpeg_out_a60 ,jpeg_out_a61 ,
	jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,jpeg_out_a66 ,jpeg_out_a67 ,
	jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,jpeg_out_a72 ,jpeg_out_a73 ,
	jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,jpeg_out_a78 ,jpeg_out_a79 ,
	jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,jpeg_out_a84 ,jpeg_out_a85 ,
	jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,jpeg_out_a90 ,jpeg_out_a91 ,
	jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,jpeg_out_a96 ,jpeg_out_a97 ,
	jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,jpeg_out_a102 ,
	jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,jpeg_out_a107 ,
	jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,jpeg_out_a112 ,
	jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,jpeg_out_a117 ,
	jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,jpeg_out_a122 ,
	jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,jpeg_out_a127 ,
	jpeg_len_out ,valid );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a64 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a65 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a66 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a67 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a68 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a69 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a70 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a71 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a72 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a73 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a74 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a75 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a76 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a77 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a78 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a79 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a80 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a81 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a82 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a83 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a84 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a85 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a86 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a87 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a88 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a89 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a90 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a91 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a92 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a93 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a94 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a95 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a96 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a97 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a98 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a99 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a100 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a101 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a102 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a103 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a104 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a105 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a106 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a107 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a108 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a109 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a110 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a111 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a112 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a113 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a114 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a115 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a116 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a117 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a118 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a119 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a120 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a121 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a122 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a123 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a124 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a125 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a126 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a127 ;	// line#=../rle.h:56
input	[11:0]	jpeg_len_in ;	// line#=../rle.h:57
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
wire		ST1_01d ;
wire		ST1_02d ;
wire		ST1_03d ;
wire		ST1_04d ;
wire		ST1_05d ;
wire		ST1_06d ;
wire		ST1_07d ;
wire		ST1_08d ;
wire		ST1_09d ;
wire		ST1_10d ;
wire		ST1_11d ;
wire		JF_01 ;
wire		lop8u_11ot ;
wire		JF_03 ;
wire		CT_33 ;
wire		RG_315 ;
wire		JF_06 ;

jpeg_fsm INST_fsm ( .clk(clk) ,.rst(rst) ,.ST1_11d(ST1_11d) ,.ST1_10d(ST1_10d) ,
	.ST1_09d(ST1_09d) ,.ST1_08d(ST1_08d) ,.ST1_07d(ST1_07d) ,.ST1_06d(ST1_06d) ,
	.ST1_05d(ST1_05d) ,.ST1_04d(ST1_04d) ,.ST1_03d(ST1_03d) ,.ST1_02d(ST1_02d) ,
	.ST1_01d(ST1_01d) ,.JF_01(JF_01) ,.lop8u_11ot(lop8u_11ot) ,.JF_03(JF_03) ,
	.CT_33(CT_33) ,.RG_315(RG_315) ,.JF_06(JF_06) );
jpeg_dat INST_dat ( .clk(clk) ,.rst(rst) ,.jpeg_in_a00(jpeg_in_a00) ,.jpeg_in_a01(jpeg_in_a01) ,
	.jpeg_in_a02(jpeg_in_a02) ,.jpeg_in_a03(jpeg_in_a03) ,.jpeg_in_a04(jpeg_in_a04) ,
	.jpeg_in_a05(jpeg_in_a05) ,.jpeg_in_a06(jpeg_in_a06) ,.jpeg_in_a07(jpeg_in_a07) ,
	.jpeg_in_a08(jpeg_in_a08) ,.jpeg_in_a09(jpeg_in_a09) ,.jpeg_in_a10(jpeg_in_a10) ,
	.jpeg_in_a11(jpeg_in_a11) ,.jpeg_in_a12(jpeg_in_a12) ,.jpeg_in_a13(jpeg_in_a13) ,
	.jpeg_in_a14(jpeg_in_a14) ,.jpeg_in_a15(jpeg_in_a15) ,.jpeg_in_a16(jpeg_in_a16) ,
	.jpeg_in_a17(jpeg_in_a17) ,.jpeg_in_a18(jpeg_in_a18) ,.jpeg_in_a19(jpeg_in_a19) ,
	.jpeg_in_a20(jpeg_in_a20) ,.jpeg_in_a21(jpeg_in_a21) ,.jpeg_in_a22(jpeg_in_a22) ,
	.jpeg_in_a23(jpeg_in_a23) ,.jpeg_in_a24(jpeg_in_a24) ,.jpeg_in_a25(jpeg_in_a25) ,
	.jpeg_in_a26(jpeg_in_a26) ,.jpeg_in_a27(jpeg_in_a27) ,.jpeg_in_a28(jpeg_in_a28) ,
	.jpeg_in_a29(jpeg_in_a29) ,.jpeg_in_a30(jpeg_in_a30) ,.jpeg_in_a31(jpeg_in_a31) ,
	.jpeg_in_a32(jpeg_in_a32) ,.jpeg_in_a33(jpeg_in_a33) ,.jpeg_in_a34(jpeg_in_a34) ,
	.jpeg_in_a35(jpeg_in_a35) ,.jpeg_in_a36(jpeg_in_a36) ,.jpeg_in_a37(jpeg_in_a37) ,
	.jpeg_in_a38(jpeg_in_a38) ,.jpeg_in_a39(jpeg_in_a39) ,.jpeg_in_a40(jpeg_in_a40) ,
	.jpeg_in_a41(jpeg_in_a41) ,.jpeg_in_a42(jpeg_in_a42) ,.jpeg_in_a43(jpeg_in_a43) ,
	.jpeg_in_a44(jpeg_in_a44) ,.jpeg_in_a45(jpeg_in_a45) ,.jpeg_in_a46(jpeg_in_a46) ,
	.jpeg_in_a47(jpeg_in_a47) ,.jpeg_in_a48(jpeg_in_a48) ,.jpeg_in_a49(jpeg_in_a49) ,
	.jpeg_in_a50(jpeg_in_a50) ,.jpeg_in_a51(jpeg_in_a51) ,.jpeg_in_a52(jpeg_in_a52) ,
	.jpeg_in_a53(jpeg_in_a53) ,.jpeg_in_a54(jpeg_in_a54) ,.jpeg_in_a55(jpeg_in_a55) ,
	.jpeg_in_a56(jpeg_in_a56) ,.jpeg_in_a57(jpeg_in_a57) ,.jpeg_in_a58(jpeg_in_a58) ,
	.jpeg_in_a59(jpeg_in_a59) ,.jpeg_in_a60(jpeg_in_a60) ,.jpeg_in_a61(jpeg_in_a61) ,
	.jpeg_in_a62(jpeg_in_a62) ,.jpeg_in_a63(jpeg_in_a63) ,.jpeg_out_a00(jpeg_out_a00) ,
	.jpeg_out_a01(jpeg_out_a01) ,.jpeg_out_a02(jpeg_out_a02) ,.jpeg_out_a03(jpeg_out_a03) ,
	.jpeg_out_a04(jpeg_out_a04) ,.jpeg_out_a05(jpeg_out_a05) ,.jpeg_out_a06(jpeg_out_a06) ,
	.jpeg_out_a07(jpeg_out_a07) ,.jpeg_out_a08(jpeg_out_a08) ,.jpeg_out_a09(jpeg_out_a09) ,
	.jpeg_out_a10(jpeg_out_a10) ,.jpeg_out_a11(jpeg_out_a11) ,.jpeg_out_a12(jpeg_out_a12) ,
	.jpeg_out_a13(jpeg_out_a13) ,.jpeg_out_a14(jpeg_out_a14) ,.jpeg_out_a15(jpeg_out_a15) ,
	.jpeg_out_a16(jpeg_out_a16) ,.jpeg_out_a17(jpeg_out_a17) ,.jpeg_out_a18(jpeg_out_a18) ,
	.jpeg_out_a19(jpeg_out_a19) ,.jpeg_out_a20(jpeg_out_a20) ,.jpeg_out_a21(jpeg_out_a21) ,
	.jpeg_out_a22(jpeg_out_a22) ,.jpeg_out_a23(jpeg_out_a23) ,.jpeg_out_a24(jpeg_out_a24) ,
	.jpeg_out_a25(jpeg_out_a25) ,.jpeg_out_a26(jpeg_out_a26) ,.jpeg_out_a27(jpeg_out_a27) ,
	.jpeg_out_a28(jpeg_out_a28) ,.jpeg_out_a29(jpeg_out_a29) ,.jpeg_out_a30(jpeg_out_a30) ,
	.jpeg_out_a31(jpeg_out_a31) ,.jpeg_out_a32(jpeg_out_a32) ,.jpeg_out_a33(jpeg_out_a33) ,
	.jpeg_out_a34(jpeg_out_a34) ,.jpeg_out_a35(jpeg_out_a35) ,.jpeg_out_a36(jpeg_out_a36) ,
	.jpeg_out_a37(jpeg_out_a37) ,.jpeg_out_a38(jpeg_out_a38) ,.jpeg_out_a39(jpeg_out_a39) ,
	.jpeg_out_a40(jpeg_out_a40) ,.jpeg_out_a41(jpeg_out_a41) ,.jpeg_out_a42(jpeg_out_a42) ,
	.jpeg_out_a43(jpeg_out_a43) ,.jpeg_out_a44(jpeg_out_a44) ,.jpeg_out_a45(jpeg_out_a45) ,
	.jpeg_out_a46(jpeg_out_a46) ,.jpeg_out_a47(jpeg_out_a47) ,.jpeg_out_a48(jpeg_out_a48) ,
	.jpeg_out_a49(jpeg_out_a49) ,.jpeg_out_a50(jpeg_out_a50) ,.jpeg_out_a51(jpeg_out_a51) ,
	.jpeg_out_a52(jpeg_out_a52) ,.jpeg_out_a53(jpeg_out_a53) ,.jpeg_out_a54(jpeg_out_a54) ,
	.jpeg_out_a55(jpeg_out_a55) ,.jpeg_out_a56(jpeg_out_a56) ,.jpeg_out_a57(jpeg_out_a57) ,
	.jpeg_out_a58(jpeg_out_a58) ,.jpeg_out_a59(jpeg_out_a59) ,.jpeg_out_a60(jpeg_out_a60) ,
	.jpeg_out_a61(jpeg_out_a61) ,.jpeg_out_a62(jpeg_out_a62) ,.jpeg_out_a63(jpeg_out_a63) ,
	.jpeg_out_a64(jpeg_out_a64) ,.jpeg_out_a65(jpeg_out_a65) ,.jpeg_out_a66(jpeg_out_a66) ,
	.jpeg_out_a67(jpeg_out_a67) ,.jpeg_out_a68(jpeg_out_a68) ,.jpeg_out_a69(jpeg_out_a69) ,
	.jpeg_out_a70(jpeg_out_a70) ,.jpeg_out_a71(jpeg_out_a71) ,.jpeg_out_a72(jpeg_out_a72) ,
	.jpeg_out_a73(jpeg_out_a73) ,.jpeg_out_a74(jpeg_out_a74) ,.jpeg_out_a75(jpeg_out_a75) ,
	.jpeg_out_a76(jpeg_out_a76) ,.jpeg_out_a77(jpeg_out_a77) ,.jpeg_out_a78(jpeg_out_a78) ,
	.jpeg_out_a79(jpeg_out_a79) ,.jpeg_out_a80(jpeg_out_a80) ,.jpeg_out_a81(jpeg_out_a81) ,
	.jpeg_out_a82(jpeg_out_a82) ,.jpeg_out_a83(jpeg_out_a83) ,.jpeg_out_a84(jpeg_out_a84) ,
	.jpeg_out_a85(jpeg_out_a85) ,.jpeg_out_a86(jpeg_out_a86) ,.jpeg_out_a87(jpeg_out_a87) ,
	.jpeg_out_a88(jpeg_out_a88) ,.jpeg_out_a89(jpeg_out_a89) ,.jpeg_out_a90(jpeg_out_a90) ,
	.jpeg_out_a91(jpeg_out_a91) ,.jpeg_out_a92(jpeg_out_a92) ,.jpeg_out_a93(jpeg_out_a93) ,
	.jpeg_out_a94(jpeg_out_a94) ,.jpeg_out_a95(jpeg_out_a95) ,.jpeg_out_a96(jpeg_out_a96) ,
	.jpeg_out_a97(jpeg_out_a97) ,.jpeg_out_a98(jpeg_out_a98) ,.jpeg_out_a99(jpeg_out_a99) ,
	.jpeg_out_a100(jpeg_out_a100) ,.jpeg_out_a101(jpeg_out_a101) ,.jpeg_out_a102(jpeg_out_a102) ,
	.jpeg_out_a103(jpeg_out_a103) ,.jpeg_out_a104(jpeg_out_a104) ,.jpeg_out_a105(jpeg_out_a105) ,
	.jpeg_out_a106(jpeg_out_a106) ,.jpeg_out_a107(jpeg_out_a107) ,.jpeg_out_a108(jpeg_out_a108) ,
	.jpeg_out_a109(jpeg_out_a109) ,.jpeg_out_a110(jpeg_out_a110) ,.jpeg_out_a111(jpeg_out_a111) ,
	.jpeg_out_a112(jpeg_out_a112) ,.jpeg_out_a113(jpeg_out_a113) ,.jpeg_out_a114(jpeg_out_a114) ,
	.jpeg_out_a115(jpeg_out_a115) ,.jpeg_out_a116(jpeg_out_a116) ,.jpeg_out_a117(jpeg_out_a117) ,
	.jpeg_out_a118(jpeg_out_a118) ,.jpeg_out_a119(jpeg_out_a119) ,.jpeg_out_a120(jpeg_out_a120) ,
	.jpeg_out_a121(jpeg_out_a121) ,.jpeg_out_a122(jpeg_out_a122) ,.jpeg_out_a123(jpeg_out_a123) ,
	.jpeg_out_a124(jpeg_out_a124) ,.jpeg_out_a125(jpeg_out_a125) ,.jpeg_out_a126(jpeg_out_a126) ,
	.jpeg_out_a127(jpeg_out_a127) ,.jpeg_len_out(jpeg_len_out) ,.valid(valid) ,
	.ST1_11d(ST1_11d) ,.ST1_10d(ST1_10d) ,.ST1_09d(ST1_09d) ,.ST1_08d(ST1_08d) ,
	.ST1_07d(ST1_07d) ,.ST1_06d(ST1_06d) ,.ST1_05d(ST1_05d) ,.ST1_04d(ST1_04d) ,
	.ST1_03d(ST1_03d) ,.ST1_02d(ST1_02d) ,.ST1_01d(ST1_01d) ,.JF_01(JF_01) ,
	.lop8u_11ot_port(lop8u_11ot) ,.JF_03(JF_03) ,.CT_33_port(CT_33) ,.RG_315_port(RG_315) ,
	.JF_06(JF_06) );

endmodule

module jpeg_fsm ( clk ,rst ,ST1_11d ,ST1_10d ,ST1_09d ,ST1_08d ,ST1_07d ,ST1_06d ,
	ST1_05d ,ST1_04d ,ST1_03d ,ST1_02d ,ST1_01d ,JF_01 ,lop8u_11ot ,JF_03 ,CT_33 ,
	RG_315 ,JF_06 );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
output		ST1_11d ;
output		ST1_10d ;
output		ST1_09d ;
output		ST1_08d ;
output		ST1_07d ;
output		ST1_06d ;
output		ST1_05d ;
output		ST1_04d ;
output		ST1_03d ;
output		ST1_02d ;
output		ST1_01d ;
input		JF_01 ;
input		lop8u_11ot ;
input		JF_03 ;
input		CT_33 ;
input		RG_315 ;
input		JF_06 ;
reg	[3:0]	B01_streg ;

parameter	ST1_01 = 4'h0 ;
parameter	ST1_02 = 4'h1 ;
parameter	ST1_03 = 4'h2 ;
parameter	ST1_04 = 4'h3 ;
parameter	ST1_05 = 4'h4 ;
parameter	ST1_06 = 4'h5 ;
parameter	ST1_07 = 4'h6 ;
parameter	ST1_08 = 4'h7 ;
parameter	ST1_09 = 4'h8 ;
parameter	ST1_10 = 4'h9 ;
parameter	ST1_11 = 4'ha ;

assign	ST1_01d = ( ( B01_streg == ST1_01 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_02d = ( ( B01_streg == ST1_02 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_03d = ( ( B01_streg == ST1_03 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_04d = ( ( B01_streg == ST1_04 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_05d = ( ( B01_streg == ST1_05 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_06d = ( ( B01_streg == ST1_06 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_07d = ( ( B01_streg == ST1_07 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_08d = ( ( B01_streg == ST1_08 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_09d = ( ( B01_streg == ST1_09 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_10d = ( ( B01_streg == ST1_10 ) ? 1'h1 : 1'h0 ) ;
assign	ST1_11d = ( ( B01_streg == ST1_11 ) ? 1'h1 : 1'h0 ) ;
always @ ( posedge clk )
	if ( !rst )
		B01_streg <= ST1_01 ;
	else
		case ( B01_streg )
		ST1_01 :
			B01_streg <= ST1_02 ;
		ST1_02 :
			if ( ( JF_01 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_03 ;
		ST1_03 :
			if ( ( lop8u_11ot != 1'h0 ) )
				B01_streg <= ST1_03 ;
			else
				B01_streg <= ST1_04 ;
		ST1_04 :
			if ( ( JF_03 != 1'h0 ) )
				B01_streg <= ST1_04 ;
			else
				B01_streg <= ST1_05 ;
		ST1_05 :
			B01_streg <= ST1_06 ;
		ST1_06 :
			B01_streg <= ST1_07 ;
		ST1_07 :
			B01_streg <= ST1_08 ;
		ST1_08 :
			if ( ( CT_33 != 1'h0 ) )
				B01_streg <= ST1_07 ;
			else
				B01_streg <= ST1_09 ;
		ST1_09 :
			if ( ( RG_315 != 1'h0 ) )
				B01_streg <= ST1_07 ;
			else
				B01_streg <= ST1_10 ;
		ST1_10 :
			B01_streg <= ST1_11 ;
		ST1_11 :
			if ( ( JF_06 != 1'h0 ) )
				B01_streg <= ST1_02 ;
			else
				B01_streg <= ST1_11 ;
		default :
			B01_streg <= ST1_01 ;
		endcase

endmodule

module jpeg_dat ( clk ,rst ,jpeg_in_a00 ,jpeg_in_a01 ,jpeg_in_a02 ,jpeg_in_a03 ,
	jpeg_in_a04 ,jpeg_in_a05 ,jpeg_in_a06 ,jpeg_in_a07 ,jpeg_in_a08 ,jpeg_in_a09 ,
	jpeg_in_a10 ,jpeg_in_a11 ,jpeg_in_a12 ,jpeg_in_a13 ,jpeg_in_a14 ,jpeg_in_a15 ,
	jpeg_in_a16 ,jpeg_in_a17 ,jpeg_in_a18 ,jpeg_in_a19 ,jpeg_in_a20 ,jpeg_in_a21 ,
	jpeg_in_a22 ,jpeg_in_a23 ,jpeg_in_a24 ,jpeg_in_a25 ,jpeg_in_a26 ,jpeg_in_a27 ,
	jpeg_in_a28 ,jpeg_in_a29 ,jpeg_in_a30 ,jpeg_in_a31 ,jpeg_in_a32 ,jpeg_in_a33 ,
	jpeg_in_a34 ,jpeg_in_a35 ,jpeg_in_a36 ,jpeg_in_a37 ,jpeg_in_a38 ,jpeg_in_a39 ,
	jpeg_in_a40 ,jpeg_in_a41 ,jpeg_in_a42 ,jpeg_in_a43 ,jpeg_in_a44 ,jpeg_in_a45 ,
	jpeg_in_a46 ,jpeg_in_a47 ,jpeg_in_a48 ,jpeg_in_a49 ,jpeg_in_a50 ,jpeg_in_a51 ,
	jpeg_in_a52 ,jpeg_in_a53 ,jpeg_in_a54 ,jpeg_in_a55 ,jpeg_in_a56 ,jpeg_in_a57 ,
	jpeg_in_a58 ,jpeg_in_a59 ,jpeg_in_a60 ,jpeg_in_a61 ,jpeg_in_a62 ,jpeg_in_a63 ,
	jpeg_out_a00 ,jpeg_out_a01 ,jpeg_out_a02 ,jpeg_out_a03 ,jpeg_out_a04 ,jpeg_out_a05 ,
	jpeg_out_a06 ,jpeg_out_a07 ,jpeg_out_a08 ,jpeg_out_a09 ,jpeg_out_a10 ,jpeg_out_a11 ,
	jpeg_out_a12 ,jpeg_out_a13 ,jpeg_out_a14 ,jpeg_out_a15 ,jpeg_out_a16 ,jpeg_out_a17 ,
	jpeg_out_a18 ,jpeg_out_a19 ,jpeg_out_a20 ,jpeg_out_a21 ,jpeg_out_a22 ,jpeg_out_a23 ,
	jpeg_out_a24 ,jpeg_out_a25 ,jpeg_out_a26 ,jpeg_out_a27 ,jpeg_out_a28 ,jpeg_out_a29 ,
	jpeg_out_a30 ,jpeg_out_a31 ,jpeg_out_a32 ,jpeg_out_a33 ,jpeg_out_a34 ,jpeg_out_a35 ,
	jpeg_out_a36 ,jpeg_out_a37 ,jpeg_out_a38 ,jpeg_out_a39 ,jpeg_out_a40 ,jpeg_out_a41 ,
	jpeg_out_a42 ,jpeg_out_a43 ,jpeg_out_a44 ,jpeg_out_a45 ,jpeg_out_a46 ,jpeg_out_a47 ,
	jpeg_out_a48 ,jpeg_out_a49 ,jpeg_out_a50 ,jpeg_out_a51 ,jpeg_out_a52 ,jpeg_out_a53 ,
	jpeg_out_a54 ,jpeg_out_a55 ,jpeg_out_a56 ,jpeg_out_a57 ,jpeg_out_a58 ,jpeg_out_a59 ,
	jpeg_out_a60 ,jpeg_out_a61 ,jpeg_out_a62 ,jpeg_out_a63 ,jpeg_out_a64 ,jpeg_out_a65 ,
	jpeg_out_a66 ,jpeg_out_a67 ,jpeg_out_a68 ,jpeg_out_a69 ,jpeg_out_a70 ,jpeg_out_a71 ,
	jpeg_out_a72 ,jpeg_out_a73 ,jpeg_out_a74 ,jpeg_out_a75 ,jpeg_out_a76 ,jpeg_out_a77 ,
	jpeg_out_a78 ,jpeg_out_a79 ,jpeg_out_a80 ,jpeg_out_a81 ,jpeg_out_a82 ,jpeg_out_a83 ,
	jpeg_out_a84 ,jpeg_out_a85 ,jpeg_out_a86 ,jpeg_out_a87 ,jpeg_out_a88 ,jpeg_out_a89 ,
	jpeg_out_a90 ,jpeg_out_a91 ,jpeg_out_a92 ,jpeg_out_a93 ,jpeg_out_a94 ,jpeg_out_a95 ,
	jpeg_out_a96 ,jpeg_out_a97 ,jpeg_out_a98 ,jpeg_out_a99 ,jpeg_out_a100 ,jpeg_out_a101 ,
	jpeg_out_a102 ,jpeg_out_a103 ,jpeg_out_a104 ,jpeg_out_a105 ,jpeg_out_a106 ,
	jpeg_out_a107 ,jpeg_out_a108 ,jpeg_out_a109 ,jpeg_out_a110 ,jpeg_out_a111 ,
	jpeg_out_a112 ,jpeg_out_a113 ,jpeg_out_a114 ,jpeg_out_a115 ,jpeg_out_a116 ,
	jpeg_out_a117 ,jpeg_out_a118 ,jpeg_out_a119 ,jpeg_out_a120 ,jpeg_out_a121 ,
	jpeg_out_a122 ,jpeg_out_a123 ,jpeg_out_a124 ,jpeg_out_a125 ,jpeg_out_a126 ,
	jpeg_out_a127 ,jpeg_len_out ,valid ,ST1_11d ,ST1_10d ,ST1_09d ,ST1_08d ,
	ST1_07d ,ST1_06d ,ST1_05d ,ST1_04d ,ST1_03d ,ST1_02d ,ST1_01d ,JF_01 ,lop8u_11ot_port ,
	JF_03 ,CT_33_port ,RG_315_port ,JF_06 );
input		clk ;	// line#=../rle.h:52
input		rst ;	// line#=../rle.h:53
input	[8:0]	jpeg_in_a00 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a01 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a02 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a03 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a04 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a05 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a06 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a07 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a08 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a09 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a10 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a11 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a12 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a13 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a14 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a15 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a16 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a17 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a18 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a19 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a20 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a21 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a22 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a23 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a24 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a25 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a26 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a27 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a28 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a29 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a30 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a31 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a32 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a33 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a34 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a35 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a36 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a37 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a38 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a39 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a40 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a41 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a42 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a43 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a44 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a45 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a46 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a47 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a48 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a49 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a50 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a51 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a52 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a53 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a54 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a55 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a56 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a57 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a58 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a59 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a60 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a61 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a62 ;	// line#=../rle.h:56
input	[8:0]	jpeg_in_a63 ;	// line#=../rle.h:56
output	[8:0]	jpeg_out_a00 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a01 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a02 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a03 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a04 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a05 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a06 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a07 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a08 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a09 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a10 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a11 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a12 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a13 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a14 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a15 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a16 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a17 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a18 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a19 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a20 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a21 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a22 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a23 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a24 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a25 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a26 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a27 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a28 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a29 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a30 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a31 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a32 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a33 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a34 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a35 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a36 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a37 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a38 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a39 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a40 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a41 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a42 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a43 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a44 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a45 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a46 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a47 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a48 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a49 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a50 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a51 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a52 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a53 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a54 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a55 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a56 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a57 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a58 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a59 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a60 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a61 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a62 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a63 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a64 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a65 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a66 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a67 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a68 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a69 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a70 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a71 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a72 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a73 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a74 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a75 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a76 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a77 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a78 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a79 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a80 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a81 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a82 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a83 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a84 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a85 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a86 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a87 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a88 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a89 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a90 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a91 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a92 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a93 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a94 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a95 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a96 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a97 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a98 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a99 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a100 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a101 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a102 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a103 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a104 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a105 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a106 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a107 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a108 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a109 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a110 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a111 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a112 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a113 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a114 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a115 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a116 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a117 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a118 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a119 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a120 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a121 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a122 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a123 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a124 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a125 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a126 ;	// line#=../rle.h:60
output	[8:0]	jpeg_out_a127 ;	// line#=../rle.h:60
output	[11:0]	jpeg_len_out ;	// line#=../rle.h:61
output		valid ;	// line#=../rle.h:62
input		ST1_11d ;
input		ST1_10d ;
input		ST1_09d ;
input		ST1_08d ;
input		ST1_07d ;
input		ST1_06d ;
input		ST1_05d ;
input		ST1_04d ;
input		ST1_03d ;
input		ST1_02d ;
input		ST1_01d ;
output		JF_01 ;
output		lop8u_11ot_port ;
output		JF_03 ;
output		CT_33_port ;
output		RG_315_port ;
output		JF_06 ;
wire		M_321 ;
wire		M_320 ;
wire		M_319 ;
wire		M_318 ;
wire		M_317 ;
wire		M_316 ;
wire		M_315 ;
wire		M_314 ;
wire		M_313 ;
wire		M_312 ;
wire		M_311 ;
wire		M_310 ;
wire		M_309 ;
wire		M_308 ;
wire		M_307 ;
wire		M_306 ;
wire		M_305 ;
wire		M_304 ;
wire		M_303 ;
wire		M_302 ;
wire		M_301 ;
wire		M_300 ;
wire		M_299 ;
wire		M_298 ;
wire		M_297 ;
wire		M_296 ;
wire		M_295 ;
wire		M_294 ;
wire		M_293 ;
wire		M_292 ;
wire		M_291 ;
wire		M_290 ;
wire		M_289 ;
wire		M_288 ;
wire		M_287 ;
wire		M_286 ;
wire		M_285 ;
wire		M_284 ;
wire		M_283 ;
wire		M_282 ;
wire		M_281 ;
wire		M_280 ;
wire		M_279 ;
wire		M_278 ;
wire		M_277 ;
wire		M_276 ;
wire		M_275 ;
wire		M_274 ;
wire		M_273 ;
wire		M_272 ;
wire		M_271 ;
wire		M_270 ;
wire		M_269 ;
wire		M_268 ;
wire		M_267 ;
wire		M_266 ;
wire		M_265 ;
wire		M_264 ;
wire		M_263 ;
wire		M_262 ;
wire		M_261 ;
wire		M_260 ;
wire		M_259 ;
wire		M_258 ;
wire		M_257 ;
wire		M_256 ;
wire		M_255 ;
wire		M_254 ;
wire		M_253 ;
wire		M_252 ;
wire		M_251 ;
wire		M_250 ;
wire		M_249 ;
wire		M_248 ;
wire		M_247 ;
wire		M_246 ;
wire		M_245 ;
wire		M_244 ;
wire		M_243 ;
wire		M_242 ;
wire		M_241 ;
wire		M_240 ;
wire		M_239 ;
wire		M_238 ;
wire		M_237 ;
wire		M_236 ;
wire		M_235 ;
wire		M_234 ;
wire		M_233 ;
wire		M_232 ;
wire		M_231 ;
wire		M_230 ;
wire		M_229 ;
wire		M_228 ;
wire		M_227 ;
wire		M_226 ;
wire		M_225 ;
wire		M_224 ;
wire		M_223 ;
wire		M_222 ;
wire		M_221 ;
wire		M_220 ;
wire		M_219 ;
wire		M_218 ;
wire		M_217 ;
wire		M_216 ;
wire		M_215 ;
wire		M_214 ;
wire		M_213 ;
wire		M_212 ;
wire		M_211 ;
wire		M_210 ;
wire		M_209 ;
wire		M_208 ;
wire		M_207 ;
wire		M_206 ;
wire		M_205 ;
wire		M_204 ;
wire		M_203 ;
wire		M_202 ;
wire		M_201 ;
wire		M_200 ;
wire		M_199 ;
wire		M_198 ;
wire		M_197 ;
wire		M_196 ;
wire		M_195 ;
wire		M_194 ;
wire		M_193 ;
wire		M_192 ;
wire		M_191 ;
wire		M_190 ;
wire		M_189 ;
wire		M_188 ;
wire		M_187 ;
wire		M_186 ;
wire		M_185 ;
wire		M_184 ;
wire		M_183 ;
wire		M_182 ;
wire		M_181 ;
wire		M_180 ;
wire		M_179 ;
wire		M_178 ;
wire		M_177 ;
wire		M_176 ;
wire		M_175 ;
wire		M_174 ;
wire		M_173 ;
wire		M_172 ;
wire		U_572 ;
wire		U_571 ;
wire		U_570 ;
wire		U_569 ;
wire		U_174 ;
wire		U_173 ;
wire		U_172 ;
wire		U_171 ;
wire		U_166 ;
wire		U_165 ;
wire		U_164 ;
wire		U_163 ;
wire		U_162 ;
wire		C_05 ;
wire		U_161 ;
wire		U_96 ;
wire		U_95 ;
wire		U_94 ;
wire		U_93 ;
wire		U_92 ;
wire		U_91 ;
wire		U_90 ;
wire		U_89 ;
wire		U_88 ;
wire		U_87 ;
wire		U_84 ;
wire		U_83 ;
wire		U_82 ;
wire		U_81 ;
wire		U_80 ;
wire		C_02 ;
wire		U_79 ;
wire		U_14 ;
wire		U_13 ;
wire		U_12 ;
wire		U_11 ;
wire		U_10 ;
wire		U_09 ;
wire		U_08 ;
wire		U_07 ;
wire		U_06 ;
wire		U_05 ;
wire		C_01 ;
wire		U_01 ;
wire	[1:0]	sub8u_7_11i2 ;
wire	[6:0]	sub8u_7_11i1 ;
wire	[6:0]	sub8u_7_11ot ;
wire	[2:0]	sub8u_71i2 ;
wire	[6:0]	sub8u_71i1 ;
wire	[6:0]	sub8u_71ot ;
wire	[31:0]	decr32s2i1 ;
wire	[31:0]	decr32s2ot ;
wire	[31:0]	decr32s1i1 ;
wire	[31:0]	decr32s1ot ;
wire	[6:0]	decr8u_71i1 ;
wire	[6:0]	decr8u_71ot ;
wire	[31:0]	incr32s3i1 ;
wire	[31:0]	incr32s3ot ;
wire	[31:0]	incr32s2i1 ;
wire	[31:0]	incr32s2ot ;
wire	[31:0]	incr32s1i1 ;
wire	[31:0]	incr32s1ot ;
wire	[7:0]	incr8u4i1 ;
wire	[7:0]	incr8u4ot ;
wire	[7:0]	incr8u3ot ;
wire	[7:0]	incr8u2i1 ;
wire	[7:0]	incr8u2ot ;
wire	[7:0]	incr8u1i1 ;
wire	[7:0]	incr8u1ot ;
wire	[3:0]	incr4s1i1 ;
wire	[3:0]	incr4s1ot ;
wire	[5:0]	lop8u_11i2 ;
wire	[5:0]	lop8u_11i1 ;
wire		lop8u_11ot ;
wire	[8:0]	sub12s_91i2 ;
wire	[8:0]	sub12s_91i1 ;
wire	[8:0]	sub12s_91ot ;
wire	[1:0]	sub8u1i2 ;
wire	[7:0]	sub8u1ot ;
wire		JF_06 ;
wire		CT_33 ;
wire		CT_32 ;
wire		CT_28 ;
wire		CT_17 ;
wire		JF_03 ;
wire		CT_12 ;
wire		JF_01 ;
wire		zz_WE2 ;
wire	[8:0]	zz_RD1 ;
wire		RG_previous_dc_en ;
wire		RG_rl_128_en ;
wire		RG_rl_129_en ;
wire		RG_rl_130_en ;
wire		RG_rl_131_en ;
wire		RG_rl_132_en ;
wire		RG_rl_133_en ;
wire		RG_rl_134_en ;
wire		RG_rl_135_en ;
wire		RG_rl_136_en ;
wire		RG_rl_137_en ;
wire		RG_rl_138_en ;
wire		RG_rl_139_en ;
wire		RG_rl_140_en ;
wire		RG_rl_141_en ;
wire		RG_rl_142_en ;
wire		RG_rl_143_en ;
wire		RG_rl_144_en ;
wire		RG_rl_145_en ;
wire		RG_rl_146_en ;
wire		RG_rl_147_en ;
wire		RG_rl_148_en ;
wire		RG_rl_149_en ;
wire		RG_rl_150_en ;
wire		RG_rl_151_en ;
wire		RG_rl_152_en ;
wire		RG_rl_153_en ;
wire		RG_rl_154_en ;
wire		RG_rl_155_en ;
wire		RG_rl_156_en ;
wire		RG_rl_157_en ;
wire		RG_rl_158_en ;
wire		RG_rl_159_en ;
wire		RG_rl_160_en ;
wire		RG_rl_161_en ;
wire		RG_rl_162_en ;
wire		RG_rl_163_en ;
wire		RG_rl_164_en ;
wire		RG_rl_165_en ;
wire		RG_rl_166_en ;
wire		RG_rl_167_en ;
wire		RG_rl_168_en ;
wire		RG_rl_169_en ;
wire		RG_rl_170_en ;
wire		RG_rl_171_en ;
wire		RG_rl_172_en ;
wire		RG_rl_173_en ;
wire		RG_rl_174_en ;
wire		RG_rl_175_en ;
wire		RG_rl_176_en ;
wire		RG_rl_177_en ;
wire		RG_rl_178_en ;
wire		RG_rl_179_en ;
wire		RG_rl_180_en ;
wire		RG_rl_181_en ;
wire		RG_rl_182_en ;
wire		RG_rl_183_en ;
wire		FF_j_en ;
wire		RG_315_en ;
wire		RG_len_01_en ;
wire		jpeg_out_a00_r_en ;
wire		jpeg_out_a01_r_en ;
wire		jpeg_out_a02_r_en ;
wire		jpeg_out_a03_r_en ;
wire		jpeg_out_a04_r_en ;
wire		jpeg_out_a05_r_en ;
wire		jpeg_out_a06_r_en ;
wire		jpeg_out_a07_r_en ;
wire		jpeg_out_a08_r_en ;
wire		jpeg_out_a09_r_en ;
wire		jpeg_out_a10_r_en ;
wire		jpeg_out_a11_r_en ;
wire		jpeg_out_a12_r_en ;
wire		jpeg_out_a13_r_en ;
wire		jpeg_out_a14_r_en ;
wire		jpeg_out_a15_r_en ;
wire		jpeg_out_a16_r_en ;
wire		jpeg_out_a17_r_en ;
wire		jpeg_out_a18_r_en ;
wire		jpeg_out_a19_r_en ;
wire		jpeg_out_a20_r_en ;
wire		jpeg_out_a21_r_en ;
wire		jpeg_out_a22_r_en ;
wire		jpeg_out_a23_r_en ;
wire		jpeg_out_a24_r_en ;
wire		jpeg_out_a25_r_en ;
wire		jpeg_out_a26_r_en ;
wire		jpeg_out_a27_r_en ;
wire		jpeg_out_a28_r_en ;
wire		jpeg_out_a29_r_en ;
wire		jpeg_out_a30_r_en ;
wire		jpeg_out_a31_r_en ;
wire		jpeg_out_a32_r_en ;
wire		jpeg_out_a33_r_en ;
wire		jpeg_out_a34_r_en ;
wire		jpeg_out_a35_r_en ;
wire		jpeg_out_a36_r_en ;
wire		jpeg_out_a37_r_en ;
wire		jpeg_out_a38_r_en ;
wire		jpeg_out_a39_r_en ;
wire		jpeg_out_a40_r_en ;
wire		jpeg_out_a41_r_en ;
wire		jpeg_out_a42_r_en ;
wire		jpeg_out_a43_r_en ;
wire		jpeg_out_a44_r_en ;
wire		jpeg_out_a45_r_en ;
wire		jpeg_out_a46_r_en ;
wire		jpeg_out_a47_r_en ;
wire		jpeg_out_a48_r_en ;
wire		jpeg_out_a49_r_en ;
wire		jpeg_out_a50_r_en ;
wire		jpeg_out_a51_r_en ;
wire		jpeg_out_a52_r_en ;
wire		jpeg_out_a53_r_en ;
wire		jpeg_out_a54_r_en ;
wire		jpeg_out_a55_r_en ;
wire		jpeg_out_a56_r_en ;
wire		jpeg_out_a57_r_en ;
wire		jpeg_out_a58_r_en ;
wire		jpeg_out_a59_r_en ;
wire		jpeg_out_a60_r_en ;
wire		jpeg_out_a61_r_en ;
wire		jpeg_out_a62_r_en ;
wire		jpeg_out_a63_r_en ;
wire		jpeg_out_a64_r_en ;
wire		jpeg_out_a65_r_en ;
wire		jpeg_out_a66_r_en ;
wire		jpeg_out_a67_r_en ;
wire		jpeg_out_a68_r_en ;
wire		jpeg_out_a69_r_en ;
wire		jpeg_out_a70_r_en ;
wire		jpeg_out_a71_r_en ;
wire		jpeg_out_a72_r_en ;
wire		jpeg_out_a73_r_en ;
wire		jpeg_out_a74_r_en ;
wire		jpeg_out_a75_r_en ;
wire		jpeg_out_a76_r_en ;
wire		jpeg_out_a77_r_en ;
wire		jpeg_out_a78_r_en ;
wire		jpeg_out_a79_r_en ;
wire		jpeg_out_a80_r_en ;
wire		jpeg_out_a81_r_en ;
wire		jpeg_out_a82_r_en ;
wire		jpeg_out_a83_r_en ;
wire		jpeg_out_a84_r_en ;
wire		jpeg_out_a85_r_en ;
wire		jpeg_out_a86_r_en ;
wire		jpeg_out_a87_r_en ;
wire		jpeg_out_a88_r_en ;
wire		jpeg_out_a89_r_en ;
wire		jpeg_out_a90_r_en ;
wire		jpeg_out_a91_r_en ;
wire		jpeg_out_a92_r_en ;
wire		jpeg_out_a93_r_en ;
wire		jpeg_out_a94_r_en ;
wire		jpeg_out_a95_r_en ;
wire		jpeg_out_a96_r_en ;
wire		jpeg_out_a97_r_en ;
wire		jpeg_out_a98_r_en ;
wire		jpeg_out_a99_r_en ;
wire		jpeg_out_a100_r_en ;
wire		jpeg_out_a101_r_en ;
wire		jpeg_out_a102_r_en ;
wire		jpeg_out_a103_r_en ;
wire		jpeg_out_a104_r_en ;
wire		jpeg_out_a105_r_en ;
wire		jpeg_out_a106_r_en ;
wire		jpeg_out_a107_r_en ;
wire		jpeg_out_a108_r_en ;
wire		jpeg_out_a109_r_en ;
wire		jpeg_out_a110_r_en ;
wire		jpeg_out_a111_r_en ;
wire		jpeg_out_a112_r_en ;
wire		jpeg_out_a113_r_en ;
wire		jpeg_out_a114_r_en ;
wire		jpeg_out_a115_r_en ;
wire		jpeg_out_a116_r_en ;
wire		jpeg_out_a117_r_en ;
wire		jpeg_out_a118_r_en ;
wire		jpeg_out_a119_r_en ;
wire		jpeg_out_a120_r_en ;
wire		jpeg_out_a121_r_en ;
wire		jpeg_out_a122_r_en ;
wire		jpeg_out_a123_r_en ;
wire		jpeg_out_a124_r_en ;
wire		jpeg_out_a125_r_en ;
wire		jpeg_out_a126_r_en ;
wire		jpeg_out_a127_r_en ;
wire		jpeg_len_out_r_en ;
wire		RG_rl_en ;
wire		RG_rl_1_en ;
wire		RG_rl_2_en ;
wire		RG_rl_3_en ;
wire		RG_rl_4_en ;
wire		RG_rl_5_en ;
wire		RG_rl_6_en ;
wire		RG_rl_7_en ;
wire		RG_rl_8_en ;
wire		RG_rl_9_en ;
wire		RG_rl_10_en ;
wire		RG_rl_11_en ;
wire		RG_rl_12_en ;
wire		RG_rl_13_en ;
wire		RG_rl_14_en ;
wire		RG_rl_15_en ;
wire		RG_rl_16_en ;
wire		RG_rl_17_en ;
wire		RG_rl_18_en ;
wire		RG_rl_19_en ;
wire		RG_rl_20_en ;
wire		RG_rl_21_en ;
wire		RG_rl_22_en ;
wire		RG_rl_23_en ;
wire		RG_rl_24_en ;
wire		RG_rl_25_en ;
wire		RG_rl_26_en ;
wire		RG_rl_27_en ;
wire		RG_rl_28_en ;
wire		RG_rl_29_en ;
wire		RG_rl_30_en ;
wire		RG_rl_31_en ;
wire		RG_rl_32_en ;
wire		RG_rl_33_en ;
wire		RG_rl_34_en ;
wire		RG_rl_35_en ;
wire		RG_rl_36_en ;
wire		RG_rl_37_en ;
wire		RG_rl_38_en ;
wire		RG_rl_39_en ;
wire		RG_rl_40_en ;
wire		RG_rl_41_en ;
wire		RG_rl_42_en ;
wire		RG_rl_43_en ;
wire		RG_rl_44_en ;
wire		RG_rl_45_en ;
wire		RG_rl_46_en ;
wire		RG_rl_47_en ;
wire		RG_rl_48_en ;
wire		RG_rl_49_en ;
wire		RG_rl_50_en ;
wire		RG_rl_51_en ;
wire		RG_rl_52_en ;
wire		RG_rl_53_en ;
wire		RG_rl_54_en ;
wire		RG_rl_55_en ;
wire		RG_rl_56_en ;
wire		RG_rl_57_en ;
wire		RG_rl_58_en ;
wire		RG_rl_59_en ;
wire		RG_rl_60_en ;
wire		RG_rl_61_en ;
wire		RG_rl_62_en ;
wire		RG_rl_63_en ;
wire		RG_rl_64_en ;
wire		RG_rl_65_en ;
wire		RG_rl_66_en ;
wire		RG_rl_67_en ;
wire		RG_rl_68_en ;
wire		RG_rl_69_en ;
wire		RG_rl_70_en ;
wire		RG_rl_71_en ;
wire		RG_rl_72_en ;
wire		RG_rl_73_en ;
wire		RG_rl_74_en ;
wire		RG_rl_75_en ;
wire		RG_rl_76_en ;
wire		RG_rl_77_en ;
wire		RG_rl_78_en ;
wire		RG_rl_79_en ;
wire		RG_rl_80_en ;
wire		RG_rl_81_en ;
wire		RG_rl_82_en ;
wire		RG_rl_83_en ;
wire		RG_rl_84_en ;
wire		RG_rl_85_en ;
wire		RG_rl_86_en ;
wire		RG_rl_87_en ;
wire		RG_rl_88_en ;
wire		RG_rl_89_en ;
wire		RG_rl_90_en ;
wire		RG_rl_91_en ;
wire		RG_rl_92_en ;
wire		RG_rl_93_en ;
wire		RG_rl_94_en ;
wire		RG_rl_95_en ;
wire		RG_rl_96_en ;
wire		RG_rl_97_en ;
wire		RG_rl_98_en ;
wire		RG_rl_99_en ;
wire		RG_rl_100_en ;
wire		RG_rl_101_en ;
wire		RG_rl_102_en ;
wire		RG_rl_103_en ;
wire		RG_rl_104_en ;
wire		RG_rl_105_en ;
wire		RG_rl_106_en ;
wire		RG_rl_107_en ;
wire		RG_rl_108_en ;
wire		RG_rl_109_en ;
wire		RG_rl_110_en ;
wire		RG_rl_111_en ;
wire		RG_rl_112_en ;
wire		RG_rl_113_en ;
wire		RG_rl_114_en ;
wire		RG_rl_115_en ;
wire		RG_rl_116_en ;
wire		RG_rl_117_en ;
wire		RG_rl_118_en ;
wire		RG_rl_119_en ;
wire		RG_rl_120_en ;
wire		RG_rl_121_en ;
wire		RG_rl_122_en ;
wire		RG_rl_123_en ;
wire		RG_rl_124_en ;
wire		RG_rl_125_en ;
wire		RG_rl_126_en ;
wire		RG_rl_127_en ;
wire		RG_rl_184_en ;
wire		RG_previous_dc_rl_en ;
wire		RG_rl_185_en ;
wire		RG_rl_186_en ;
wire		RG_rl_187_en ;
wire		RG_rl_188_en ;
wire		RG_rl_189_en ;
wire		RG_rl_190_en ;
wire		RG_rl_191_en ;
wire		RG_rl_192_en ;
wire		RG_rl_193_en ;
wire		RG_rl_194_en ;
wire		RG_rl_195_en ;
wire		RG_rl_196_en ;
wire		RG_rl_197_en ;
wire		RG_rl_198_en ;
wire		RG_rl_199_en ;
wire		RG_rl_200_en ;
wire		RG_rl_201_en ;
wire		RG_rl_202_en ;
wire		RG_rl_203_en ;
wire		RG_rl_204_en ;
wire		RG_rl_205_en ;
wire		RG_rl_206_en ;
wire		RG_rl_207_en ;
wire		RG_rl_208_en ;
wire		RG_rl_209_en ;
wire		RG_rl_210_en ;
wire		RG_rl_211_en ;
wire		RG_rl_212_en ;
wire		RG_rl_213_en ;
wire		RG_rl_214_en ;
wire		RG_rl_215_en ;
wire		RG_rl_216_en ;
wire		RG_rl_217_en ;
wire		RG_rl_218_en ;
wire		RG_rl_219_en ;
wire		RG_rl_220_en ;
wire		RG_rl_221_en ;
wire		RG_rl_222_en ;
wire		RG_rl_223_en ;
wire		RG_rl_224_en ;
wire		RG_rl_225_en ;
wire		RG_rl_226_en ;
wire		RG_rl_227_en ;
wire		RG_rl_228_en ;
wire		RG_rl_229_en ;
wire		RG_rl_230_en ;
wire		RG_rl_231_en ;
wire		RG_rl_232_en ;
wire		RG_rl_233_en ;
wire		RG_rl_234_en ;
wire		RG_rl_235_en ;
wire		RG_rl_236_en ;
wire		RG_rl_237_en ;
wire		RG_rl_238_en ;
wire		RG_rl_239_en ;
wire		RG_rl_240_en ;
wire		RG_rl_241_en ;
wire		RG_i_k_01_en ;
wire		RG_i_j_01_en ;
wire		RG_quantized_block_rl_en ;
wire		RG_quantized_block_rl_1_en ;
wire		RG_quantized_block_rl_2_en ;
wire		RG_quantized_block_rl_3_en ;
wire		RG_quantized_block_rl_4_en ;
wire		RG_quantized_block_rl_5_en ;
wire		RG_quantized_block_rl_6_en ;
wire		RG_quantized_block_rl_7_en ;
wire		RG_quantized_block_rl_8_en ;
wire		RG_quantized_block_rl_9_en ;
wire		RG_quantized_block_rl_10_en ;
wire		RG_quantized_block_rl_11_en ;
wire		RG_quantized_block_rl_12_en ;
wire		RG_quantized_block_rl_13_en ;
wire		RG_quantized_block_rl_14_en ;
wire		RG_quantized_block_rl_15_en ;
wire		RG_quantized_block_rl_16_en ;
wire		RG_quantized_block_rl_17_en ;
wire		RG_quantized_block_rl_18_en ;
wire		RG_quantized_block_rl_19_en ;
wire		RG_quantized_block_rl_20_en ;
wire		RG_quantized_block_rl_21_en ;
wire		RG_quantized_block_rl_22_en ;
wire		RG_quantized_block_rl_23_en ;
wire		RG_quantized_block_rl_24_en ;
wire		RG_quantized_block_rl_25_en ;
wire		RG_quantized_block_rl_26_en ;
wire		RG_quantized_block_rl_27_en ;
wire		RG_quantized_block_rl_28_en ;
wire		RG_quantized_block_rl_29_en ;
wire		RG_quantized_block_rl_30_en ;
wire		RG_quantized_block_rl_31_en ;
wire		RG_quantized_block_rl_32_en ;
wire		RG_quantized_block_rl_33_en ;
wire		RG_quantized_block_rl_34_en ;
wire		RG_quantized_block_rl_35_en ;
wire		RG_quantized_block_rl_36_en ;
wire		RG_quantized_block_rl_37_en ;
wire		RG_quantized_block_rl_38_en ;
wire		RG_quantized_block_rl_39_en ;
wire		RG_quantized_block_rl_40_en ;
wire		RG_quantized_block_rl_41_en ;
wire		RG_quantized_block_rl_42_en ;
wire		RG_quantized_block_rl_43_en ;
wire		RG_quantized_block_rl_44_en ;
wire		RG_quantized_block_rl_45_en ;
wire		RG_quantized_block_rl_46_en ;
wire		RG_quantized_block_rl_47_en ;
wire		RG_quantized_block_rl_48_en ;
wire		RG_quantized_block_rl_49_en ;
wire		RG_quantized_block_rl_50_en ;
wire		RG_quantized_block_rl_51_en ;
wire		RG_quantized_block_rl_52_en ;
wire		RG_quantized_block_rl_53_en ;
wire		RG_quantized_block_rl_54_en ;
wire		RG_quantized_block_rl_55_en ;
wire		RG_quantized_block_rl_56_en ;
wire		RG_quantized_block_rl_57_en ;
wire		RG_quantized_block_rl_58_en ;
wire		RG_quantized_block_rl_59_en ;
wire		RG_quantized_block_rl_60_en ;
wire		RG_quantized_block_rl_61_en ;
wire		RG_quantized_block_rl_62_en ;
wire		RL_previous_dc_quantized_block_en ;
wire		RG_k_01_en ;
wire		FF_d_01_en ;
wire		FF_i_en ;
wire		RG_rl_242_en ;
wire		RG_rl_243_en ;
wire		RG_rl_244_en ;
wire		RG_rl_245_en ;
wire		RG_rl_246_en ;
wire		RG_previous_dc_rl_1_en ;
wire		RG_len_en ;
wire		FF_len_en ;
wire		valid_r_en ;
reg	RG_M_14_d10_c7 ;
reg	RG_M_14_d10_c6 ;
reg	RG_M_14_d10_c5 ;
reg	RG_M_14_d10_c4 ;
reg	RG_M_14_d10_c3 ;
reg	RG_M_14_d10_c2 ;
reg	RG_M_14_d10_c1 ;
reg	RG_M_14_d10_c0 ;
reg	[8:0]	RG_rl_a127_d9_c7 ;
reg	[8:0]	RG_rl_a127_d9_c0 ;
reg	[8:0]	RG_rl_a126_d9_c7 ;
reg	[8:0]	RG_rl_a126_d9_c0 ;
reg	[8:0]	RG_rl_a125_d9_c7 ;
reg	[8:0]	RG_rl_a125_d9_c0 ;
reg	[8:0]	RG_rl_a124_d9_c7 ;
reg	[8:0]	RG_rl_a124_d9_c0 ;
reg	[8:0]	RG_rl_a123_d9_c7 ;
reg	[8:0]	RG_rl_a123_d9_c0 ;
reg	[8:0]	RG_rl_a122_d9_c7 ;
reg	[8:0]	RG_rl_a122_d9_c0 ;
reg	[8:0]	RG_rl_a121_d9_c7 ;
reg	[8:0]	RG_rl_a121_d9_c0 ;
reg	[8:0]	RG_rl_a120_d9_c7 ;
reg	[8:0]	RG_rl_a120_d9_c0 ;
reg	[8:0]	RG_rl_a119_d9_c7 ;
reg	[8:0]	RG_rl_a119_d9_c0 ;
reg	[8:0]	RG_rl_a118_d9_c7 ;
reg	[8:0]	RG_rl_a118_d9_c0 ;
reg	[8:0]	RG_rl_a117_d9_c7 ;
reg	[8:0]	RG_rl_a117_d9_c0 ;
reg	[8:0]	RG_rl_a116_d9_c7 ;
reg	[8:0]	RG_rl_a116_d9_c0 ;
reg	[8:0]	RG_rl_a115_d9_c7 ;
reg	[8:0]	RG_rl_a115_d9_c0 ;
reg	[8:0]	RG_rl_a114_d9_c7 ;
reg	[8:0]	RG_rl_a114_d9_c0 ;
reg	[8:0]	RG_rl_a113_d9_c7 ;
reg	[8:0]	RG_rl_a113_d9_c0 ;
reg	[8:0]	RG_rl_a112_d9_c7 ;
reg	[8:0]	RG_rl_a112_d9_c0 ;
reg	[8:0]	RG_rl_a111_d9_c6 ;
reg	[8:0]	RG_rl_a111_d9_c0 ;
reg	[8:0]	RG_rl_a110_d9_c6 ;
reg	[8:0]	RG_rl_a110_d9_c0 ;
reg	[8:0]	RG_rl_a109_d9_c6 ;
reg	[8:0]	RG_rl_a109_d9_c0 ;
reg	[8:0]	RG_rl_a108_d9_c6 ;
reg	[8:0]	RG_rl_a108_d9_c0 ;
reg	[8:0]	RG_rl_a107_d9_c6 ;
reg	[8:0]	RG_rl_a107_d9_c0 ;
reg	[8:0]	RG_rl_a106_d9_c6 ;
reg	[8:0]	RG_rl_a106_d9_c0 ;
reg	[8:0]	RG_rl_a105_d9_c6 ;
reg	[8:0]	RG_rl_a105_d9_c0 ;
reg	[8:0]	RG_rl_a104_d9_c6 ;
reg	[8:0]	RG_rl_a104_d9_c0 ;
reg	[8:0]	RG_rl_a103_d9_c6 ;
reg	[8:0]	RG_rl_a103_d9_c0 ;
reg	[8:0]	RG_rl_a102_d9_c6 ;
reg	[8:0]	RG_rl_a102_d9_c0 ;
reg	[8:0]	RG_rl_a101_d9_c6 ;
reg	[8:0]	RG_rl_a101_d9_c0 ;
reg	[8:0]	RG_rl_a100_d9_c6 ;
reg	[8:0]	RG_rl_a100_d9_c0 ;
reg	[8:0]	RG_rl_a99_d9_c6 ;
reg	[8:0]	RG_rl_a99_d9_c0 ;
reg	[8:0]	RG_rl_a98_d9_c6 ;
reg	[8:0]	RG_rl_a98_d9_c0 ;
reg	[8:0]	RG_rl_a97_d9_c6 ;
reg	[8:0]	RG_rl_a97_d9_c0 ;
reg	[8:0]	RG_rl_a96_d9_c6 ;
reg	[8:0]	RG_rl_a96_d9_c0 ;
reg	[8:0]	RG_rl_a95_d9_c5 ;
reg	[8:0]	RG_rl_a95_d9_c0 ;
reg	[8:0]	RG_rl_a94_d9_c5 ;
reg	[8:0]	RG_rl_a94_d9_c0 ;
reg	[8:0]	RG_rl_a93_d9_c5 ;
reg	[8:0]	RG_rl_a93_d9_c0 ;
reg	[8:0]	RG_rl_a92_d9_c5 ;
reg	[8:0]	RG_rl_a92_d9_c0 ;
reg	[8:0]	RG_rl_a91_d9_c5 ;
reg	[8:0]	RG_rl_a91_d9_c0 ;
reg	[8:0]	RG_rl_a90_d9_c5 ;
reg	[8:0]	RG_rl_a90_d9_c0 ;
reg	[8:0]	RG_rl_a89_d9_c5 ;
reg	[8:0]	RG_rl_a89_d9_c0 ;
reg	[8:0]	RG_rl_a88_d9_c5 ;
reg	[8:0]	RG_rl_a88_d9_c0 ;
reg	[8:0]	RG_rl_a87_d9_c5 ;
reg	[8:0]	RG_rl_a87_d9_c0 ;
reg	[8:0]	RG_rl_a86_d9_c5 ;
reg	[8:0]	RG_rl_a86_d9_c0 ;
reg	[8:0]	RG_rl_a85_d9_c5 ;
reg	[8:0]	RG_rl_a85_d9_c0 ;
reg	[8:0]	RG_rl_a84_d9_c5 ;
reg	[8:0]	RG_rl_a84_d9_c0 ;
reg	[8:0]	RG_rl_a83_d9_c5 ;
reg	[8:0]	RG_rl_a83_d9_c0 ;
reg	[8:0]	RG_rl_a82_d9_c5 ;
reg	[8:0]	RG_rl_a82_d9_c0 ;
reg	[8:0]	RG_rl_a81_d9_c5 ;
reg	[8:0]	RG_rl_a81_d9_c0 ;
reg	[8:0]	RG_rl_a80_d9_c5 ;
reg	[8:0]	RG_rl_a80_d9_c0 ;
reg	[8:0]	RG_rl_a79_d9_c4 ;
reg	[8:0]	RG_rl_a79_d9_c0 ;
reg	[8:0]	RG_rl_a78_d9_c4 ;
reg	[8:0]	RG_rl_a78_d9_c0 ;
reg	[8:0]	RG_rl_a77_d9_c4 ;
reg	[8:0]	RG_rl_a77_d9_c0 ;
reg	[8:0]	RG_rl_a76_d9_c4 ;
reg	[8:0]	RG_rl_a76_d9_c0 ;
reg	[8:0]	RG_rl_a75_d9_c4 ;
reg	[8:0]	RG_rl_a75_d9_c0 ;
reg	[8:0]	RG_rl_a74_d9_c4 ;
reg	[8:0]	RG_rl_a74_d9_c0 ;
reg	[8:0]	RG_rl_a73_d9_c4 ;
reg	[8:0]	RG_rl_a73_d9_c0 ;
reg	[8:0]	RG_rl_a72_d9_c4 ;
reg	[8:0]	RG_rl_a72_d9_c0 ;
reg	[8:0]	RG_rl_a71_d9_c4 ;
reg	[8:0]	RG_rl_a71_d9_c0 ;
reg	[8:0]	RG_rl_a70_d9_c4 ;
reg	[8:0]	RG_rl_a70_d9_c0 ;
reg	[8:0]	RG_rl_a69_d9_c4 ;
reg	[8:0]	RG_rl_a69_d9_c0 ;
reg	[8:0]	RG_rl_a68_d9_c4 ;
reg	[8:0]	RG_rl_a68_d9_c0 ;
reg	[8:0]	RG_rl_a67_d9_c4 ;
reg	[8:0]	RG_rl_a67_d9_c0 ;
reg	[8:0]	RG_rl_a66_d9_c4 ;
reg	[8:0]	RG_rl_a66_d9_c0 ;
reg	[8:0]	RG_rl_a65_d9_c4 ;
reg	[8:0]	RG_rl_a65_d9_c0 ;
reg	[8:0]	RG_rl_a64_d9_c4 ;
reg	[8:0]	RG_rl_a64_d9_c0 ;
reg	[8:0]	RG_rl_a63_d9_c3 ;
reg	[8:0]	RG_rl_a63_d9_c0 ;
reg	[8:0]	RG_rl_a62_d9_c3 ;
reg	[8:0]	RG_rl_a62_d9_c0 ;
reg	[8:0]	RG_rl_a61_d9_c3 ;
reg	[8:0]	RG_rl_a61_d9_c0 ;
reg	[8:0]	RG_rl_a60_d9_c3 ;
reg	[8:0]	RG_rl_a60_d9_c0 ;
reg	[8:0]	RG_rl_a59_d9_c3 ;
reg	[8:0]	RG_rl_a59_d9_c0 ;
reg	[8:0]	RG_rl_a58_d9_c3 ;
reg	[8:0]	RG_rl_a58_d9_c0 ;
reg	[8:0]	RG_rl_a57_d9_c3 ;
reg	[8:0]	RG_rl_a57_d9_c0 ;
reg	[8:0]	RG_rl_a56_d9_c3 ;
reg	[8:0]	RG_rl_a56_d9_c0 ;
reg	[8:0]	RG_rl_a55_d9_c3 ;
reg	[8:0]	RG_rl_a55_d9_c0 ;
reg	[8:0]	RG_rl_a54_d9_c3 ;
reg	[8:0]	RG_rl_a54_d9_c0 ;
reg	[8:0]	RG_rl_a53_d9_c3 ;
reg	[8:0]	RG_rl_a53_d9_c0 ;
reg	[8:0]	RG_rl_a52_d9_c3 ;
reg	[8:0]	RG_rl_a52_d9_c0 ;
reg	[8:0]	RG_rl_a51_d9_c3 ;
reg	[8:0]	RG_rl_a51_d9_c0 ;
reg	[8:0]	RG_rl_a50_d9_c3 ;
reg	[8:0]	RG_rl_a50_d9_c0 ;
reg	[8:0]	RG_rl_a49_d9_c3 ;
reg	[8:0]	RG_rl_a49_d9_c0 ;
reg	[8:0]	RG_rl_a48_d9_c3 ;
reg	[8:0]	RG_rl_a48_d9_c0 ;
reg	[8:0]	RG_rl_a47_d9_c2 ;
reg	[8:0]	RG_rl_a47_d9_c0 ;
reg	[8:0]	RG_rl_a46_d9_c2 ;
reg	[8:0]	RG_rl_a46_d9_c0 ;
reg	[8:0]	RG_rl_a45_d9_c2 ;
reg	[8:0]	RG_rl_a45_d9_c0 ;
reg	[8:0]	RG_rl_a44_d9_c2 ;
reg	[8:0]	RG_rl_a44_d9_c0 ;
reg	[8:0]	RG_rl_a43_d9_c2 ;
reg	[8:0]	RG_rl_a43_d9_c0 ;
reg	[8:0]	RG_rl_a42_d9_c2 ;
reg	[8:0]	RG_rl_a42_d9_c0 ;
reg	[8:0]	RG_rl_a41_d9_c2 ;
reg	[8:0]	RG_rl_a41_d9_c0 ;
reg	[8:0]	RG_rl_a40_d9_c2 ;
reg	[8:0]	RG_rl_a40_d9_c0 ;
reg	[8:0]	RG_rl_a39_d9_c2 ;
reg	[8:0]	RG_rl_a39_d9_c0 ;
reg	[8:0]	RG_rl_a38_d9_c2 ;
reg	[8:0]	RG_rl_a38_d9_c0 ;
reg	[8:0]	RG_rl_a37_d9_c2 ;
reg	[8:0]	RG_rl_a37_d9_c0 ;
reg	[8:0]	RG_rl_a36_d9_c2 ;
reg	[8:0]	RG_rl_a36_d9_c0 ;
reg	[8:0]	RG_rl_a35_d9_c2 ;
reg	[8:0]	RG_rl_a35_d9_c0 ;
reg	[8:0]	RG_rl_a34_d9_c2 ;
reg	[8:0]	RG_rl_a34_d9_c0 ;
reg	[8:0]	RG_rl_a33_d9_c2 ;
reg	[8:0]	RG_rl_a33_d9_c0 ;
reg	[8:0]	RG_rl_a32_d9_c2 ;
reg	[8:0]	RG_rl_a32_d9_c0 ;
reg	[8:0]	RG_rl_a31_d9_c1 ;
reg	[8:0]	RG_rl_a31_d9_c0 ;
reg	[8:0]	RG_rl_a30_d9_c1 ;
reg	[8:0]	RG_rl_a30_d9_c0 ;
reg	[8:0]	RG_rl_a29_d9_c1 ;
reg	[8:0]	RG_rl_a29_d9_c0 ;
reg	[8:0]	RG_rl_a28_d9_c1 ;
reg	[8:0]	RG_rl_a28_d9_c0 ;
reg	[8:0]	RG_rl_a27_d9_c1 ;
reg	[8:0]	RG_rl_a27_d9_c0 ;
reg	[8:0]	RG_rl_a26_d9_c1 ;
reg	[8:0]	RG_rl_a26_d9_c0 ;
reg	[8:0]	RG_rl_a25_d9_c1 ;
reg	[8:0]	RG_rl_a25_d9_c0 ;
reg	[8:0]	RG_rl_a24_d9_c1 ;
reg	[8:0]	RG_rl_a24_d9_c0 ;
reg	[8:0]	RG_rl_a23_d9_c1 ;
reg	[8:0]	RG_rl_a23_d9_c0 ;
reg	[8:0]	RG_rl_a22_d9_c1 ;
reg	[8:0]	RG_rl_a22_d9_c0 ;
reg	[8:0]	RG_rl_a21_d9_c1 ;
reg	[8:0]	RG_rl_a21_d9_c0 ;
reg	[8:0]	RG_rl_a20_d9_c1 ;
reg	[8:0]	RG_rl_a20_d9_c0 ;
reg	[8:0]	RG_rl_a19_d9_c1 ;
reg	[8:0]	RG_rl_a19_d9_c0 ;
reg	[8:0]	RG_rl_a18_d9_c1 ;
reg	[8:0]	RG_rl_a18_d9_c0 ;
reg	[8:0]	RG_rl_a17_d9_c1 ;
reg	[8:0]	RG_rl_a17_d9_c0 ;
reg	[8:0]	RG_rl_a16_d9_c1 ;
reg	[8:0]	RG_rl_a16_d9_c0 ;
reg	[8:0]	RG_rl_a15_d9_c1 ;
reg	[8:0]	RG_rl_a15_d9_c0 ;
reg	[8:0]	RG_rl_a14_d9_c1 ;
reg	[8:0]	RG_rl_a14_d9_c0 ;
reg	[8:0]	RG_rl_a13_d9_c1 ;
reg	[8:0]	RG_rl_a13_d9_c0 ;
reg	[8:0]	RG_rl_a12_d9_c1 ;
reg	[8:0]	RG_rl_a12_d9_c0 ;
reg	[8:0]	RG_rl_a11_d9_c1 ;
reg	[8:0]	RG_rl_a11_d9_c0 ;
reg	[8:0]	RG_rl_a10_d9_c1 ;
reg	[8:0]	RG_rl_a10_d9_c0 ;
reg	[8:0]	RG_rl_a09_d9_c1 ;
reg	[8:0]	RG_rl_a09_d9_c0 ;
reg	[8:0]	RG_rl_a08_d9_c1 ;
reg	[8:0]	RG_rl_a08_d9_c0 ;
reg	[8:0]	RG_rl_a07_d9_c1 ;
reg	[8:0]	RG_rl_a07_d9_c0 ;
reg	[8:0]	RG_rl_a06_d9_c1 ;
reg	[8:0]	RG_rl_a06_d9_c0 ;
reg	[8:0]	RG_rl_a05_d9_c1 ;
reg	[8:0]	RG_rl_a05_d9_c0 ;
reg	[8:0]	RG_rl_a04_d9_c1 ;
reg	[8:0]	RG_rl_a04_d9_c0 ;
reg	[8:0]	RG_rl_a03_d9_c1 ;
reg	[8:0]	RG_rl_a03_d9_c0 ;
reg	[8:0]	RG_rl_a02_d9_c1 ;
reg	[8:0]	RG_rl_a02_d9_c0 ;
reg	[8:0]	RG_rl_a01_d9_c1 ;
reg	[8:0]	RG_rl_a01_d9_c0 ;
reg	[8:0]	RG_rl_a00_d9_c1 ;
reg	[8:0]	RG_rl_a00_d9_c0 ;
reg	[8:0]	RG_rl ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_1 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_2 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_3 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_4 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_5 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_6 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_7 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_8 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_9 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_10 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_11 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_12 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_13 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_14 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_15 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_16 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_17 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_18 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_19 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_20 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_21 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_22 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_23 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_24 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_25 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_26 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_27 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_28 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_29 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_30 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_31 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_32 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_33 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_34 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_35 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_36 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_37 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_38 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_39 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_40 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_41 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_42 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_43 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_44 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_45 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_46 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_47 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_48 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_49 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_50 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_51 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_52 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_53 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_54 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_55 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_56 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_57 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_58 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_59 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_60 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_61 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_62 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_63 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_64 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_65 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_66 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_67 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_68 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_69 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_70 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_71 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_72 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_73 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_74 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_75 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_76 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_77 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_78 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_79 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_80 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_81 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_82 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_83 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_84 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_85 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_86 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_87 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_88 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_89 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_90 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_91 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_92 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_93 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_94 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_95 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_96 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_97 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_98 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_99 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_100 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_101 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_102 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_103 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_104 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_105 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_106 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_107 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_108 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_109 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_110 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_111 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_112 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_113 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_114 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_115 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_116 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_117 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_118 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_119 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_120 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_121 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_122 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_123 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_124 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_125 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_126 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_127 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_previous_dc ;	// line#=../rle.h:66
reg	[8:0]	RG_rl_128 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_129 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_130 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_131 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_132 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_133 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_134 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_135 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_136 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_137 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_138 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_139 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_140 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_141 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_142 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_143 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_144 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_145 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_146 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_147 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_148 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_149 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_150 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_151 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_152 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_153 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_154 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_155 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_156 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_157 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_158 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_159 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_160 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_161 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_162 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_163 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_164 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_165 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_166 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_167 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_168 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_169 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_170 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_171 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_172 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_173 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_174 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_175 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_176 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_177 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_178 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_179 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_180 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_181 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_182 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_183 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_184 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_previous_dc_rl ;	// line#=../rle.h:66 ../rle.cpp:23
reg	[8:0]	RG_rl_185 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_186 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_187 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_188 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_189 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_190 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_191 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_192 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_193 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_194 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_195 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_196 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_197 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_198 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_199 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_200 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_201 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_202 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_203 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_204 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_205 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_206 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_207 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_208 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_209 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_210 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_211 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_212 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_213 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_214 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_215 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_216 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_217 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_218 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_219 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_220 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_221 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_222 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_223 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_224 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_225 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_226 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_227 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_228 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_229 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_230 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_231 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_232 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_233 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_234 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_235 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_236 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_237 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_238 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_239 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_240 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_241 ;	// line#=../rle.cpp:23
reg	[3:0]	RG_j ;	// line#=../rle.cpp:27
reg	[31:0]	RG_i_k_01 ;	// line#=../rle.cpp:25,105
reg	[31:0]	RG_i_j_01 ;	// line#=../rle.cpp:25,105
reg	[8:0]	RG_quantized_block_rl ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_1 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_2 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_3 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_4 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_5 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_6 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_7 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_8 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_9 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_10 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_11 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_12 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_13 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_14 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_15 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_16 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_17 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_18 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_19 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_20 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_21 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_22 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_23 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_24 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_25 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_26 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_27 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_28 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_29 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_30 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_31 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_32 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_33 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_34 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_35 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_36 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_37 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_38 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_39 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_40 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_41 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_42 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_43 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_44 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_45 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_46 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_47 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_48 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_49 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_50 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_51 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_52 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_53 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_54 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_55 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_56 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_57 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_58 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_59 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_60 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_61 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RG_quantized_block_rl_62 ;	// line#=../rle.cpp:22,23
reg	[8:0]	RL_previous_dc_quantized_block ;	// line#=../rle.cpp:22,23 ../rle.h:66
reg	[6:0]	RG_k_01 ;	// line#=../rle.cpp:105
reg	FF_d_01 ;	// line#=../rle.cpp:105
reg	FF_j ;	// line#=../rle.cpp:27
reg	FF_i ;	// line#=../rle.cpp:25
reg	RG_315 ;
reg	[8:0]	RG_rl_242 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_243 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_244 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_245 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_rl_246 ;	// line#=../rle.cpp:23
reg	[8:0]	RG_previous_dc_rl_1 ;	// line#=../rle.cpp:23 ../rle.h:66
reg	[7:0]	RG_len_01 ;	// line#=../rle.cpp:24
reg	[6:0]	RG_323 ;
reg	RG_324 ;
reg	RG_325 ;
reg	RG_326 ;
reg	RG_327 ;
reg	RG_328 ;
reg	RG_329 ;
reg	RG_330 ;
reg	RG_331 ;
reg	RG_332 ;
reg	RG_333 ;
reg	RG_334 ;
reg	RG_335 ;
reg	RG_336 ;
reg	RG_337 ;
reg	RG_338 ;
reg	RG_339 ;
reg	RG_340 ;
reg	RG_341 ;
reg	RG_342 ;
reg	RG_343 ;
reg	RG_344 ;
reg	RG_345 ;
reg	RG_346 ;
reg	RG_347 ;
reg	RG_348 ;
reg	RG_349 ;
reg	RG_350 ;
reg	RG_351 ;
reg	RG_352 ;
reg	RG_353 ;
reg	RG_354 ;
reg	RG_355 ;
reg	RG_356 ;
reg	RG_357 ;
reg	RG_358 ;
reg	RG_359 ;
reg	RG_360 ;
reg	RG_361 ;
reg	RG_362 ;
reg	RG_363 ;
reg	RG_364 ;
reg	RG_365 ;
reg	RG_366 ;
reg	RG_367 ;
reg	RG_368 ;
reg	RG_369 ;
reg	RG_370 ;
reg	RG_371 ;
reg	RG_372 ;
reg	RG_373 ;
reg	RG_374 ;
reg	RG_375 ;
reg	RG_376 ;
reg	RG_377 ;
reg	RG_378 ;
reg	RG_379 ;
reg	RG_380 ;
reg	RG_381 ;
reg	RG_382 ;
reg	RG_383 ;
reg	RG_384 ;
reg	RG_385 ;
reg	[7:0]	RG_len ;	// line#=../rle.cpp:24
reg	RG_387 ;
reg	RG_388 ;
reg	RG_389 ;
reg	RG_390 ;
reg	RG_391 ;
reg	RG_392 ;
reg	RG_393 ;
reg	RG_394 ;
reg	RG_395 ;
reg	RG_396 ;
reg	RG_397 ;
reg	RG_398 ;
reg	RG_399 ;
reg	RG_400 ;
reg	RG_401 ;
reg	RG_402 ;
reg	RG_403 ;
reg	RG_404 ;
reg	RG_405 ;
reg	RG_406 ;
reg	RG_407 ;
reg	RG_408 ;
reg	RG_409 ;
reg	RG_410 ;
reg	RG_411 ;
reg	RG_412 ;
reg	RG_413 ;
reg	RG_414 ;
reg	RG_415 ;
reg	RG_416 ;
reg	RG_417 ;
reg	RG_418 ;
reg	RG_419 ;
reg	RG_420 ;
reg	RG_421 ;
reg	RG_422 ;
reg	RG_423 ;
reg	RG_424 ;
reg	RG_425 ;
reg	RG_426 ;
reg	RG_427 ;
reg	RG_428 ;
reg	RG_429 ;
reg	RG_430 ;
reg	RG_431 ;
reg	RG_432 ;
reg	RG_433 ;
reg	RG_434 ;
reg	RG_435 ;
reg	RG_436 ;
reg	RG_437 ;
reg	RG_438 ;
reg	RG_439 ;
reg	RG_440 ;
reg	RG_441 ;
reg	RG_442 ;
reg	RG_443 ;
reg	RG_444 ;
reg	RG_445 ;
reg	RG_446 ;
reg	RG_447 ;
reg	RG_448 ;
reg	RG_449 ;
reg	RG_450 ;
reg	RG_451 ;
reg	FF_len ;	// line#=../rle.cpp:24
reg	[8:0]	jpeg_out_a00_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a01_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a02_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a03_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a04_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a05_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a06_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a07_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a08_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a09_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a10_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a11_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a12_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a13_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a14_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a15_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a16_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a17_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a18_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a19_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a20_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a21_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a22_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a23_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a24_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a25_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a26_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a27_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a28_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a29_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a30_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a31_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a32_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a33_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a34_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a35_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a36_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a37_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a38_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a39_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a40_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a41_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a42_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a43_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a44_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a45_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a46_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a47_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a48_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a49_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a50_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a51_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a52_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a53_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a54_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a55_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a56_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a57_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a58_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a59_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a60_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a61_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a62_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a63_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a64_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a65_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a66_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a67_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a68_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a69_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a70_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a71_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a72_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a73_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a74_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a75_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a76_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a77_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a78_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a79_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a80_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a81_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a82_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a83_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a84_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a85_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a86_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a87_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a88_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a89_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a90_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a91_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a92_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a93_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a94_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a95_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a96_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a97_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a98_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a99_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a100_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a101_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a102_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a103_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a104_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a105_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a106_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a107_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a108_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a109_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a110_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a111_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a112_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a113_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a114_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a115_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a116_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a117_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a118_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a119_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a120_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a121_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a122_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a123_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a124_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a125_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a126_r ;	// line#=../rle.h:60
reg	[8:0]	jpeg_out_a127_r ;	// line#=../rle.h:60
reg	[11:0]	jpeg_len_out_r ;	// line#=../rle.h:61
reg	valid_r ;	// line#=../rle.h:62
reg	M_01_t1 ;
reg	[8:0]	TR_12 ;
reg	[8:0]	TR_13 ;
reg	[8:0]	TR_14 ;
reg	[8:0]	TR_15 ;
reg	[8:0]	TR_16 ;
reg	[8:0]	TR_17 ;
reg	[8:0]	TR_18 ;
reg	[8:0]	TR_19 ;
reg	[8:0]	TR_20 ;
reg	[8:0]	TR_21 ;
reg	[8:0]	TR_22 ;
reg	[8:0]	TR_23 ;
reg	[8:0]	TR_24 ;
reg	[8:0]	TR_25 ;
reg	[8:0]	TR_26 ;
reg	[8:0]	TR_27 ;
reg	[8:0]	TR_28 ;
reg	[8:0]	TR_29 ;
reg	[8:0]	TR_30 ;
reg	[8:0]	TR_31 ;
reg	[8:0]	TR_32 ;
reg	[8:0]	TR_33 ;
reg	[8:0]	TR_34 ;
reg	[8:0]	TR_35 ;
reg	[8:0]	TR_36 ;
reg	[8:0]	TR_37 ;
reg	[8:0]	TR_38 ;
reg	[8:0]	TR_39 ;
reg	[8:0]	TR_40 ;
reg	[8:0]	TR_41 ;
reg	[8:0]	TR_42 ;
reg	[8:0]	TR_43 ;
reg	[8:0]	TR_44 ;
reg	[8:0]	TR_45 ;
reg	[8:0]	TR_46 ;
reg	[8:0]	TR_47 ;
reg	[8:0]	TR_48 ;
reg	[8:0]	TR_49 ;
reg	[8:0]	TR_50 ;
reg	[8:0]	TR_51 ;
reg	[8:0]	TR_52 ;
reg	[8:0]	TR_53 ;
reg	[8:0]	TR_54 ;
reg	[8:0]	TR_55 ;
reg	[8:0]	TR_56 ;
reg	[8:0]	TR_57 ;
reg	[8:0]	TR_58 ;
reg	[8:0]	TR_59 ;
reg	[8:0]	TR_60 ;
reg	[8:0]	TR_61 ;
reg	[8:0]	TR_62 ;
reg	[8:0]	TR_63 ;
reg	[8:0]	TR_64 ;
reg	[8:0]	TR_65 ;
reg	[8:0]	TR_66 ;
reg	[8:0]	TR_67 ;
reg	[8:0]	TR_68 ;
reg	[8:0]	TR_69 ;
reg	[8:0]	TR_70 ;
reg	[8:0]	TR_71 ;
reg	[8:0]	TR_72 ;
reg	[8:0]	TR_73 ;
reg	[8:0]	TR_74 ;
reg	[8:0]	TR_75 ;
reg	[8:0]	TR_76 ;
reg	[8:0]	TR_77 ;
reg	[8:0]	TR_78 ;
reg	[8:0]	TR_79 ;
reg	[8:0]	TR_80 ;
reg	[8:0]	TR_81 ;
reg	[8:0]	TR_82 ;
reg	[8:0]	TR_83 ;
reg	[8:0]	TR_84 ;
reg	[8:0]	TR_85 ;
reg	[8:0]	TR_86 ;
reg	[8:0]	TR_87 ;
reg	[8:0]	TR_88 ;
reg	[8:0]	TR_89 ;
reg	[8:0]	TR_90 ;
reg	[8:0]	TR_91 ;
reg	[8:0]	TR_92 ;
reg	[8:0]	TR_93 ;
reg	[8:0]	TR_94 ;
reg	[8:0]	TR_95 ;
reg	[8:0]	TR_96 ;
reg	[8:0]	TR_97 ;
reg	[8:0]	TR_98 ;
reg	[8:0]	TR_99 ;
reg	[8:0]	TR_100 ;
reg	[8:0]	TR_101 ;
reg	[8:0]	TR_102 ;
reg	[8:0]	TR_103 ;
reg	[8:0]	TR_104 ;
reg	[8:0]	TR_105 ;
reg	[8:0]	TR_106 ;
reg	[8:0]	TR_107 ;
reg	[8:0]	TR_108 ;
reg	[8:0]	TR_109 ;
reg	[8:0]	TR_110 ;
reg	[8:0]	TR_111 ;
reg	[8:0]	TR_112 ;
reg	[8:0]	TR_113 ;
reg	[8:0]	TR_114 ;
reg	[8:0]	TR_115 ;
reg	[8:0]	TR_116 ;
reg	[8:0]	TR_117 ;
reg	[8:0]	TR_118 ;
reg	[8:0]	TR_119 ;
reg	[8:0]	TR_120 ;
reg	[8:0]	TR_121 ;
reg	[8:0]	TR_122 ;
reg	[8:0]	TR_123 ;
reg	[8:0]	TR_124 ;
reg	[8:0]	TR_125 ;
reg	[8:0]	TR_126 ;
reg	[8:0]	TR_127 ;
reg	[8:0]	TR_128 ;
reg	[8:0]	TR_129 ;
reg	[8:0]	TR_130 ;
reg	[8:0]	TR_131 ;
reg	[8:0]	TR_132 ;
reg	[8:0]	TR_133 ;
reg	[8:0]	TR_134 ;
reg	[8:0]	TR_135 ;
reg	[8:0]	TR_136 ;
reg	[8:0]	TR_137 ;
reg	[8:0]	TR_138 ;
reg	[8:0]	TR_11 ;
reg	[8:0]	RG_rl_a00_d9_c0_t ;
reg	[8:0]	RG_rl_a01_d9_c0_t ;
reg	[8:0]	RG_rl_a02_d9_c0_t ;
reg	[8:0]	RG_rl_a03_d9_c0_t ;
reg	[8:0]	RG_rl_a04_d9_c0_t ;
reg	[8:0]	RG_rl_a05_d9_c0_t ;
reg	[8:0]	RG_rl_a06_d9_c0_t ;
reg	[8:0]	RG_rl_a07_d9_c0_t ;
reg	[8:0]	RG_rl_a08_d9_c0_t ;
reg	[8:0]	RG_rl_a09_d9_c0_t ;
reg	[8:0]	RG_rl_a10_d9_c0_t ;
reg	[8:0]	RG_rl_a11_d9_c0_t ;
reg	[8:0]	RG_rl_a12_d9_c0_t ;
reg	[8:0]	RG_rl_a13_d9_c0_t ;
reg	[8:0]	RG_rl_a14_d9_c0_t ;
reg	[8:0]	RG_rl_a15_d9_c0_t ;
reg	[8:0]	RG_rl_a16_d9_c1_t ;
reg	[8:0]	RG_rl_a17_d9_c1_t ;
reg	[8:0]	RG_rl_a18_d9_c1_t ;
reg	[8:0]	RG_rl_a19_d9_c1_t ;
reg	[8:0]	RG_rl_a20_d9_c1_t ;
reg	[8:0]	RG_rl_a21_d9_c1_t ;
reg	[8:0]	RG_rl_a22_d9_c1_t ;
reg	[8:0]	RG_rl_a23_d9_c1_t ;
reg	[8:0]	RG_rl_a24_d9_c1_t ;
reg	[8:0]	RG_rl_a25_d9_c1_t ;
reg	[8:0]	RG_rl_a26_d9_c1_t ;
reg	[8:0]	RG_rl_a27_d9_c1_t ;
reg	[8:0]	RG_rl_a28_d9_c1_t ;
reg	[8:0]	RG_rl_a29_d9_c1_t ;
reg	[8:0]	RG_rl_a30_d9_c1_t ;
reg	[8:0]	RG_rl_a31_d9_c1_t ;
reg	[8:0]	RG_rl_a32_d9_c2_t ;
reg	[8:0]	RG_rl_a33_d9_c2_t ;
reg	[8:0]	RG_rl_a34_d9_c2_t ;
reg	[8:0]	RG_rl_a35_d9_c2_t ;
reg	[8:0]	RG_rl_a36_d9_c2_t ;
reg	[8:0]	RG_rl_a37_d9_c2_t ;
reg	[8:0]	RG_rl_a38_d9_c2_t ;
reg	[8:0]	RG_rl_a39_d9_c2_t ;
reg	[8:0]	RG_rl_a40_d9_c2_t ;
reg	[8:0]	RG_rl_a41_d9_c2_t ;
reg	[8:0]	RG_rl_a42_d9_c2_t ;
reg	[8:0]	RG_rl_a43_d9_c2_t ;
reg	[8:0]	RG_rl_a44_d9_c2_t ;
reg	[8:0]	RG_rl_a45_d9_c2_t ;
reg	[8:0]	RG_rl_a46_d9_c2_t ;
reg	[8:0]	RG_rl_a47_d9_c2_t ;
reg	[8:0]	RG_rl_a48_d9_c3_t ;
reg	[8:0]	RG_rl_a49_d9_c3_t ;
reg	[8:0]	RG_rl_a50_d9_c3_t ;
reg	[8:0]	RG_rl_a51_d9_c3_t ;
reg	[8:0]	RG_rl_a52_d9_c3_t ;
reg	[8:0]	RG_rl_a53_d9_c3_t ;
reg	[8:0]	RG_rl_a54_d9_c3_t ;
reg	[8:0]	RG_rl_a55_d9_c3_t ;
reg	[8:0]	RG_rl_a56_d9_c3_t ;
reg	[8:0]	RG_rl_a57_d9_c3_t ;
reg	[8:0]	RG_rl_a58_d9_c3_t ;
reg	[8:0]	RG_rl_a59_d9_c3_t ;
reg	[8:0]	RG_rl_a60_d9_c3_t ;
reg	[8:0]	RG_rl_a61_d9_c3_t ;
reg	[8:0]	RG_rl_a62_d9_c3_t ;
reg	[8:0]	RG_rl_a63_d9_c3_t ;
reg	[8:0]	RG_rl_a64_d9_c4_t ;
reg	[8:0]	RG_rl_a65_d9_c4_t ;
reg	[8:0]	RG_rl_a66_d9_c4_t ;
reg	[8:0]	RG_rl_a67_d9_c4_t ;
reg	[8:0]	RG_rl_a68_d9_c4_t ;
reg	[8:0]	RG_rl_a69_d9_c4_t ;
reg	[8:0]	RG_rl_a70_d9_c4_t ;
reg	[8:0]	RG_rl_a71_d9_c4_t ;
reg	[8:0]	RG_rl_a72_d9_c4_t ;
reg	[8:0]	RG_rl_a73_d9_c4_t ;
reg	[8:0]	RG_rl_a74_d9_c4_t ;
reg	[8:0]	RG_rl_a75_d9_c4_t ;
reg	[8:0]	RG_rl_a76_d9_c4_t ;
reg	[8:0]	RG_rl_a77_d9_c4_t ;
reg	[8:0]	RG_rl_a78_d9_c4_t ;
reg	[8:0]	RG_rl_a79_d9_c4_t ;
reg	[8:0]	RG_rl_a80_d9_c5_t ;
reg	[8:0]	RG_rl_a81_d9_c5_t ;
reg	[8:0]	RG_rl_a82_d9_c5_t ;
reg	[8:0]	RG_rl_a83_d9_c5_t ;
reg	[8:0]	RG_rl_a84_d9_c5_t ;
reg	[8:0]	RG_rl_a85_d9_c5_t ;
reg	[8:0]	RG_rl_a86_d9_c5_t ;
reg	[8:0]	RG_rl_a87_d9_c5_t ;
reg	[8:0]	RG_rl_a88_d9_c5_t ;
reg	[8:0]	RG_rl_a89_d9_c5_t ;
reg	[8:0]	RG_rl_a90_d9_c5_t ;
reg	[8:0]	RG_rl_a91_d9_c5_t ;
reg	[8:0]	RG_rl_a92_d9_c5_t ;
reg	[8:0]	RG_rl_a93_d9_c5_t ;
reg	[8:0]	RG_rl_a94_d9_c5_t ;
reg	[8:0]	RG_rl_a95_d9_c5_t ;
reg	[8:0]	RG_rl_a96_d9_c6_t ;
reg	[8:0]	RG_rl_a97_d9_c6_t ;
reg	[8:0]	RG_rl_a98_d9_c6_t ;
reg	[8:0]	RG_rl_a99_d9_c6_t ;
reg	[8:0]	RG_rl_a100_d9_c6_t ;
reg	[8:0]	RG_rl_a101_d9_c6_t ;
reg	[8:0]	RG_rl_a102_d9_c6_t ;
reg	[8:0]	RG_rl_a103_d9_c6_t ;
reg	[8:0]	RG_rl_a104_d9_c6_t ;
reg	[8:0]	RG_rl_a105_d9_c6_t ;
reg	[8:0]	RG_rl_a106_d9_c6_t ;
reg	[8:0]	RG_rl_a107_d9_c6_t ;
reg	[8:0]	RG_rl_a108_d9_c6_t ;
reg	[8:0]	RG_rl_a109_d9_c6_t ;
reg	[8:0]	RG_rl_a110_d9_c6_t ;
reg	[8:0]	RG_rl_a111_d9_c6_t ;
reg	[8:0]	RG_rl_a112_d9_c7_t ;
reg	[8:0]	RG_rl_a113_d9_c7_t ;
reg	[8:0]	RG_rl_a114_d9_c7_t ;
reg	[8:0]	RG_rl_a115_d9_c7_t ;
reg	[8:0]	RG_rl_a116_d9_c7_t ;
reg	[8:0]	RG_rl_a117_d9_c7_t ;
reg	[8:0]	RG_rl_a118_d9_c7_t ;
reg	[8:0]	RG_rl_a119_d9_c7_t ;
reg	[8:0]	RG_rl_a120_d9_c7_t ;
reg	[8:0]	RG_rl_a121_d9_c7_t ;
reg	[8:0]	RG_rl_a122_d9_c7_t ;
reg	[8:0]	RG_rl_a123_d9_c7_t ;
reg	[8:0]	RG_rl_a124_d9_c7_t ;
reg	[8:0]	RG_rl_a125_d9_c7_t ;
reg	[8:0]	RG_rl_a126_d9_c7_t ;
reg	[8:0]	RG_rl_a127_d9_c7_t ;
reg	[8:0]	rl_a00_t5 ;
reg	[8:0]	rl_a01_t5 ;
reg	[8:0]	rl_a02_t5 ;
reg	[8:0]	rl_a03_t5 ;
reg	[8:0]	rl_a04_t5 ;
reg	[8:0]	rl_a05_t5 ;
reg	[8:0]	rl_a06_t5 ;
reg	[8:0]	rl_a07_t5 ;
reg	[8:0]	rl_a08_t5 ;
reg	[8:0]	rl_a09_t5 ;
reg	[8:0]	rl_a10_t5 ;
reg	[8:0]	rl_a11_t5 ;
reg	[8:0]	rl_a12_t5 ;
reg	[8:0]	rl_a13_t5 ;
reg	[8:0]	rl_a14_t5 ;
reg	[8:0]	rl_a15_t5 ;
reg	[8:0]	rl_a16_t5 ;
reg	[8:0]	rl_a17_t5 ;
reg	[8:0]	rl_a18_t5 ;
reg	[8:0]	rl_a19_t5 ;
reg	[8:0]	rl_a20_t5 ;
reg	[8:0]	rl_a21_t5 ;
reg	[8:0]	rl_a22_t5 ;
reg	[8:0]	rl_a23_t5 ;
reg	[8:0]	rl_a24_t5 ;
reg	[8:0]	rl_a25_t5 ;
reg	[8:0]	rl_a26_t5 ;
reg	[8:0]	rl_a27_t5 ;
reg	[8:0]	rl_a28_t5 ;
reg	[8:0]	rl_a29_t5 ;
reg	[8:0]	rl_a30_t5 ;
reg	[8:0]	rl_a31_t5 ;
reg	[8:0]	rl_a32_t5 ;
reg	[8:0]	rl_a33_t5 ;
reg	[8:0]	rl_a34_t5 ;
reg	[8:0]	rl_a35_t5 ;
reg	[8:0]	rl_a36_t5 ;
reg	[8:0]	rl_a37_t5 ;
reg	[8:0]	rl_a38_t5 ;
reg	[8:0]	rl_a39_t5 ;
reg	[8:0]	rl_a40_t5 ;
reg	[8:0]	rl_a41_t5 ;
reg	[8:0]	rl_a42_t5 ;
reg	[8:0]	rl_a43_t5 ;
reg	[8:0]	rl_a44_t5 ;
reg	[8:0]	rl_a45_t5 ;
reg	[8:0]	rl_a46_t5 ;
reg	[8:0]	rl_a47_t5 ;
reg	[8:0]	rl_a48_t5 ;
reg	[8:0]	rl_a49_t5 ;
reg	[8:0]	rl_a50_t5 ;
reg	[8:0]	rl_a51_t5 ;
reg	[8:0]	rl_a52_t5 ;
reg	[8:0]	rl_a53_t5 ;
reg	[8:0]	rl_a54_t5 ;
reg	[8:0]	rl_a55_t5 ;
reg	[8:0]	rl_a56_t5 ;
reg	[8:0]	rl_a57_t5 ;
reg	[8:0]	rl_a58_t5 ;
reg	[8:0]	rl_a59_t5 ;
reg	[8:0]	rl_a60_t5 ;
reg	[8:0]	rl_a61_t5 ;
reg	[8:0]	rl_a62_t5 ;
reg	[8:0]	rl_a63_t5 ;
reg	[8:0]	rl_a64_t5 ;
reg	[8:0]	rl_a65_t5 ;
reg	[8:0]	rl_a66_t5 ;
reg	[8:0]	rl_a67_t5 ;
reg	[8:0]	rl_a68_t5 ;
reg	[8:0]	rl_a69_t5 ;
reg	[8:0]	rl_a70_t5 ;
reg	[8:0]	rl_a71_t5 ;
reg	[8:0]	rl_a72_t5 ;
reg	[8:0]	rl_a73_t5 ;
reg	[8:0]	rl_a74_t5 ;
reg	[8:0]	rl_a75_t5 ;
reg	[8:0]	rl_a76_t5 ;
reg	[8:0]	rl_a77_t5 ;
reg	[8:0]	rl_a78_t5 ;
reg	[8:0]	rl_a79_t5 ;
reg	[8:0]	rl_a80_t5 ;
reg	[8:0]	rl_a81_t5 ;
reg	[8:0]	rl_a82_t5 ;
reg	[8:0]	rl_a83_t5 ;
reg	[8:0]	rl_a84_t5 ;
reg	[8:0]	rl_a85_t5 ;
reg	[8:0]	rl_a86_t5 ;
reg	[8:0]	rl_a87_t5 ;
reg	[8:0]	rl_a88_t5 ;
reg	[8:0]	rl_a89_t5 ;
reg	[8:0]	rl_a90_t5 ;
reg	[8:0]	rl_a91_t5 ;
reg	[8:0]	rl_a92_t5 ;
reg	[8:0]	rl_a93_t5 ;
reg	[8:0]	rl_a94_t5 ;
reg	[8:0]	rl_a95_t5 ;
reg	[8:0]	rl_a96_t5 ;
reg	[8:0]	rl_a97_t5 ;
reg	[8:0]	rl_a98_t5 ;
reg	[8:0]	rl_a99_t5 ;
reg	[8:0]	rl_a100_t5 ;
reg	[8:0]	rl_a101_t5 ;
reg	[8:0]	rl_a102_t5 ;
reg	[8:0]	rl_a103_t5 ;
reg	[8:0]	rl_a104_t5 ;
reg	[8:0]	rl_a105_t5 ;
reg	[8:0]	rl_a106_t5 ;
reg	[8:0]	rl_a107_t5 ;
reg	[8:0]	rl_a108_t5 ;
reg	[8:0]	rl_a109_t5 ;
reg	[8:0]	rl_a110_t5 ;
reg	[8:0]	rl_a111_t5 ;
reg	[8:0]	rl_a112_t5 ;
reg	[8:0]	rl_a113_t5 ;
reg	[8:0]	rl_a114_t5 ;
reg	[8:0]	rl_a115_t5 ;
reg	[8:0]	rl_a116_t5 ;
reg	[8:0]	rl_a117_t5 ;
reg	[8:0]	rl_a118_t5 ;
reg	[8:0]	rl_a119_t5 ;
reg	[8:0]	rl_a120_t5 ;
reg	[8:0]	rl_a121_t5 ;
reg	[8:0]	rl_a122_t5 ;
reg	[8:0]	rl_a123_t5 ;
reg	[8:0]	rl_a124_t5 ;
reg	[8:0]	rl_a125_t5 ;
reg	[8:0]	rl_a126_t5 ;
reg	[8:0]	rl_a127_t5 ;
reg	RG_M_14_d10_c0_t ;
reg	RG_M_14_d10_c1_t ;
reg	RG_M_14_d10_c2_t ;
reg	RG_M_14_d10_c3_t ;
reg	RG_M_14_d10_c4_t ;
reg	RG_M_14_d10_c5_t ;
reg	RG_M_14_d10_c6_t ;
reg	RG_M_14_d10_c7_t ;
reg	M_14_t128 ;
reg	M_15_t128 ;
reg	[8:0]	RG_rl_t ;
reg	RG_rl_t_c1 ;
reg	[8:0]	RG_rl_t1 ;
reg	[8:0]	RG_rl_1_t ;
reg	RG_rl_1_t_c1 ;
reg	[8:0]	RG_rl_1_t1 ;
reg	[8:0]	RG_rl_2_t ;
reg	RG_rl_2_t_c1 ;
reg	[8:0]	RG_rl_2_t1 ;
reg	[8:0]	RG_rl_3_t ;
reg	RG_rl_3_t_c1 ;
reg	[8:0]	RG_rl_3_t1 ;
reg	[8:0]	RG_rl_4_t ;
reg	RG_rl_4_t_c1 ;
reg	[8:0]	RG_rl_4_t1 ;
reg	[8:0]	RG_rl_5_t ;
reg	RG_rl_5_t_c1 ;
reg	[8:0]	RG_rl_5_t1 ;
reg	[8:0]	RG_rl_6_t ;
reg	RG_rl_6_t_c1 ;
reg	[8:0]	RG_rl_6_t1 ;
reg	[8:0]	RG_rl_7_t ;
reg	RG_rl_7_t_c1 ;
reg	[8:0]	RG_rl_7_t1 ;
reg	[8:0]	RG_rl_8_t ;
reg	RG_rl_8_t_c1 ;
reg	[8:0]	RG_rl_8_t1 ;
reg	[8:0]	RG_rl_9_t ;
reg	RG_rl_9_t_c1 ;
reg	[8:0]	RG_rl_9_t1 ;
reg	[8:0]	RG_rl_10_t ;
reg	RG_rl_10_t_c1 ;
reg	[8:0]	RG_rl_10_t1 ;
reg	[8:0]	RG_rl_11_t ;
reg	RG_rl_11_t_c1 ;
reg	[8:0]	RG_rl_11_t1 ;
reg	[8:0]	RG_rl_12_t ;
reg	RG_rl_12_t_c1 ;
reg	[8:0]	RG_rl_12_t1 ;
reg	[8:0]	RG_rl_13_t ;
reg	RG_rl_13_t_c1 ;
reg	[8:0]	RG_rl_13_t1 ;
reg	[8:0]	RG_rl_14_t ;
reg	RG_rl_14_t_c1 ;
reg	[8:0]	RG_rl_14_t1 ;
reg	[8:0]	RG_rl_15_t ;
reg	RG_rl_15_t_c1 ;
reg	[8:0]	RG_rl_15_t1 ;
reg	[8:0]	RG_rl_16_t ;
reg	RG_rl_16_t_c1 ;
reg	[8:0]	RG_rl_16_t1 ;
reg	[8:0]	RG_rl_17_t ;
reg	RG_rl_17_t_c1 ;
reg	[8:0]	RG_rl_17_t1 ;
reg	[8:0]	RG_rl_18_t ;
reg	RG_rl_18_t_c1 ;
reg	[8:0]	RG_rl_18_t1 ;
reg	[8:0]	RG_rl_19_t ;
reg	RG_rl_19_t_c1 ;
reg	[8:0]	RG_rl_19_t1 ;
reg	[8:0]	RG_rl_20_t ;
reg	RG_rl_20_t_c1 ;
reg	[8:0]	RG_rl_20_t1 ;
reg	[8:0]	RG_rl_21_t ;
reg	RG_rl_21_t_c1 ;
reg	[8:0]	RG_rl_21_t1 ;
reg	[8:0]	RG_rl_22_t ;
reg	RG_rl_22_t_c1 ;
reg	[8:0]	RG_rl_22_t1 ;
reg	[8:0]	RG_rl_23_t ;
reg	RG_rl_23_t_c1 ;
reg	[8:0]	RG_rl_23_t1 ;
reg	[8:0]	RG_rl_24_t ;
reg	RG_rl_24_t_c1 ;
reg	[8:0]	RG_rl_24_t1 ;
reg	[8:0]	RG_rl_25_t ;
reg	RG_rl_25_t_c1 ;
reg	[8:0]	RG_rl_25_t1 ;
reg	[8:0]	RG_rl_26_t ;
reg	RG_rl_26_t_c1 ;
reg	[8:0]	RG_rl_26_t1 ;
reg	[8:0]	RG_rl_27_t ;
reg	RG_rl_27_t_c1 ;
reg	[8:0]	RG_rl_27_t1 ;
reg	[8:0]	RG_rl_28_t ;
reg	RG_rl_28_t_c1 ;
reg	[8:0]	RG_rl_28_t1 ;
reg	[8:0]	RG_rl_29_t ;
reg	RG_rl_29_t_c1 ;
reg	[8:0]	RG_rl_29_t1 ;
reg	[8:0]	RG_rl_30_t ;
reg	RG_rl_30_t_c1 ;
reg	[8:0]	RG_rl_30_t1 ;
reg	[8:0]	RG_rl_31_t ;
reg	RG_rl_31_t_c1 ;
reg	[8:0]	RG_rl_31_t1 ;
reg	[8:0]	RG_rl_32_t ;
reg	RG_rl_32_t_c1 ;
reg	[8:0]	RG_rl_32_t1 ;
reg	[8:0]	RG_rl_33_t ;
reg	RG_rl_33_t_c1 ;
reg	[8:0]	RG_rl_33_t1 ;
reg	[8:0]	RG_rl_34_t ;
reg	RG_rl_34_t_c1 ;
reg	[8:0]	RG_rl_34_t1 ;
reg	[8:0]	RG_rl_35_t ;
reg	RG_rl_35_t_c1 ;
reg	[8:0]	RG_rl_35_t1 ;
reg	[8:0]	RG_rl_36_t ;
reg	RG_rl_36_t_c1 ;
reg	[8:0]	RG_rl_36_t1 ;
reg	[8:0]	RG_rl_37_t ;
reg	RG_rl_37_t_c1 ;
reg	[8:0]	RG_rl_37_t1 ;
reg	[8:0]	RG_rl_38_t ;
reg	RG_rl_38_t_c1 ;
reg	[8:0]	RG_rl_38_t1 ;
reg	[8:0]	RG_rl_39_t ;
reg	RG_rl_39_t_c1 ;
reg	[8:0]	RG_rl_39_t1 ;
reg	[8:0]	RG_rl_40_t ;
reg	RG_rl_40_t_c1 ;
reg	[8:0]	RG_rl_40_t1 ;
reg	[8:0]	RG_rl_41_t ;
reg	RG_rl_41_t_c1 ;
reg	[8:0]	RG_rl_41_t1 ;
reg	[8:0]	RG_rl_42_t ;
reg	RG_rl_42_t_c1 ;
reg	[8:0]	RG_rl_42_t1 ;
reg	[8:0]	RG_rl_43_t ;
reg	RG_rl_43_t_c1 ;
reg	[8:0]	RG_rl_43_t1 ;
reg	[8:0]	RG_rl_44_t ;
reg	RG_rl_44_t_c1 ;
reg	[8:0]	RG_rl_44_t1 ;
reg	[8:0]	RG_rl_45_t ;
reg	RG_rl_45_t_c1 ;
reg	[8:0]	RG_rl_45_t1 ;
reg	[8:0]	RG_rl_46_t ;
reg	RG_rl_46_t_c1 ;
reg	[8:0]	RG_rl_46_t1 ;
reg	[8:0]	RG_rl_47_t ;
reg	RG_rl_47_t_c1 ;
reg	[8:0]	RG_rl_47_t1 ;
reg	[8:0]	RG_rl_48_t ;
reg	RG_rl_48_t_c1 ;
reg	[8:0]	RG_rl_48_t1 ;
reg	[8:0]	RG_rl_49_t ;
reg	RG_rl_49_t_c1 ;
reg	[8:0]	RG_rl_49_t1 ;
reg	[8:0]	RG_rl_50_t ;
reg	RG_rl_50_t_c1 ;
reg	[8:0]	RG_rl_50_t1 ;
reg	[8:0]	RG_rl_51_t ;
reg	RG_rl_51_t_c1 ;
reg	[8:0]	RG_rl_51_t1 ;
reg	[8:0]	RG_rl_52_t ;
reg	RG_rl_52_t_c1 ;
reg	[8:0]	RG_rl_52_t1 ;
reg	[8:0]	RG_rl_53_t ;
reg	RG_rl_53_t_c1 ;
reg	[8:0]	RG_rl_53_t1 ;
reg	[8:0]	RG_rl_54_t ;
reg	RG_rl_54_t_c1 ;
reg	[8:0]	RG_rl_54_t1 ;
reg	[8:0]	RG_rl_55_t ;
reg	RG_rl_55_t_c1 ;
reg	[8:0]	RG_rl_55_t1 ;
reg	[8:0]	RG_rl_56_t ;
reg	RG_rl_56_t_c1 ;
reg	[8:0]	RG_rl_56_t1 ;
reg	[8:0]	RG_rl_57_t ;
reg	RG_rl_57_t_c1 ;
reg	[8:0]	RG_rl_57_t1 ;
reg	[8:0]	RG_rl_58_t ;
reg	RG_rl_58_t_c1 ;
reg	[8:0]	RG_rl_58_t1 ;
reg	[8:0]	RG_rl_59_t ;
reg	RG_rl_59_t_c1 ;
reg	[8:0]	RG_rl_59_t1 ;
reg	[8:0]	RG_rl_60_t ;
reg	RG_rl_60_t_c1 ;
reg	[8:0]	RG_rl_60_t1 ;
reg	[8:0]	RG_rl_61_t ;
reg	RG_rl_61_t_c1 ;
reg	[8:0]	RG_rl_61_t1 ;
reg	[8:0]	RG_rl_62_t ;
reg	RG_rl_62_t_c1 ;
reg	[8:0]	RG_rl_62_t1 ;
reg	[8:0]	RG_rl_63_t ;
reg	RG_rl_63_t_c1 ;
reg	[8:0]	RG_rl_63_t1 ;
reg	[8:0]	RG_rl_64_t ;
reg	RG_rl_64_t_c1 ;
reg	[8:0]	RG_rl_64_t1 ;
reg	[8:0]	RG_rl_65_t ;
reg	RG_rl_65_t_c1 ;
reg	[8:0]	RG_rl_65_t1 ;
reg	[8:0]	RG_rl_66_t ;
reg	RG_rl_66_t_c1 ;
reg	[8:0]	RG_rl_66_t1 ;
reg	[8:0]	RG_rl_67_t ;
reg	RG_rl_67_t_c1 ;
reg	[8:0]	RG_rl_67_t1 ;
reg	[8:0]	RG_rl_68_t ;
reg	RG_rl_68_t_c1 ;
reg	[8:0]	RG_rl_68_t1 ;
reg	[8:0]	RG_rl_69_t ;
reg	RG_rl_69_t_c1 ;
reg	[8:0]	RG_rl_69_t1 ;
reg	[8:0]	RG_rl_70_t ;
reg	RG_rl_70_t_c1 ;
reg	[8:0]	RG_rl_70_t1 ;
reg	[8:0]	RG_rl_71_t ;
reg	RG_rl_71_t_c1 ;
reg	[8:0]	RG_rl_71_t1 ;
reg	[8:0]	RG_rl_72_t ;
reg	RG_rl_72_t_c1 ;
reg	[8:0]	RG_rl_72_t1 ;
reg	[8:0]	RG_rl_73_t ;
reg	RG_rl_73_t_c1 ;
reg	[8:0]	RG_rl_73_t1 ;
reg	[8:0]	RG_rl_74_t ;
reg	RG_rl_74_t_c1 ;
reg	[8:0]	RG_rl_74_t1 ;
reg	[8:0]	RG_rl_75_t ;
reg	RG_rl_75_t_c1 ;
reg	[8:0]	RG_rl_75_t1 ;
reg	[8:0]	RG_rl_76_t ;
reg	RG_rl_76_t_c1 ;
reg	[8:0]	RG_rl_76_t1 ;
reg	[8:0]	RG_rl_77_t ;
reg	RG_rl_77_t_c1 ;
reg	[8:0]	RG_rl_77_t1 ;
reg	[8:0]	RG_rl_78_t ;
reg	RG_rl_78_t_c1 ;
reg	[8:0]	RG_rl_78_t1 ;
reg	[8:0]	RG_rl_79_t ;
reg	RG_rl_79_t_c1 ;
reg	[8:0]	RG_rl_79_t1 ;
reg	[8:0]	RG_rl_80_t ;
reg	RG_rl_80_t_c1 ;
reg	[8:0]	RG_rl_80_t1 ;
reg	[8:0]	RG_rl_81_t ;
reg	RG_rl_81_t_c1 ;
reg	[8:0]	RG_rl_81_t1 ;
reg	[8:0]	RG_rl_82_t ;
reg	RG_rl_82_t_c1 ;
reg	[8:0]	RG_rl_82_t1 ;
reg	[8:0]	RG_rl_83_t ;
reg	RG_rl_83_t_c1 ;
reg	[8:0]	RG_rl_83_t1 ;
reg	[8:0]	RG_rl_84_t ;
reg	RG_rl_84_t_c1 ;
reg	[8:0]	RG_rl_84_t1 ;
reg	[8:0]	RG_rl_85_t ;
reg	RG_rl_85_t_c1 ;
reg	[8:0]	RG_rl_85_t1 ;
reg	[8:0]	RG_rl_86_t ;
reg	RG_rl_86_t_c1 ;
reg	[8:0]	RG_rl_86_t1 ;
reg	[8:0]	RG_rl_87_t ;
reg	RG_rl_87_t_c1 ;
reg	[8:0]	RG_rl_87_t1 ;
reg	[8:0]	RG_rl_88_t ;
reg	RG_rl_88_t_c1 ;
reg	[8:0]	RG_rl_88_t1 ;
reg	[8:0]	RG_rl_89_t ;
reg	RG_rl_89_t_c1 ;
reg	[8:0]	RG_rl_89_t1 ;
reg	[8:0]	RG_rl_90_t ;
reg	RG_rl_90_t_c1 ;
reg	[8:0]	RG_rl_90_t1 ;
reg	[8:0]	RG_rl_91_t ;
reg	RG_rl_91_t_c1 ;
reg	[8:0]	RG_rl_91_t1 ;
reg	[8:0]	RG_rl_92_t ;
reg	RG_rl_92_t_c1 ;
reg	[8:0]	RG_rl_92_t1 ;
reg	[8:0]	RG_rl_93_t ;
reg	RG_rl_93_t_c1 ;
reg	[8:0]	RG_rl_93_t1 ;
reg	[8:0]	RG_rl_94_t ;
reg	RG_rl_94_t_c1 ;
reg	[8:0]	RG_rl_94_t1 ;
reg	[8:0]	RG_rl_95_t ;
reg	RG_rl_95_t_c1 ;
reg	[8:0]	RG_rl_95_t1 ;
reg	[8:0]	RG_rl_96_t ;
reg	RG_rl_96_t_c1 ;
reg	[8:0]	RG_rl_96_t1 ;
reg	[8:0]	RG_rl_97_t ;
reg	RG_rl_97_t_c1 ;
reg	[8:0]	RG_rl_97_t1 ;
reg	[8:0]	RG_rl_98_t ;
reg	RG_rl_98_t_c1 ;
reg	[8:0]	RG_rl_98_t1 ;
reg	[8:0]	RG_rl_99_t ;
reg	RG_rl_99_t_c1 ;
reg	[8:0]	RG_rl_99_t1 ;
reg	[8:0]	RG_rl_100_t ;
reg	RG_rl_100_t_c1 ;
reg	[8:0]	RG_rl_100_t1 ;
reg	[8:0]	RG_rl_101_t ;
reg	RG_rl_101_t_c1 ;
reg	[8:0]	RG_rl_101_t1 ;
reg	[8:0]	RG_rl_102_t ;
reg	RG_rl_102_t_c1 ;
reg	[8:0]	RG_rl_102_t1 ;
reg	[8:0]	RG_rl_103_t ;
reg	RG_rl_103_t_c1 ;
reg	[8:0]	RG_rl_103_t1 ;
reg	[8:0]	RG_rl_104_t ;
reg	RG_rl_104_t_c1 ;
reg	[8:0]	RG_rl_104_t1 ;
reg	[8:0]	RG_rl_105_t ;
reg	RG_rl_105_t_c1 ;
reg	[8:0]	RG_rl_105_t1 ;
reg	[8:0]	RG_rl_106_t ;
reg	RG_rl_106_t_c1 ;
reg	[8:0]	RG_rl_106_t1 ;
reg	[8:0]	RG_rl_107_t ;
reg	RG_rl_107_t_c1 ;
reg	[8:0]	RG_rl_107_t1 ;
reg	[8:0]	RG_rl_108_t ;
reg	RG_rl_108_t_c1 ;
reg	[8:0]	RG_rl_108_t1 ;
reg	[8:0]	RG_rl_109_t ;
reg	RG_rl_109_t_c1 ;
reg	[8:0]	RG_rl_109_t1 ;
reg	[8:0]	RG_rl_110_t ;
reg	RG_rl_110_t_c1 ;
reg	[8:0]	RG_rl_110_t1 ;
reg	[8:0]	RG_rl_111_t ;
reg	RG_rl_111_t_c1 ;
reg	[8:0]	RG_rl_111_t1 ;
reg	[8:0]	RG_rl_112_t ;
reg	RG_rl_112_t_c1 ;
reg	[8:0]	RG_rl_112_t1 ;
reg	[8:0]	RG_rl_113_t ;
reg	RG_rl_113_t_c1 ;
reg	[8:0]	RG_rl_113_t1 ;
reg	[8:0]	RG_rl_114_t ;
reg	RG_rl_114_t_c1 ;
reg	[8:0]	RG_rl_114_t1 ;
reg	[8:0]	RG_rl_115_t ;
reg	RG_rl_115_t_c1 ;
reg	[8:0]	RG_rl_115_t1 ;
reg	[8:0]	RG_rl_116_t ;
reg	RG_rl_116_t_c1 ;
reg	[8:0]	RG_rl_116_t1 ;
reg	[8:0]	RG_rl_117_t ;
reg	RG_rl_117_t_c1 ;
reg	[8:0]	RG_rl_117_t1 ;
reg	[8:0]	RG_rl_118_t ;
reg	RG_rl_118_t_c1 ;
reg	[8:0]	RG_rl_118_t1 ;
reg	[8:0]	RG_rl_119_t ;
reg	RG_rl_119_t_c1 ;
reg	[8:0]	RG_rl_119_t1 ;
reg	[8:0]	RG_rl_120_t ;
reg	RG_rl_120_t_c1 ;
reg	[8:0]	RG_rl_120_t1 ;
reg	[8:0]	RG_rl_121_t ;
reg	RG_rl_121_t_c1 ;
reg	[8:0]	RG_rl_121_t1 ;
reg	[8:0]	RG_rl_122_t ;
reg	RG_rl_122_t_c1 ;
reg	[8:0]	RG_rl_122_t1 ;
reg	[8:0]	RG_rl_123_t ;
reg	RG_rl_123_t_c1 ;
reg	[8:0]	RG_rl_123_t1 ;
reg	[8:0]	RG_rl_124_t ;
reg	RG_rl_124_t_c1 ;
reg	[8:0]	RG_rl_124_t1 ;
reg	[8:0]	RG_rl_125_t ;
reg	RG_rl_125_t_c1 ;
reg	[8:0]	RG_rl_125_t1 ;
reg	[8:0]	RG_rl_126_t ;
reg	RG_rl_126_t_c1 ;
reg	[8:0]	RG_rl_126_t1 ;
reg	[8:0]	RG_rl_127_t ;
reg	RG_rl_127_t_c1 ;
reg	[8:0]	RG_rl_127_t1 ;
reg	[8:0]	RG_rl_184_t ;
reg	RG_rl_184_t_c1 ;
reg	[8:0]	RG_previous_dc_rl_t ;
reg	RG_previous_dc_rl_t_c1 ;
reg	[8:0]	RG_rl_185_t ;
reg	RG_rl_185_t_c1 ;
reg	[8:0]	RG_rl_186_t ;
reg	RG_rl_186_t_c1 ;
reg	[8:0]	RG_rl_187_t ;
reg	RG_rl_187_t_c1 ;
reg	[8:0]	RG_rl_188_t ;
reg	RG_rl_188_t_c1 ;
reg	[8:0]	RG_rl_189_t ;
reg	RG_rl_189_t_c1 ;
reg	[8:0]	RG_rl_190_t ;
reg	RG_rl_190_t_c1 ;
reg	[8:0]	RG_rl_191_t ;
reg	RG_rl_191_t_c1 ;
reg	[8:0]	RG_rl_192_t ;
reg	RG_rl_192_t_c1 ;
reg	[8:0]	RG_rl_193_t ;
reg	RG_rl_193_t_c1 ;
reg	[8:0]	RG_rl_194_t ;
reg	RG_rl_194_t_c1 ;
reg	[8:0]	RG_rl_195_t ;
reg	RG_rl_195_t_c1 ;
reg	[8:0]	RG_rl_196_t ;
reg	RG_rl_196_t_c1 ;
reg	[8:0]	RG_rl_197_t ;
reg	RG_rl_197_t_c1 ;
reg	[8:0]	RG_rl_198_t ;
reg	RG_rl_198_t_c1 ;
reg	[8:0]	RG_rl_199_t ;
reg	RG_rl_199_t_c1 ;
reg	[8:0]	RG_rl_200_t ;
reg	RG_rl_200_t_c1 ;
reg	[8:0]	RG_rl_201_t ;
reg	RG_rl_201_t_c1 ;
reg	[8:0]	RG_rl_202_t ;
reg	RG_rl_202_t_c1 ;
reg	[8:0]	RG_rl_203_t ;
reg	RG_rl_203_t_c1 ;
reg	[8:0]	RG_rl_204_t ;
reg	RG_rl_204_t_c1 ;
reg	[8:0]	RG_rl_205_t ;
reg	RG_rl_205_t_c1 ;
reg	[8:0]	RG_rl_206_t ;
reg	RG_rl_206_t_c1 ;
reg	[8:0]	RG_rl_207_t ;
reg	RG_rl_207_t_c1 ;
reg	[8:0]	RG_rl_208_t ;
reg	RG_rl_208_t_c1 ;
reg	[8:0]	RG_rl_209_t ;
reg	RG_rl_209_t_c1 ;
reg	[8:0]	RG_rl_210_t ;
reg	RG_rl_210_t_c1 ;
reg	[8:0]	RG_rl_211_t ;
reg	RG_rl_211_t_c1 ;
reg	[8:0]	RG_rl_212_t ;
reg	RG_rl_212_t_c1 ;
reg	[8:0]	RG_rl_213_t ;
reg	RG_rl_213_t_c1 ;
reg	[8:0]	RG_rl_214_t ;
reg	RG_rl_214_t_c1 ;
reg	[8:0]	RG_rl_215_t ;
reg	RG_rl_215_t_c1 ;
reg	[8:0]	RG_rl_216_t ;
reg	RG_rl_216_t_c1 ;
reg	[8:0]	RG_rl_217_t ;
reg	RG_rl_217_t_c1 ;
reg	[8:0]	RG_rl_218_t ;
reg	RG_rl_218_t_c1 ;
reg	[8:0]	RG_rl_219_t ;
reg	RG_rl_219_t_c1 ;
reg	[8:0]	RG_rl_220_t ;
reg	RG_rl_220_t_c1 ;
reg	[8:0]	RG_rl_221_t ;
reg	RG_rl_221_t_c1 ;
reg	[8:0]	RG_rl_222_t ;
reg	RG_rl_222_t_c1 ;
reg	[8:0]	RG_rl_223_t ;
reg	RG_rl_223_t_c1 ;
reg	[8:0]	RG_rl_224_t ;
reg	RG_rl_224_t_c1 ;
reg	[8:0]	RG_rl_225_t ;
reg	RG_rl_225_t_c1 ;
reg	[8:0]	RG_rl_226_t ;
reg	RG_rl_226_t_c1 ;
reg	[8:0]	RG_rl_227_t ;
reg	RG_rl_227_t_c1 ;
reg	[8:0]	RG_rl_228_t ;
reg	RG_rl_228_t_c1 ;
reg	[8:0]	RG_rl_229_t ;
reg	RG_rl_229_t_c1 ;
reg	[8:0]	RG_rl_230_t ;
reg	RG_rl_230_t_c1 ;
reg	[8:0]	RG_rl_231_t ;
reg	RG_rl_231_t_c1 ;
reg	[8:0]	RG_rl_232_t ;
reg	RG_rl_232_t_c1 ;
reg	[8:0]	RG_rl_233_t ;
reg	RG_rl_233_t_c1 ;
reg	[8:0]	RG_rl_234_t ;
reg	RG_rl_234_t_c1 ;
reg	[8:0]	RG_rl_235_t ;
reg	RG_rl_235_t_c1 ;
reg	[8:0]	RG_rl_236_t ;
reg	RG_rl_236_t_c1 ;
reg	[8:0]	RG_rl_237_t ;
reg	RG_rl_237_t_c1 ;
reg	[8:0]	RG_rl_238_t ;
reg	RG_rl_238_t_c1 ;
reg	[8:0]	RG_rl_239_t ;
reg	RG_rl_239_t_c1 ;
reg	[8:0]	RG_rl_240_t ;
reg	RG_rl_240_t_c1 ;
reg	[8:0]	RG_rl_241_t ;
reg	RG_rl_241_t_c1 ;
reg	[3:0]	RG_j_t ;
reg	[2:0]	TR_01 ;
reg	[31:0]	RG_i_k_01_t ;
reg	RG_i_k_01_t_c1 ;
reg	RG_i_k_01_t_c2 ;
reg	RG_i_k_01_t_c3 ;
reg	TR_02 ;
reg	[31:0]	RG_i_j_01_t ;
reg	RG_i_j_01_t_c1 ;
reg	RG_i_j_01_t_c2 ;
reg	RG_i_j_01_t_c3 ;
reg	[8:0]	RG_quantized_block_rl_t ;
reg	RG_quantized_block_rl_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_1_t ;
reg	RG_quantized_block_rl_1_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_2_t ;
reg	RG_quantized_block_rl_2_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_3_t ;
reg	RG_quantized_block_rl_3_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_4_t ;
reg	RG_quantized_block_rl_4_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_5_t ;
reg	RG_quantized_block_rl_5_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_6_t ;
reg	RG_quantized_block_rl_6_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_7_t ;
reg	RG_quantized_block_rl_7_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_8_t ;
reg	RG_quantized_block_rl_8_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_9_t ;
reg	RG_quantized_block_rl_9_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_10_t ;
reg	RG_quantized_block_rl_10_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_11_t ;
reg	RG_quantized_block_rl_11_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_12_t ;
reg	RG_quantized_block_rl_12_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_13_t ;
reg	RG_quantized_block_rl_13_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_14_t ;
reg	RG_quantized_block_rl_14_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_15_t ;
reg	RG_quantized_block_rl_15_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_16_t ;
reg	RG_quantized_block_rl_16_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_17_t ;
reg	RG_quantized_block_rl_17_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_18_t ;
reg	RG_quantized_block_rl_18_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_19_t ;
reg	RG_quantized_block_rl_19_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_20_t ;
reg	RG_quantized_block_rl_20_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_21_t ;
reg	RG_quantized_block_rl_21_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_22_t ;
reg	RG_quantized_block_rl_22_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_23_t ;
reg	RG_quantized_block_rl_23_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_24_t ;
reg	RG_quantized_block_rl_24_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_25_t ;
reg	RG_quantized_block_rl_25_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_26_t ;
reg	RG_quantized_block_rl_26_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_27_t ;
reg	RG_quantized_block_rl_27_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_28_t ;
reg	RG_quantized_block_rl_28_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_29_t ;
reg	RG_quantized_block_rl_29_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_30_t ;
reg	RG_quantized_block_rl_30_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_31_t ;
reg	RG_quantized_block_rl_31_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_32_t ;
reg	RG_quantized_block_rl_32_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_33_t ;
reg	RG_quantized_block_rl_33_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_34_t ;
reg	RG_quantized_block_rl_34_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_35_t ;
reg	RG_quantized_block_rl_35_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_36_t ;
reg	RG_quantized_block_rl_36_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_37_t ;
reg	RG_quantized_block_rl_37_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_38_t ;
reg	RG_quantized_block_rl_38_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_39_t ;
reg	RG_quantized_block_rl_39_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_40_t ;
reg	RG_quantized_block_rl_40_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_41_t ;
reg	RG_quantized_block_rl_41_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_42_t ;
reg	RG_quantized_block_rl_42_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_43_t ;
reg	RG_quantized_block_rl_43_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_44_t ;
reg	RG_quantized_block_rl_44_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_45_t ;
reg	RG_quantized_block_rl_45_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_46_t ;
reg	RG_quantized_block_rl_46_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_47_t ;
reg	RG_quantized_block_rl_47_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_48_t ;
reg	RG_quantized_block_rl_48_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_49_t ;
reg	RG_quantized_block_rl_49_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_50_t ;
reg	RG_quantized_block_rl_50_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_51_t ;
reg	RG_quantized_block_rl_51_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_52_t ;
reg	RG_quantized_block_rl_52_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_53_t ;
reg	RG_quantized_block_rl_53_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_54_t ;
reg	RG_quantized_block_rl_54_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_55_t ;
reg	RG_quantized_block_rl_55_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_56_t ;
reg	RG_quantized_block_rl_56_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_57_t ;
reg	RG_quantized_block_rl_57_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_58_t ;
reg	RG_quantized_block_rl_58_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_59_t ;
reg	RG_quantized_block_rl_59_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_60_t ;
reg	RG_quantized_block_rl_60_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_61_t ;
reg	RG_quantized_block_rl_61_t_c1 ;
reg	[8:0]	RG_quantized_block_rl_62_t ;
reg	RG_quantized_block_rl_62_t_c1 ;
reg	[8:0]	RL_previous_dc_quantized_block_t ;
reg	[6:0]	RG_k_01_t ;
reg	RG_k_01_t_c1 ;
reg	FF_d_01_t ;
reg	FF_d_01_t_c1 ;
reg	FF_d_01_t_c2 ;
reg	FF_i_t ;
reg	[8:0]	RG_rl_242_t ;
reg	RG_rl_242_t_c1 ;
reg	[8:0]	RG_rl_243_t ;
reg	RG_rl_243_t_c1 ;
reg	[8:0]	RG_rl_244_t ;
reg	RG_rl_244_t_c1 ;
reg	[8:0]	RG_rl_245_t ;
reg	RG_rl_245_t_c1 ;
reg	[8:0]	RG_rl_246_t ;
reg	RG_rl_246_t_c1 ;
reg	[8:0]	RG_previous_dc_rl_1_t ;
reg	RG_previous_dc_rl_1_t_c1 ;
reg	RG_previous_dc_rl_1_t_c2 ;
reg	[7:0]	RG_len_t ;
reg	FF_len_t ;
reg	[31:0]	i2_t1 ;
reg	i2_t1_c1 ;
reg	[7:0]	len1_t3 ;
reg	len1_t3_c1 ;
reg	[8:0]	rl_a00_t4 ;
reg	rl_a00_t4_c1 ;
reg	[8:0]	rl_a00_t4_t1 ;
reg	[8:0]	rl_a01_t4 ;
reg	rl_a01_t4_c1 ;
reg	[8:0]	rl_a01_t4_t1 ;
reg	[8:0]	rl_a02_t4 ;
reg	rl_a02_t4_c1 ;
reg	[8:0]	rl_a02_t4_t1 ;
reg	[8:0]	rl_a03_t4 ;
reg	rl_a03_t4_c1 ;
reg	[8:0]	rl_a03_t4_t1 ;
reg	[8:0]	rl_a04_t4 ;
reg	rl_a04_t4_c1 ;
reg	[8:0]	rl_a04_t4_t1 ;
reg	[8:0]	rl_a05_t4 ;
reg	rl_a05_t4_c1 ;
reg	[8:0]	rl_a05_t4_t1 ;
reg	[8:0]	rl_a06_t4 ;
reg	rl_a06_t4_c1 ;
reg	[8:0]	rl_a06_t4_t1 ;
reg	[8:0]	rl_a07_t4 ;
reg	rl_a07_t4_c1 ;
reg	[8:0]	rl_a07_t4_t1 ;
reg	[8:0]	rl_a08_t4 ;
reg	rl_a08_t4_c1 ;
reg	[8:0]	rl_a08_t4_t1 ;
reg	[8:0]	rl_a09_t4 ;
reg	rl_a09_t4_c1 ;
reg	[8:0]	rl_a09_t4_t1 ;
reg	[8:0]	rl_a10_t4 ;
reg	rl_a10_t4_c1 ;
reg	[8:0]	rl_a10_t4_t1 ;
reg	[8:0]	rl_a11_t4 ;
reg	rl_a11_t4_c1 ;
reg	[8:0]	rl_a11_t4_t1 ;
reg	[8:0]	rl_a12_t4 ;
reg	rl_a12_t4_c1 ;
reg	[8:0]	rl_a12_t4_t1 ;
reg	[8:0]	rl_a13_t4 ;
reg	rl_a13_t4_c1 ;
reg	[8:0]	rl_a13_t4_t1 ;
reg	[8:0]	rl_a14_t4 ;
reg	rl_a14_t4_c1 ;
reg	[8:0]	rl_a14_t4_t1 ;
reg	[8:0]	rl_a15_t4 ;
reg	rl_a15_t4_c1 ;
reg	[8:0]	rl_a15_t4_t1 ;
reg	[8:0]	rl_a16_t4 ;
reg	rl_a16_t4_c1 ;
reg	[8:0]	rl_a16_t4_t1 ;
reg	[8:0]	rl_a17_t4 ;
reg	rl_a17_t4_c1 ;
reg	[8:0]	rl_a17_t4_t1 ;
reg	[8:0]	rl_a18_t4 ;
reg	rl_a18_t4_c1 ;
reg	[8:0]	rl_a18_t4_t1 ;
reg	[8:0]	rl_a19_t4 ;
reg	rl_a19_t4_c1 ;
reg	[8:0]	rl_a19_t4_t1 ;
reg	[8:0]	rl_a20_t4 ;
reg	rl_a20_t4_c1 ;
reg	[8:0]	rl_a20_t4_t1 ;
reg	[8:0]	rl_a21_t4 ;
reg	rl_a21_t4_c1 ;
reg	[8:0]	rl_a21_t4_t1 ;
reg	[8:0]	rl_a22_t4 ;
reg	rl_a22_t4_c1 ;
reg	[8:0]	rl_a22_t4_t1 ;
reg	[8:0]	rl_a23_t4 ;
reg	rl_a23_t4_c1 ;
reg	[8:0]	rl_a23_t4_t1 ;
reg	[8:0]	rl_a24_t4 ;
reg	rl_a24_t4_c1 ;
reg	[8:0]	rl_a24_t4_t1 ;
reg	[8:0]	rl_a25_t4 ;
reg	rl_a25_t4_c1 ;
reg	[8:0]	rl_a25_t4_t1 ;
reg	[8:0]	rl_a26_t4 ;
reg	rl_a26_t4_c1 ;
reg	[8:0]	rl_a26_t4_t1 ;
reg	[8:0]	rl_a27_t4 ;
reg	rl_a27_t4_c1 ;
reg	[8:0]	rl_a27_t4_t1 ;
reg	[8:0]	rl_a28_t4 ;
reg	rl_a28_t4_c1 ;
reg	[8:0]	rl_a28_t4_t1 ;
reg	[8:0]	rl_a29_t4 ;
reg	rl_a29_t4_c1 ;
reg	[8:0]	rl_a29_t4_t1 ;
reg	[8:0]	rl_a30_t4 ;
reg	rl_a30_t4_c1 ;
reg	[8:0]	rl_a30_t4_t1 ;
reg	[8:0]	rl_a31_t4 ;
reg	rl_a31_t4_c1 ;
reg	[8:0]	rl_a31_t4_t1 ;
reg	[8:0]	rl_a32_t4 ;
reg	rl_a32_t4_c1 ;
reg	[8:0]	rl_a32_t4_t1 ;
reg	[8:0]	rl_a33_t4 ;
reg	rl_a33_t4_c1 ;
reg	[8:0]	rl_a33_t4_t1 ;
reg	[8:0]	rl_a34_t4 ;
reg	rl_a34_t4_c1 ;
reg	[8:0]	rl_a34_t4_t1 ;
reg	[8:0]	rl_a35_t4 ;
reg	rl_a35_t4_c1 ;
reg	[8:0]	rl_a35_t4_t1 ;
reg	[8:0]	rl_a36_t4 ;
reg	rl_a36_t4_c1 ;
reg	[8:0]	rl_a36_t4_t1 ;
reg	[8:0]	rl_a37_t4 ;
reg	rl_a37_t4_c1 ;
reg	[8:0]	rl_a37_t4_t1 ;
reg	[8:0]	rl_a38_t4 ;
reg	rl_a38_t4_c1 ;
reg	[8:0]	rl_a38_t4_t1 ;
reg	[8:0]	rl_a39_t4 ;
reg	rl_a39_t4_c1 ;
reg	[8:0]	rl_a39_t4_t1 ;
reg	[8:0]	rl_a40_t4 ;
reg	rl_a40_t4_c1 ;
reg	[8:0]	rl_a40_t4_t1 ;
reg	[8:0]	rl_a41_t4 ;
reg	rl_a41_t4_c1 ;
reg	[8:0]	rl_a41_t4_t1 ;
reg	[8:0]	rl_a42_t4 ;
reg	rl_a42_t4_c1 ;
reg	[8:0]	rl_a42_t4_t1 ;
reg	[8:0]	rl_a43_t4 ;
reg	rl_a43_t4_c1 ;
reg	[8:0]	rl_a43_t4_t1 ;
reg	[8:0]	rl_a44_t4 ;
reg	rl_a44_t4_c1 ;
reg	[8:0]	rl_a44_t4_t1 ;
reg	[8:0]	rl_a45_t4 ;
reg	rl_a45_t4_c1 ;
reg	[8:0]	rl_a45_t4_t1 ;
reg	[8:0]	rl_a46_t4 ;
reg	rl_a46_t4_c1 ;
reg	[8:0]	rl_a46_t4_t1 ;
reg	[8:0]	rl_a47_t4 ;
reg	rl_a47_t4_c1 ;
reg	[8:0]	rl_a47_t4_t1 ;
reg	[8:0]	rl_a48_t4 ;
reg	rl_a48_t4_c1 ;
reg	[8:0]	rl_a48_t4_t1 ;
reg	[8:0]	rl_a49_t4 ;
reg	rl_a49_t4_c1 ;
reg	[8:0]	rl_a49_t4_t1 ;
reg	[8:0]	rl_a50_t4 ;
reg	rl_a50_t4_c1 ;
reg	[8:0]	rl_a50_t4_t1 ;
reg	[8:0]	rl_a51_t4 ;
reg	rl_a51_t4_c1 ;
reg	[8:0]	rl_a51_t4_t1 ;
reg	[8:0]	rl_a52_t4 ;
reg	rl_a52_t4_c1 ;
reg	[8:0]	rl_a52_t4_t1 ;
reg	[8:0]	rl_a53_t4 ;
reg	rl_a53_t4_c1 ;
reg	[8:0]	rl_a53_t4_t1 ;
reg	[8:0]	rl_a54_t4 ;
reg	rl_a54_t4_c1 ;
reg	[8:0]	rl_a54_t4_t1 ;
reg	[8:0]	rl_a55_t4 ;
reg	rl_a55_t4_c1 ;
reg	[8:0]	rl_a55_t4_t1 ;
reg	[8:0]	rl_a56_t4 ;
reg	rl_a56_t4_c1 ;
reg	[8:0]	rl_a56_t4_t1 ;
reg	[8:0]	rl_a57_t4 ;
reg	rl_a57_t4_c1 ;
reg	[8:0]	rl_a57_t4_t1 ;
reg	[8:0]	rl_a58_t4 ;
reg	rl_a58_t4_c1 ;
reg	[8:0]	rl_a58_t4_t1 ;
reg	[8:0]	rl_a59_t4 ;
reg	rl_a59_t4_c1 ;
reg	[8:0]	rl_a59_t4_t1 ;
reg	[8:0]	rl_a60_t4 ;
reg	rl_a60_t4_c1 ;
reg	[8:0]	rl_a60_t4_t1 ;
reg	[8:0]	rl_a61_t4 ;
reg	rl_a61_t4_c1 ;
reg	[8:0]	rl_a61_t4_t1 ;
reg	[8:0]	rl_a62_t4 ;
reg	rl_a62_t4_c1 ;
reg	[8:0]	rl_a62_t4_t1 ;
reg	[8:0]	rl_a63_t4 ;
reg	rl_a63_t4_c1 ;
reg	[8:0]	rl_a63_t4_t1 ;
reg	[8:0]	rl_a64_t4 ;
reg	rl_a64_t4_c1 ;
reg	[8:0]	rl_a64_t4_t1 ;
reg	[8:0]	rl_a65_t4 ;
reg	rl_a65_t4_c1 ;
reg	[8:0]	rl_a65_t4_t1 ;
reg	[8:0]	rl_a66_t4 ;
reg	rl_a66_t4_c1 ;
reg	[8:0]	rl_a66_t4_t1 ;
reg	[8:0]	rl_a67_t4 ;
reg	rl_a67_t4_c1 ;
reg	[8:0]	rl_a67_t4_t1 ;
reg	[8:0]	rl_a68_t4 ;
reg	rl_a68_t4_c1 ;
reg	[8:0]	rl_a68_t4_t1 ;
reg	[8:0]	rl_a69_t4 ;
reg	rl_a69_t4_c1 ;
reg	[8:0]	rl_a69_t4_t1 ;
reg	[8:0]	rl_a70_t4 ;
reg	rl_a70_t4_c1 ;
reg	[8:0]	rl_a70_t4_t1 ;
reg	[8:0]	rl_a71_t4 ;
reg	rl_a71_t4_c1 ;
reg	[8:0]	rl_a71_t4_t1 ;
reg	[8:0]	rl_a72_t4 ;
reg	rl_a72_t4_c1 ;
reg	[8:0]	rl_a72_t4_t1 ;
reg	[8:0]	rl_a73_t4 ;
reg	rl_a73_t4_c1 ;
reg	[8:0]	rl_a73_t4_t1 ;
reg	[8:0]	rl_a74_t4 ;
reg	rl_a74_t4_c1 ;
reg	[8:0]	rl_a74_t4_t1 ;
reg	[8:0]	rl_a75_t4 ;
reg	rl_a75_t4_c1 ;
reg	[8:0]	rl_a75_t4_t1 ;
reg	[8:0]	rl_a76_t4 ;
reg	rl_a76_t4_c1 ;
reg	[8:0]	rl_a76_t4_t1 ;
reg	[8:0]	rl_a77_t4 ;
reg	rl_a77_t4_c1 ;
reg	[8:0]	rl_a77_t4_t1 ;
reg	[8:0]	rl_a78_t4 ;
reg	rl_a78_t4_c1 ;
reg	[8:0]	rl_a78_t4_t1 ;
reg	[8:0]	rl_a79_t4 ;
reg	rl_a79_t4_c1 ;
reg	[8:0]	rl_a79_t4_t1 ;
reg	[8:0]	rl_a80_t4 ;
reg	rl_a80_t4_c1 ;
reg	[8:0]	rl_a80_t4_t1 ;
reg	[8:0]	rl_a81_t4 ;
reg	rl_a81_t4_c1 ;
reg	[8:0]	rl_a81_t4_t1 ;
reg	[8:0]	rl_a82_t4 ;
reg	rl_a82_t4_c1 ;
reg	[8:0]	rl_a82_t4_t1 ;
reg	[8:0]	rl_a83_t4 ;
reg	rl_a83_t4_c1 ;
reg	[8:0]	rl_a83_t4_t1 ;
reg	[8:0]	rl_a84_t4 ;
reg	rl_a84_t4_c1 ;
reg	[8:0]	rl_a84_t4_t1 ;
reg	[8:0]	rl_a85_t4 ;
reg	rl_a85_t4_c1 ;
reg	[8:0]	rl_a85_t4_t1 ;
reg	[8:0]	rl_a86_t4 ;
reg	rl_a86_t4_c1 ;
reg	[8:0]	rl_a86_t4_t1 ;
reg	[8:0]	rl_a87_t4 ;
reg	rl_a87_t4_c1 ;
reg	[8:0]	rl_a87_t4_t1 ;
reg	[8:0]	rl_a88_t4 ;
reg	rl_a88_t4_c1 ;
reg	[8:0]	rl_a88_t4_t1 ;
reg	[8:0]	rl_a89_t4 ;
reg	rl_a89_t4_c1 ;
reg	[8:0]	rl_a89_t4_t1 ;
reg	[8:0]	rl_a90_t4 ;
reg	rl_a90_t4_c1 ;
reg	[8:0]	rl_a90_t4_t1 ;
reg	[8:0]	rl_a91_t4 ;
reg	rl_a91_t4_c1 ;
reg	[8:0]	rl_a91_t4_t1 ;
reg	[8:0]	rl_a92_t4 ;
reg	rl_a92_t4_c1 ;
reg	[8:0]	rl_a92_t4_t1 ;
reg	[8:0]	rl_a93_t4 ;
reg	rl_a93_t4_c1 ;
reg	[8:0]	rl_a93_t4_t1 ;
reg	[8:0]	rl_a94_t4 ;
reg	rl_a94_t4_c1 ;
reg	[8:0]	rl_a94_t4_t1 ;
reg	[8:0]	rl_a95_t4 ;
reg	rl_a95_t4_c1 ;
reg	[8:0]	rl_a95_t4_t1 ;
reg	[8:0]	rl_a96_t4 ;
reg	rl_a96_t4_c1 ;
reg	[8:0]	rl_a96_t4_t1 ;
reg	[8:0]	rl_a97_t4 ;
reg	rl_a97_t4_c1 ;
reg	[8:0]	rl_a97_t4_t1 ;
reg	[8:0]	rl_a98_t4 ;
reg	rl_a98_t4_c1 ;
reg	[8:0]	rl_a98_t4_t1 ;
reg	[8:0]	rl_a99_t4 ;
reg	rl_a99_t4_c1 ;
reg	[8:0]	rl_a99_t4_t1 ;
reg	[8:0]	rl_a100_t4 ;
reg	rl_a100_t4_c1 ;
reg	[8:0]	rl_a100_t4_t1 ;
reg	[8:0]	rl_a101_t4 ;
reg	rl_a101_t4_c1 ;
reg	[8:0]	rl_a101_t4_t1 ;
reg	[8:0]	rl_a102_t4 ;
reg	rl_a102_t4_c1 ;
reg	[8:0]	rl_a102_t4_t1 ;
reg	[8:0]	rl_a103_t4 ;
reg	rl_a103_t4_c1 ;
reg	[8:0]	rl_a103_t4_t1 ;
reg	[8:0]	rl_a104_t4 ;
reg	rl_a104_t4_c1 ;
reg	[8:0]	rl_a104_t4_t1 ;
reg	[8:0]	rl_a105_t4 ;
reg	rl_a105_t4_c1 ;
reg	[8:0]	rl_a105_t4_t1 ;
reg	[8:0]	rl_a106_t4 ;
reg	rl_a106_t4_c1 ;
reg	[8:0]	rl_a106_t4_t1 ;
reg	[8:0]	rl_a107_t4 ;
reg	rl_a107_t4_c1 ;
reg	[8:0]	rl_a107_t4_t1 ;
reg	[8:0]	rl_a108_t4 ;
reg	rl_a108_t4_c1 ;
reg	[8:0]	rl_a108_t4_t1 ;
reg	[8:0]	rl_a109_t4 ;
reg	rl_a109_t4_c1 ;
reg	[8:0]	rl_a109_t4_t1 ;
reg	[8:0]	rl_a110_t4 ;
reg	rl_a110_t4_c1 ;
reg	[8:0]	rl_a110_t4_t1 ;
reg	[8:0]	rl_a111_t4 ;
reg	rl_a111_t4_c1 ;
reg	[8:0]	rl_a111_t4_t1 ;
reg	[8:0]	rl_a112_t4 ;
reg	rl_a112_t4_c1 ;
reg	[8:0]	rl_a112_t4_t1 ;
reg	[8:0]	rl_a113_t4 ;
reg	rl_a113_t4_c1 ;
reg	[8:0]	rl_a113_t4_t1 ;
reg	[8:0]	rl_a114_t4 ;
reg	rl_a114_t4_c1 ;
reg	[8:0]	rl_a114_t4_t1 ;
reg	[8:0]	rl_a115_t4 ;
reg	rl_a115_t4_c1 ;
reg	[8:0]	rl_a115_t4_t1 ;
reg	[8:0]	rl_a116_t4 ;
reg	rl_a116_t4_c1 ;
reg	[8:0]	rl_a116_t4_t1 ;
reg	[8:0]	rl_a117_t4 ;
reg	rl_a117_t4_c1 ;
reg	[8:0]	rl_a117_t4_t1 ;
reg	[8:0]	rl_a118_t4 ;
reg	rl_a118_t4_c1 ;
reg	[8:0]	rl_a118_t4_t1 ;
reg	[8:0]	rl_a119_t4 ;
reg	rl_a119_t4_c1 ;
reg	[8:0]	rl_a119_t4_t1 ;
reg	[8:0]	rl_a120_t4 ;
reg	rl_a120_t4_c1 ;
reg	[8:0]	rl_a120_t4_t1 ;
reg	[8:0]	rl_a121_t4 ;
reg	rl_a121_t4_c1 ;
reg	[8:0]	rl_a121_t4_t1 ;
reg	[8:0]	rl_a122_t4 ;
reg	rl_a122_t4_c1 ;
reg	[8:0]	rl_a122_t4_t1 ;
reg	[8:0]	rl_a123_t4 ;
reg	rl_a123_t4_c1 ;
reg	[8:0]	rl_a123_t4_t1 ;
reg	[8:0]	rl_a124_t4 ;
reg	rl_a124_t4_c1 ;
reg	[8:0]	rl_a124_t4_t1 ;
reg	[8:0]	rl_a125_t4 ;
reg	rl_a125_t4_c1 ;
reg	[8:0]	rl_a125_t4_t1 ;
reg	[8:0]	rl_a126_t4 ;
reg	rl_a126_t4_c1 ;
reg	[8:0]	rl_a126_t4_t1 ;
reg	[8:0]	rl_a127_t4 ;
reg	rl_a127_t4_c1 ;
reg	[8:0]	rl_a127_t4_t1 ;
reg	M_02_t ;
reg	M_02_t_c1 ;
reg	M_02_t_t1 ;
reg	M_03_t128 ;
reg	M_03_t128_t1 ;
reg	valid_r_t ;
reg	[7:0]	sub8u1i1 ;
reg	sub8u1i1_c1 ;
reg	[7:0]	incr8u3i1 ;
reg	incr8u3i1_c1 ;
reg	incr8u3i1_c2 ;
reg	[5:0]	zz_RA1 ;
reg	zz_RA1_c1 ;
reg	[8:0]	TR_03 ;
reg	[8:0]	TR_04 ;
reg	[8:0]	TR_05 ;
reg	[8:0]	TR_06 ;
reg	[8:0]	TR_07 ;
reg	[8:0]	TR_08 ;
reg	[8:0]	TR_09 ;
reg	[8:0]	TR_10 ;
reg	[8:0]	zz_WD2 ;

jpeg_sub8u_7_1 INST_sub8u_7_1_1 ( .i1(sub8u_7_11i1) ,.i2(sub8u_7_11i2) ,.o1(sub8u_7_11ot) );	// line#=../rle.cpp:83,84
jpeg_sub8u_7 INST_sub8u_7_1 ( .i1(sub8u_71i1) ,.i2(sub8u_71i2) ,.o1(sub8u_71ot) );	// line#=../rle.cpp:83,84
jpeg_decr32s INST_decr32s_1 ( .i1(decr32s1i1) ,.o1(decr32s1ot) );	// line#=../rle.cpp:124,155
jpeg_decr32s INST_decr32s_2 ( .i1(decr32s2i1) ,.o1(decr32s2ot) );	// line#=../rle.cpp:130,161
jpeg_decr8u_7 INST_decr8u_7_1 ( .i1(decr8u_71i1) ,.o1(decr8u_71ot) );	// line#=../rle.cpp:77,78
jpeg_incr32s INST_incr32s_1 ( .i1(incr32s1i1) ,.o1(incr32s1ot) );	// line#=../rle.cpp:64,119,129,150,160
jpeg_incr32s INST_incr32s_2 ( .i1(incr32s2i1) ,.o1(incr32s2ot) );	// line#=../rle.cpp:63,114,125,145,156
jpeg_incr32s INST_incr32s_3 ( .i1(incr32s3i1) ,.o1(incr32s3ot) );	// line#=../rle.cpp:74
jpeg_incr8u INST_incr8u_1 ( .i1(incr8u1i1) ,.o1(incr8u1ot) );	// line#=../rle.cpp:68,73,79
jpeg_incr8u INST_incr8u_2 ( .i1(incr8u2i1) ,.o1(incr8u2ot) );	// line#=../rle.cpp:69
jpeg_incr8u INST_incr8u_3 ( .i1(incr8u3i1) ,.o1(incr8u3ot) );	// line#=../rle.cpp:74,111,142
jpeg_incr8u INST_incr8u_4 ( .i1(incr8u4i1) ,.o1(incr8u4ot) );	// line#=../rle.cpp:80
jpeg_incr4s INST_incr4s_1 ( .i1(incr4s1i1) ,.o1(incr4s1ot) );	// line#=../rle.cpp:34
jpeg_lop8u_1 INST_lop8u_1_1 ( .i1(lop8u_11i1) ,.i2(lop8u_11i2) ,.o1(lop8u_11ot) );	// line#=../rle.cpp:109,110
assign	lop8u_11ot_port = lop8u_11ot ;
jpeg_sub12s_9 INST_sub12s_9_1 ( .i1(sub12s_91i1) ,.i2(sub12s_91i2) ,.o1(sub12s_91ot) );	// line#=../rle.cpp:52
jpeg_sub8u INST_sub8u_1 ( .i1(sub8u1i1) ,.i2(sub8u1i2) ,.o1(sub8u1ot) );	// line#=../rle.cpp:77,78,86
assign	jpeg_out_a00 = jpeg_out_a00_r ;	// line#=../rle.h:60
assign	jpeg_out_a01 = jpeg_out_a01_r ;	// line#=../rle.h:60
assign	jpeg_out_a02 = jpeg_out_a02_r ;	// line#=../rle.h:60
assign	jpeg_out_a03 = jpeg_out_a03_r ;	// line#=../rle.h:60
assign	jpeg_out_a04 = jpeg_out_a04_r ;	// line#=../rle.h:60
assign	jpeg_out_a05 = jpeg_out_a05_r ;	// line#=../rle.h:60
assign	jpeg_out_a06 = jpeg_out_a06_r ;	// line#=../rle.h:60
assign	jpeg_out_a07 = jpeg_out_a07_r ;	// line#=../rle.h:60
assign	jpeg_out_a08 = jpeg_out_a08_r ;	// line#=../rle.h:60
assign	jpeg_out_a09 = jpeg_out_a09_r ;	// line#=../rle.h:60
assign	jpeg_out_a10 = jpeg_out_a10_r ;	// line#=../rle.h:60
assign	jpeg_out_a11 = jpeg_out_a11_r ;	// line#=../rle.h:60
assign	jpeg_out_a12 = jpeg_out_a12_r ;	// line#=../rle.h:60
assign	jpeg_out_a13 = jpeg_out_a13_r ;	// line#=../rle.h:60
assign	jpeg_out_a14 = jpeg_out_a14_r ;	// line#=../rle.h:60
assign	jpeg_out_a15 = jpeg_out_a15_r ;	// line#=../rle.h:60
assign	jpeg_out_a16 = jpeg_out_a16_r ;	// line#=../rle.h:60
assign	jpeg_out_a17 = jpeg_out_a17_r ;	// line#=../rle.h:60
assign	jpeg_out_a18 = jpeg_out_a18_r ;	// line#=../rle.h:60
assign	jpeg_out_a19 = jpeg_out_a19_r ;	// line#=../rle.h:60
assign	jpeg_out_a20 = jpeg_out_a20_r ;	// line#=../rle.h:60
assign	jpeg_out_a21 = jpeg_out_a21_r ;	// line#=../rle.h:60
assign	jpeg_out_a22 = jpeg_out_a22_r ;	// line#=../rle.h:60
assign	jpeg_out_a23 = jpeg_out_a23_r ;	// line#=../rle.h:60
assign	jpeg_out_a24 = jpeg_out_a24_r ;	// line#=../rle.h:60
assign	jpeg_out_a25 = jpeg_out_a25_r ;	// line#=../rle.h:60
assign	jpeg_out_a26 = jpeg_out_a26_r ;	// line#=../rle.h:60
assign	jpeg_out_a27 = jpeg_out_a27_r ;	// line#=../rle.h:60
assign	jpeg_out_a28 = jpeg_out_a28_r ;	// line#=../rle.h:60
assign	jpeg_out_a29 = jpeg_out_a29_r ;	// line#=../rle.h:60
assign	jpeg_out_a30 = jpeg_out_a30_r ;	// line#=../rle.h:60
assign	jpeg_out_a31 = jpeg_out_a31_r ;	// line#=../rle.h:60
assign	jpeg_out_a32 = jpeg_out_a32_r ;	// line#=../rle.h:60
assign	jpeg_out_a33 = jpeg_out_a33_r ;	// line#=../rle.h:60
assign	jpeg_out_a34 = jpeg_out_a34_r ;	// line#=../rle.h:60
assign	jpeg_out_a35 = jpeg_out_a35_r ;	// line#=../rle.h:60
assign	jpeg_out_a36 = jpeg_out_a36_r ;	// line#=../rle.h:60
assign	jpeg_out_a37 = jpeg_out_a37_r ;	// line#=../rle.h:60
assign	jpeg_out_a38 = jpeg_out_a38_r ;	// line#=../rle.h:60
assign	jpeg_out_a39 = jpeg_out_a39_r ;	// line#=../rle.h:60
assign	jpeg_out_a40 = jpeg_out_a40_r ;	// line#=../rle.h:60
assign	jpeg_out_a41 = jpeg_out_a41_r ;	// line#=../rle.h:60
assign	jpeg_out_a42 = jpeg_out_a42_r ;	// line#=../rle.h:60
assign	jpeg_out_a43 = jpeg_out_a43_r ;	// line#=../rle.h:60
assign	jpeg_out_a44 = jpeg_out_a44_r ;	// line#=../rle.h:60
assign	jpeg_out_a45 = jpeg_out_a45_r ;	// line#=../rle.h:60
assign	jpeg_out_a46 = jpeg_out_a46_r ;	// line#=../rle.h:60
assign	jpeg_out_a47 = jpeg_out_a47_r ;	// line#=../rle.h:60
assign	jpeg_out_a48 = jpeg_out_a48_r ;	// line#=../rle.h:60
assign	jpeg_out_a49 = jpeg_out_a49_r ;	// line#=../rle.h:60
assign	jpeg_out_a50 = jpeg_out_a50_r ;	// line#=../rle.h:60
assign	jpeg_out_a51 = jpeg_out_a51_r ;	// line#=../rle.h:60
assign	jpeg_out_a52 = jpeg_out_a52_r ;	// line#=../rle.h:60
assign	jpeg_out_a53 = jpeg_out_a53_r ;	// line#=../rle.h:60
assign	jpeg_out_a54 = jpeg_out_a54_r ;	// line#=../rle.h:60
assign	jpeg_out_a55 = jpeg_out_a55_r ;	// line#=../rle.h:60
assign	jpeg_out_a56 = jpeg_out_a56_r ;	// line#=../rle.h:60
assign	jpeg_out_a57 = jpeg_out_a57_r ;	// line#=../rle.h:60
assign	jpeg_out_a58 = jpeg_out_a58_r ;	// line#=../rle.h:60
assign	jpeg_out_a59 = jpeg_out_a59_r ;	// line#=../rle.h:60
assign	jpeg_out_a60 = jpeg_out_a60_r ;	// line#=../rle.h:60
assign	jpeg_out_a61 = jpeg_out_a61_r ;	// line#=../rle.h:60
assign	jpeg_out_a62 = jpeg_out_a62_r ;	// line#=../rle.h:60
assign	jpeg_out_a63 = jpeg_out_a63_r ;	// line#=../rle.h:60
assign	jpeg_out_a64 = jpeg_out_a64_r ;	// line#=../rle.h:60
assign	jpeg_out_a65 = jpeg_out_a65_r ;	// line#=../rle.h:60
assign	jpeg_out_a66 = jpeg_out_a66_r ;	// line#=../rle.h:60
assign	jpeg_out_a67 = jpeg_out_a67_r ;	// line#=../rle.h:60
assign	jpeg_out_a68 = jpeg_out_a68_r ;	// line#=../rle.h:60
assign	jpeg_out_a69 = jpeg_out_a69_r ;	// line#=../rle.h:60
assign	jpeg_out_a70 = jpeg_out_a70_r ;	// line#=../rle.h:60
assign	jpeg_out_a71 = jpeg_out_a71_r ;	// line#=../rle.h:60
assign	jpeg_out_a72 = jpeg_out_a72_r ;	// line#=../rle.h:60
assign	jpeg_out_a73 = jpeg_out_a73_r ;	// line#=../rle.h:60
assign	jpeg_out_a74 = jpeg_out_a74_r ;	// line#=../rle.h:60
assign	jpeg_out_a75 = jpeg_out_a75_r ;	// line#=../rle.h:60
assign	jpeg_out_a76 = jpeg_out_a76_r ;	// line#=../rle.h:60
assign	jpeg_out_a77 = jpeg_out_a77_r ;	// line#=../rle.h:60
assign	jpeg_out_a78 = jpeg_out_a78_r ;	// line#=../rle.h:60
assign	jpeg_out_a79 = jpeg_out_a79_r ;	// line#=../rle.h:60
assign	jpeg_out_a80 = jpeg_out_a80_r ;	// line#=../rle.h:60
assign	jpeg_out_a81 = jpeg_out_a81_r ;	// line#=../rle.h:60
assign	jpeg_out_a82 = jpeg_out_a82_r ;	// line#=../rle.h:60
assign	jpeg_out_a83 = jpeg_out_a83_r ;	// line#=../rle.h:60
assign	jpeg_out_a84 = jpeg_out_a84_r ;	// line#=../rle.h:60
assign	jpeg_out_a85 = jpeg_out_a85_r ;	// line#=../rle.h:60
assign	jpeg_out_a86 = jpeg_out_a86_r ;	// line#=../rle.h:60
assign	jpeg_out_a87 = jpeg_out_a87_r ;	// line#=../rle.h:60
assign	jpeg_out_a88 = jpeg_out_a88_r ;	// line#=../rle.h:60
assign	jpeg_out_a89 = jpeg_out_a89_r ;	// line#=../rle.h:60
assign	jpeg_out_a90 = jpeg_out_a90_r ;	// line#=../rle.h:60
assign	jpeg_out_a91 = jpeg_out_a91_r ;	// line#=../rle.h:60
assign	jpeg_out_a92 = jpeg_out_a92_r ;	// line#=../rle.h:60
assign	jpeg_out_a93 = jpeg_out_a93_r ;	// line#=../rle.h:60
assign	jpeg_out_a94 = jpeg_out_a94_r ;	// line#=../rle.h:60
assign	jpeg_out_a95 = jpeg_out_a95_r ;	// line#=../rle.h:60
assign	jpeg_out_a96 = jpeg_out_a96_r ;	// line#=../rle.h:60
assign	jpeg_out_a97 = jpeg_out_a97_r ;	// line#=../rle.h:60
assign	jpeg_out_a98 = jpeg_out_a98_r ;	// line#=../rle.h:60
assign	jpeg_out_a99 = jpeg_out_a99_r ;	// line#=../rle.h:60
assign	jpeg_out_a100 = jpeg_out_a100_r ;	// line#=../rle.h:60
assign	jpeg_out_a101 = jpeg_out_a101_r ;	// line#=../rle.h:60
assign	jpeg_out_a102 = jpeg_out_a102_r ;	// line#=../rle.h:60
assign	jpeg_out_a103 = jpeg_out_a103_r ;	// line#=../rle.h:60
assign	jpeg_out_a104 = jpeg_out_a104_r ;	// line#=../rle.h:60
assign	jpeg_out_a105 = jpeg_out_a105_r ;	// line#=../rle.h:60
assign	jpeg_out_a106 = jpeg_out_a106_r ;	// line#=../rle.h:60
assign	jpeg_out_a107 = jpeg_out_a107_r ;	// line#=../rle.h:60
assign	jpeg_out_a108 = jpeg_out_a108_r ;	// line#=../rle.h:60
assign	jpeg_out_a109 = jpeg_out_a109_r ;	// line#=../rle.h:60
assign	jpeg_out_a110 = jpeg_out_a110_r ;	// line#=../rle.h:60
assign	jpeg_out_a111 = jpeg_out_a111_r ;	// line#=../rle.h:60
assign	jpeg_out_a112 = jpeg_out_a112_r ;	// line#=../rle.h:60
assign	jpeg_out_a113 = jpeg_out_a113_r ;	// line#=../rle.h:60
assign	jpeg_out_a114 = jpeg_out_a114_r ;	// line#=../rle.h:60
assign	jpeg_out_a115 = jpeg_out_a115_r ;	// line#=../rle.h:60
assign	jpeg_out_a116 = jpeg_out_a116_r ;	// line#=../rle.h:60
assign	jpeg_out_a117 = jpeg_out_a117_r ;	// line#=../rle.h:60
assign	jpeg_out_a118 = jpeg_out_a118_r ;	// line#=../rle.h:60
assign	jpeg_out_a119 = jpeg_out_a119_r ;	// line#=../rle.h:60
assign	jpeg_out_a120 = jpeg_out_a120_r ;	// line#=../rle.h:60
assign	jpeg_out_a121 = jpeg_out_a121_r ;	// line#=../rle.h:60
assign	jpeg_out_a122 = jpeg_out_a122_r ;	// line#=../rle.h:60
assign	jpeg_out_a123 = jpeg_out_a123_r ;	// line#=../rle.h:60
assign	jpeg_out_a124 = jpeg_out_a124_r ;	// line#=../rle.h:60
assign	jpeg_out_a125 = jpeg_out_a125_r ;	// line#=../rle.h:60
assign	jpeg_out_a126 = jpeg_out_a126_r ;	// line#=../rle.h:60
assign	jpeg_out_a127 = jpeg_out_a127_r ;	// line#=../rle.h:60
assign	jpeg_len_out = jpeg_len_out_r ;	// line#=../rle.h:61
assign	valid = valid_r ;	// line#=../rle.h:62
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_323 <= decr8u_71ot ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_324 <= 1'h0 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_325 <= M_190 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_326 <= M_191 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_327 <= M_192 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_328 <= M_193 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_329 <= M_194 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_330 <= M_195 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_331 <= M_196 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_332 <= M_197 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_333 <= M_198 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_334 <= M_199 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_335 <= M_200 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_336 <= M_201 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_337 <= M_202 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_338 <= M_203 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_339 <= M_204 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_340 <= M_205 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_341 <= M_206 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_342 <= M_207 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_343 <= M_208 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_344 <= M_209 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_345 <= M_210 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_346 <= M_211 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_347 <= M_212 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_348 <= M_213 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_349 <= M_214 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_350 <= M_215 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_351 <= M_216 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_352 <= M_217 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_353 <= M_218 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_354 <= M_219 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_355 <= M_220 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_356 <= M_221 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_357 <= M_222 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_358 <= M_223 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_359 <= M_224 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_360 <= M_225 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_361 <= M_226 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_362 <= M_227 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_363 <= M_228 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_364 <= M_229 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_365 <= M_230 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_366 <= M_231 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_367 <= M_232 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_368 <= M_233 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_369 <= M_234 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_370 <= M_235 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_371 <= M_236 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_372 <= M_237 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_373 <= M_238 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_374 <= M_239 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_375 <= M_240 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_376 <= M_241 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_377 <= M_242 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_378 <= M_243 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_379 <= M_244 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_380 <= M_245 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_381 <= M_246 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_382 <= M_247 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_383 <= M_248 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_384 <= M_249 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_385 <= M_250 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_387 <= M_251 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_388 <= M_252 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_389 <= M_253 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_390 <= M_254 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_391 <= M_255 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_392 <= M_256 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_393 <= M_257 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_394 <= M_258 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_395 <= M_259 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_396 <= M_260 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_397 <= M_261 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_398 <= M_262 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_399 <= M_263 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_400 <= M_264 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_401 <= M_265 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_402 <= M_266 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_403 <= M_267 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_404 <= M_268 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_405 <= M_269 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_406 <= M_270 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_407 <= M_271 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_408 <= M_272 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_409 <= M_273 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_410 <= M_274 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_411 <= M_275 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_412 <= M_276 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_413 <= M_277 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_414 <= M_278 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_415 <= M_279 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_416 <= M_280 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_417 <= M_281 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_418 <= M_282 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_419 <= M_283 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_420 <= M_284 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_421 <= M_285 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_422 <= M_286 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_423 <= M_287 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_424 <= M_288 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_425 <= M_289 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_426 <= M_290 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_427 <= M_291 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_428 <= M_292 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_429 <= M_293 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_430 <= M_294 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_431 <= M_295 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_432 <= M_296 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_433 <= M_297 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_434 <= M_298 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_435 <= M_299 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_436 <= M_300 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_437 <= M_301 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_438 <= M_302 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_439 <= M_303 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_440 <= M_304 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_441 <= M_305 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_442 <= M_306 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_443 <= M_307 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_444 <= M_308 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_445 <= M_309 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_446 <= M_310 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_447 <= M_311 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_448 <= M_312 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_449 <= M_313 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_450 <= M_314 ;
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_451 <= M_315 ;
assign	CT_12 = ( ( ~|RG_i_j_01 ) & M_172 ) ;	// line#=../rle.cpp:117,118
assign	M_172 = ~|{ ( RG_i_k_01 [31] & RG_i_k_01 [0] ) , ~RG_i_k_01 [0] } ;	// line#=../rle.cpp:117,118,140,141,148
										// ,149
assign	CT_17 = ( ( ~|{ RG_i_j_01 [31:3] , ~RG_i_j_01 [2:0] } ) & M_172 ) ;	// line#=../rle.cpp:140,141,148,149
assign	CT_28 = ( RG_i_j_01 [31] | ( ~|RG_i_j_01 [30:6] ) ) ;	// line#=../rle.cpp:61,62
always @ ( zz_RD1 or FF_i )	// line#=../rle.cpp:61,62
	case ( FF_i )
	1'h1 :
		M_01_t1 = ~|zz_RD1 ;	// line#=../rle.cpp:61,62
	1'h0 :
		M_01_t1 = 1'h0 ;	// line#=../rle.cpp:61,62
	default :
		M_01_t1 = 1'hx ;
	endcase
always @ ( RG_rl_184 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_12 = 9'h000 ;	// line#=../rle.cpp:68
	7'h01 :
		TR_12 = RG_rl_184 ;
	7'h02 :
		TR_12 = RG_rl_184 ;
	7'h03 :
		TR_12 = RG_rl_184 ;
	7'h04 :
		TR_12 = RG_rl_184 ;
	7'h05 :
		TR_12 = RG_rl_184 ;
	7'h06 :
		TR_12 = RG_rl_184 ;
	7'h07 :
		TR_12 = RG_rl_184 ;
	7'h08 :
		TR_12 = RG_rl_184 ;
	7'h09 :
		TR_12 = RG_rl_184 ;
	7'h0a :
		TR_12 = RG_rl_184 ;
	7'h0b :
		TR_12 = RG_rl_184 ;
	7'h0c :
		TR_12 = RG_rl_184 ;
	7'h0d :
		TR_12 = RG_rl_184 ;
	7'h0e :
		TR_12 = RG_rl_184 ;
	7'h0f :
		TR_12 = RG_rl_184 ;
	7'h10 :
		TR_12 = RG_rl_184 ;
	7'h11 :
		TR_12 = RG_rl_184 ;
	7'h12 :
		TR_12 = RG_rl_184 ;
	7'h13 :
		TR_12 = RG_rl_184 ;
	7'h14 :
		TR_12 = RG_rl_184 ;
	7'h15 :
		TR_12 = RG_rl_184 ;
	7'h16 :
		TR_12 = RG_rl_184 ;
	7'h17 :
		TR_12 = RG_rl_184 ;
	7'h18 :
		TR_12 = RG_rl_184 ;
	7'h19 :
		TR_12 = RG_rl_184 ;
	7'h1a :
		TR_12 = RG_rl_184 ;
	7'h1b :
		TR_12 = RG_rl_184 ;
	7'h1c :
		TR_12 = RG_rl_184 ;
	7'h1d :
		TR_12 = RG_rl_184 ;
	7'h1e :
		TR_12 = RG_rl_184 ;
	7'h1f :
		TR_12 = RG_rl_184 ;
	7'h20 :
		TR_12 = RG_rl_184 ;
	7'h21 :
		TR_12 = RG_rl_184 ;
	7'h22 :
		TR_12 = RG_rl_184 ;
	7'h23 :
		TR_12 = RG_rl_184 ;
	7'h24 :
		TR_12 = RG_rl_184 ;
	7'h25 :
		TR_12 = RG_rl_184 ;
	7'h26 :
		TR_12 = RG_rl_184 ;
	7'h27 :
		TR_12 = RG_rl_184 ;
	7'h28 :
		TR_12 = RG_rl_184 ;
	7'h29 :
		TR_12 = RG_rl_184 ;
	7'h2a :
		TR_12 = RG_rl_184 ;
	7'h2b :
		TR_12 = RG_rl_184 ;
	7'h2c :
		TR_12 = RG_rl_184 ;
	7'h2d :
		TR_12 = RG_rl_184 ;
	7'h2e :
		TR_12 = RG_rl_184 ;
	7'h2f :
		TR_12 = RG_rl_184 ;
	7'h30 :
		TR_12 = RG_rl_184 ;
	7'h31 :
		TR_12 = RG_rl_184 ;
	7'h32 :
		TR_12 = RG_rl_184 ;
	7'h33 :
		TR_12 = RG_rl_184 ;
	7'h34 :
		TR_12 = RG_rl_184 ;
	7'h35 :
		TR_12 = RG_rl_184 ;
	7'h36 :
		TR_12 = RG_rl_184 ;
	7'h37 :
		TR_12 = RG_rl_184 ;
	7'h38 :
		TR_12 = RG_rl_184 ;
	7'h39 :
		TR_12 = RG_rl_184 ;
	7'h3a :
		TR_12 = RG_rl_184 ;
	7'h3b :
		TR_12 = RG_rl_184 ;
	7'h3c :
		TR_12 = RG_rl_184 ;
	7'h3d :
		TR_12 = RG_rl_184 ;
	7'h3e :
		TR_12 = RG_rl_184 ;
	7'h3f :
		TR_12 = RG_rl_184 ;
	7'h40 :
		TR_12 = RG_rl_184 ;
	7'h41 :
		TR_12 = RG_rl_184 ;
	7'h42 :
		TR_12 = RG_rl_184 ;
	7'h43 :
		TR_12 = RG_rl_184 ;
	7'h44 :
		TR_12 = RG_rl_184 ;
	7'h45 :
		TR_12 = RG_rl_184 ;
	7'h46 :
		TR_12 = RG_rl_184 ;
	7'h47 :
		TR_12 = RG_rl_184 ;
	7'h48 :
		TR_12 = RG_rl_184 ;
	7'h49 :
		TR_12 = RG_rl_184 ;
	7'h4a :
		TR_12 = RG_rl_184 ;
	7'h4b :
		TR_12 = RG_rl_184 ;
	7'h4c :
		TR_12 = RG_rl_184 ;
	7'h4d :
		TR_12 = RG_rl_184 ;
	7'h4e :
		TR_12 = RG_rl_184 ;
	7'h4f :
		TR_12 = RG_rl_184 ;
	7'h50 :
		TR_12 = RG_rl_184 ;
	7'h51 :
		TR_12 = RG_rl_184 ;
	7'h52 :
		TR_12 = RG_rl_184 ;
	7'h53 :
		TR_12 = RG_rl_184 ;
	7'h54 :
		TR_12 = RG_rl_184 ;
	7'h55 :
		TR_12 = RG_rl_184 ;
	7'h56 :
		TR_12 = RG_rl_184 ;
	7'h57 :
		TR_12 = RG_rl_184 ;
	7'h58 :
		TR_12 = RG_rl_184 ;
	7'h59 :
		TR_12 = RG_rl_184 ;
	7'h5a :
		TR_12 = RG_rl_184 ;
	7'h5b :
		TR_12 = RG_rl_184 ;
	7'h5c :
		TR_12 = RG_rl_184 ;
	7'h5d :
		TR_12 = RG_rl_184 ;
	7'h5e :
		TR_12 = RG_rl_184 ;
	7'h5f :
		TR_12 = RG_rl_184 ;
	7'h60 :
		TR_12 = RG_rl_184 ;
	7'h61 :
		TR_12 = RG_rl_184 ;
	7'h62 :
		TR_12 = RG_rl_184 ;
	7'h63 :
		TR_12 = RG_rl_184 ;
	7'h64 :
		TR_12 = RG_rl_184 ;
	7'h65 :
		TR_12 = RG_rl_184 ;
	7'h66 :
		TR_12 = RG_rl_184 ;
	7'h67 :
		TR_12 = RG_rl_184 ;
	7'h68 :
		TR_12 = RG_rl_184 ;
	7'h69 :
		TR_12 = RG_rl_184 ;
	7'h6a :
		TR_12 = RG_rl_184 ;
	7'h6b :
		TR_12 = RG_rl_184 ;
	7'h6c :
		TR_12 = RG_rl_184 ;
	7'h6d :
		TR_12 = RG_rl_184 ;
	7'h6e :
		TR_12 = RG_rl_184 ;
	7'h6f :
		TR_12 = RG_rl_184 ;
	7'h70 :
		TR_12 = RG_rl_184 ;
	7'h71 :
		TR_12 = RG_rl_184 ;
	7'h72 :
		TR_12 = RG_rl_184 ;
	7'h73 :
		TR_12 = RG_rl_184 ;
	7'h74 :
		TR_12 = RG_rl_184 ;
	7'h75 :
		TR_12 = RG_rl_184 ;
	7'h76 :
		TR_12 = RG_rl_184 ;
	7'h77 :
		TR_12 = RG_rl_184 ;
	7'h78 :
		TR_12 = RG_rl_184 ;
	7'h79 :
		TR_12 = RG_rl_184 ;
	7'h7a :
		TR_12 = RG_rl_184 ;
	7'h7b :
		TR_12 = RG_rl_184 ;
	7'h7c :
		TR_12 = RG_rl_184 ;
	7'h7d :
		TR_12 = RG_rl_184 ;
	7'h7e :
		TR_12 = RG_rl_184 ;
	7'h7f :
		TR_12 = RG_rl_184 ;
	default :
		TR_12 = 9'hx ;
	endcase
always @ ( RG_previous_dc_rl or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_13 = RG_previous_dc_rl ;
	7'h01 :
		TR_13 = 9'h000 ;	// line#=../rle.cpp:68
	7'h02 :
		TR_13 = RG_previous_dc_rl ;
	7'h03 :
		TR_13 = RG_previous_dc_rl ;
	7'h04 :
		TR_13 = RG_previous_dc_rl ;
	7'h05 :
		TR_13 = RG_previous_dc_rl ;
	7'h06 :
		TR_13 = RG_previous_dc_rl ;
	7'h07 :
		TR_13 = RG_previous_dc_rl ;
	7'h08 :
		TR_13 = RG_previous_dc_rl ;
	7'h09 :
		TR_13 = RG_previous_dc_rl ;
	7'h0a :
		TR_13 = RG_previous_dc_rl ;
	7'h0b :
		TR_13 = RG_previous_dc_rl ;
	7'h0c :
		TR_13 = RG_previous_dc_rl ;
	7'h0d :
		TR_13 = RG_previous_dc_rl ;
	7'h0e :
		TR_13 = RG_previous_dc_rl ;
	7'h0f :
		TR_13 = RG_previous_dc_rl ;
	7'h10 :
		TR_13 = RG_previous_dc_rl ;
	7'h11 :
		TR_13 = RG_previous_dc_rl ;
	7'h12 :
		TR_13 = RG_previous_dc_rl ;
	7'h13 :
		TR_13 = RG_previous_dc_rl ;
	7'h14 :
		TR_13 = RG_previous_dc_rl ;
	7'h15 :
		TR_13 = RG_previous_dc_rl ;
	7'h16 :
		TR_13 = RG_previous_dc_rl ;
	7'h17 :
		TR_13 = RG_previous_dc_rl ;
	7'h18 :
		TR_13 = RG_previous_dc_rl ;
	7'h19 :
		TR_13 = RG_previous_dc_rl ;
	7'h1a :
		TR_13 = RG_previous_dc_rl ;
	7'h1b :
		TR_13 = RG_previous_dc_rl ;
	7'h1c :
		TR_13 = RG_previous_dc_rl ;
	7'h1d :
		TR_13 = RG_previous_dc_rl ;
	7'h1e :
		TR_13 = RG_previous_dc_rl ;
	7'h1f :
		TR_13 = RG_previous_dc_rl ;
	7'h20 :
		TR_13 = RG_previous_dc_rl ;
	7'h21 :
		TR_13 = RG_previous_dc_rl ;
	7'h22 :
		TR_13 = RG_previous_dc_rl ;
	7'h23 :
		TR_13 = RG_previous_dc_rl ;
	7'h24 :
		TR_13 = RG_previous_dc_rl ;
	7'h25 :
		TR_13 = RG_previous_dc_rl ;
	7'h26 :
		TR_13 = RG_previous_dc_rl ;
	7'h27 :
		TR_13 = RG_previous_dc_rl ;
	7'h28 :
		TR_13 = RG_previous_dc_rl ;
	7'h29 :
		TR_13 = RG_previous_dc_rl ;
	7'h2a :
		TR_13 = RG_previous_dc_rl ;
	7'h2b :
		TR_13 = RG_previous_dc_rl ;
	7'h2c :
		TR_13 = RG_previous_dc_rl ;
	7'h2d :
		TR_13 = RG_previous_dc_rl ;
	7'h2e :
		TR_13 = RG_previous_dc_rl ;
	7'h2f :
		TR_13 = RG_previous_dc_rl ;
	7'h30 :
		TR_13 = RG_previous_dc_rl ;
	7'h31 :
		TR_13 = RG_previous_dc_rl ;
	7'h32 :
		TR_13 = RG_previous_dc_rl ;
	7'h33 :
		TR_13 = RG_previous_dc_rl ;
	7'h34 :
		TR_13 = RG_previous_dc_rl ;
	7'h35 :
		TR_13 = RG_previous_dc_rl ;
	7'h36 :
		TR_13 = RG_previous_dc_rl ;
	7'h37 :
		TR_13 = RG_previous_dc_rl ;
	7'h38 :
		TR_13 = RG_previous_dc_rl ;
	7'h39 :
		TR_13 = RG_previous_dc_rl ;
	7'h3a :
		TR_13 = RG_previous_dc_rl ;
	7'h3b :
		TR_13 = RG_previous_dc_rl ;
	7'h3c :
		TR_13 = RG_previous_dc_rl ;
	7'h3d :
		TR_13 = RG_previous_dc_rl ;
	7'h3e :
		TR_13 = RG_previous_dc_rl ;
	7'h3f :
		TR_13 = RG_previous_dc_rl ;
	7'h40 :
		TR_13 = RG_previous_dc_rl ;
	7'h41 :
		TR_13 = RG_previous_dc_rl ;
	7'h42 :
		TR_13 = RG_previous_dc_rl ;
	7'h43 :
		TR_13 = RG_previous_dc_rl ;
	7'h44 :
		TR_13 = RG_previous_dc_rl ;
	7'h45 :
		TR_13 = RG_previous_dc_rl ;
	7'h46 :
		TR_13 = RG_previous_dc_rl ;
	7'h47 :
		TR_13 = RG_previous_dc_rl ;
	7'h48 :
		TR_13 = RG_previous_dc_rl ;
	7'h49 :
		TR_13 = RG_previous_dc_rl ;
	7'h4a :
		TR_13 = RG_previous_dc_rl ;
	7'h4b :
		TR_13 = RG_previous_dc_rl ;
	7'h4c :
		TR_13 = RG_previous_dc_rl ;
	7'h4d :
		TR_13 = RG_previous_dc_rl ;
	7'h4e :
		TR_13 = RG_previous_dc_rl ;
	7'h4f :
		TR_13 = RG_previous_dc_rl ;
	7'h50 :
		TR_13 = RG_previous_dc_rl ;
	7'h51 :
		TR_13 = RG_previous_dc_rl ;
	7'h52 :
		TR_13 = RG_previous_dc_rl ;
	7'h53 :
		TR_13 = RG_previous_dc_rl ;
	7'h54 :
		TR_13 = RG_previous_dc_rl ;
	7'h55 :
		TR_13 = RG_previous_dc_rl ;
	7'h56 :
		TR_13 = RG_previous_dc_rl ;
	7'h57 :
		TR_13 = RG_previous_dc_rl ;
	7'h58 :
		TR_13 = RG_previous_dc_rl ;
	7'h59 :
		TR_13 = RG_previous_dc_rl ;
	7'h5a :
		TR_13 = RG_previous_dc_rl ;
	7'h5b :
		TR_13 = RG_previous_dc_rl ;
	7'h5c :
		TR_13 = RG_previous_dc_rl ;
	7'h5d :
		TR_13 = RG_previous_dc_rl ;
	7'h5e :
		TR_13 = RG_previous_dc_rl ;
	7'h5f :
		TR_13 = RG_previous_dc_rl ;
	7'h60 :
		TR_13 = RG_previous_dc_rl ;
	7'h61 :
		TR_13 = RG_previous_dc_rl ;
	7'h62 :
		TR_13 = RG_previous_dc_rl ;
	7'h63 :
		TR_13 = RG_previous_dc_rl ;
	7'h64 :
		TR_13 = RG_previous_dc_rl ;
	7'h65 :
		TR_13 = RG_previous_dc_rl ;
	7'h66 :
		TR_13 = RG_previous_dc_rl ;
	7'h67 :
		TR_13 = RG_previous_dc_rl ;
	7'h68 :
		TR_13 = RG_previous_dc_rl ;
	7'h69 :
		TR_13 = RG_previous_dc_rl ;
	7'h6a :
		TR_13 = RG_previous_dc_rl ;
	7'h6b :
		TR_13 = RG_previous_dc_rl ;
	7'h6c :
		TR_13 = RG_previous_dc_rl ;
	7'h6d :
		TR_13 = RG_previous_dc_rl ;
	7'h6e :
		TR_13 = RG_previous_dc_rl ;
	7'h6f :
		TR_13 = RG_previous_dc_rl ;
	7'h70 :
		TR_13 = RG_previous_dc_rl ;
	7'h71 :
		TR_13 = RG_previous_dc_rl ;
	7'h72 :
		TR_13 = RG_previous_dc_rl ;
	7'h73 :
		TR_13 = RG_previous_dc_rl ;
	7'h74 :
		TR_13 = RG_previous_dc_rl ;
	7'h75 :
		TR_13 = RG_previous_dc_rl ;
	7'h76 :
		TR_13 = RG_previous_dc_rl ;
	7'h77 :
		TR_13 = RG_previous_dc_rl ;
	7'h78 :
		TR_13 = RG_previous_dc_rl ;
	7'h79 :
		TR_13 = RG_previous_dc_rl ;
	7'h7a :
		TR_13 = RG_previous_dc_rl ;
	7'h7b :
		TR_13 = RG_previous_dc_rl ;
	7'h7c :
		TR_13 = RG_previous_dc_rl ;
	7'h7d :
		TR_13 = RG_previous_dc_rl ;
	7'h7e :
		TR_13 = RG_previous_dc_rl ;
	7'h7f :
		TR_13 = RG_previous_dc_rl ;
	default :
		TR_13 = 9'hx ;
	endcase
always @ ( RG_rl_185 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_14 = RG_rl_185 ;
	7'h01 :
		TR_14 = RG_rl_185 ;
	7'h02 :
		TR_14 = 9'h000 ;	// line#=../rle.cpp:68
	7'h03 :
		TR_14 = RG_rl_185 ;
	7'h04 :
		TR_14 = RG_rl_185 ;
	7'h05 :
		TR_14 = RG_rl_185 ;
	7'h06 :
		TR_14 = RG_rl_185 ;
	7'h07 :
		TR_14 = RG_rl_185 ;
	7'h08 :
		TR_14 = RG_rl_185 ;
	7'h09 :
		TR_14 = RG_rl_185 ;
	7'h0a :
		TR_14 = RG_rl_185 ;
	7'h0b :
		TR_14 = RG_rl_185 ;
	7'h0c :
		TR_14 = RG_rl_185 ;
	7'h0d :
		TR_14 = RG_rl_185 ;
	7'h0e :
		TR_14 = RG_rl_185 ;
	7'h0f :
		TR_14 = RG_rl_185 ;
	7'h10 :
		TR_14 = RG_rl_185 ;
	7'h11 :
		TR_14 = RG_rl_185 ;
	7'h12 :
		TR_14 = RG_rl_185 ;
	7'h13 :
		TR_14 = RG_rl_185 ;
	7'h14 :
		TR_14 = RG_rl_185 ;
	7'h15 :
		TR_14 = RG_rl_185 ;
	7'h16 :
		TR_14 = RG_rl_185 ;
	7'h17 :
		TR_14 = RG_rl_185 ;
	7'h18 :
		TR_14 = RG_rl_185 ;
	7'h19 :
		TR_14 = RG_rl_185 ;
	7'h1a :
		TR_14 = RG_rl_185 ;
	7'h1b :
		TR_14 = RG_rl_185 ;
	7'h1c :
		TR_14 = RG_rl_185 ;
	7'h1d :
		TR_14 = RG_rl_185 ;
	7'h1e :
		TR_14 = RG_rl_185 ;
	7'h1f :
		TR_14 = RG_rl_185 ;
	7'h20 :
		TR_14 = RG_rl_185 ;
	7'h21 :
		TR_14 = RG_rl_185 ;
	7'h22 :
		TR_14 = RG_rl_185 ;
	7'h23 :
		TR_14 = RG_rl_185 ;
	7'h24 :
		TR_14 = RG_rl_185 ;
	7'h25 :
		TR_14 = RG_rl_185 ;
	7'h26 :
		TR_14 = RG_rl_185 ;
	7'h27 :
		TR_14 = RG_rl_185 ;
	7'h28 :
		TR_14 = RG_rl_185 ;
	7'h29 :
		TR_14 = RG_rl_185 ;
	7'h2a :
		TR_14 = RG_rl_185 ;
	7'h2b :
		TR_14 = RG_rl_185 ;
	7'h2c :
		TR_14 = RG_rl_185 ;
	7'h2d :
		TR_14 = RG_rl_185 ;
	7'h2e :
		TR_14 = RG_rl_185 ;
	7'h2f :
		TR_14 = RG_rl_185 ;
	7'h30 :
		TR_14 = RG_rl_185 ;
	7'h31 :
		TR_14 = RG_rl_185 ;
	7'h32 :
		TR_14 = RG_rl_185 ;
	7'h33 :
		TR_14 = RG_rl_185 ;
	7'h34 :
		TR_14 = RG_rl_185 ;
	7'h35 :
		TR_14 = RG_rl_185 ;
	7'h36 :
		TR_14 = RG_rl_185 ;
	7'h37 :
		TR_14 = RG_rl_185 ;
	7'h38 :
		TR_14 = RG_rl_185 ;
	7'h39 :
		TR_14 = RG_rl_185 ;
	7'h3a :
		TR_14 = RG_rl_185 ;
	7'h3b :
		TR_14 = RG_rl_185 ;
	7'h3c :
		TR_14 = RG_rl_185 ;
	7'h3d :
		TR_14 = RG_rl_185 ;
	7'h3e :
		TR_14 = RG_rl_185 ;
	7'h3f :
		TR_14 = RG_rl_185 ;
	7'h40 :
		TR_14 = RG_rl_185 ;
	7'h41 :
		TR_14 = RG_rl_185 ;
	7'h42 :
		TR_14 = RG_rl_185 ;
	7'h43 :
		TR_14 = RG_rl_185 ;
	7'h44 :
		TR_14 = RG_rl_185 ;
	7'h45 :
		TR_14 = RG_rl_185 ;
	7'h46 :
		TR_14 = RG_rl_185 ;
	7'h47 :
		TR_14 = RG_rl_185 ;
	7'h48 :
		TR_14 = RG_rl_185 ;
	7'h49 :
		TR_14 = RG_rl_185 ;
	7'h4a :
		TR_14 = RG_rl_185 ;
	7'h4b :
		TR_14 = RG_rl_185 ;
	7'h4c :
		TR_14 = RG_rl_185 ;
	7'h4d :
		TR_14 = RG_rl_185 ;
	7'h4e :
		TR_14 = RG_rl_185 ;
	7'h4f :
		TR_14 = RG_rl_185 ;
	7'h50 :
		TR_14 = RG_rl_185 ;
	7'h51 :
		TR_14 = RG_rl_185 ;
	7'h52 :
		TR_14 = RG_rl_185 ;
	7'h53 :
		TR_14 = RG_rl_185 ;
	7'h54 :
		TR_14 = RG_rl_185 ;
	7'h55 :
		TR_14 = RG_rl_185 ;
	7'h56 :
		TR_14 = RG_rl_185 ;
	7'h57 :
		TR_14 = RG_rl_185 ;
	7'h58 :
		TR_14 = RG_rl_185 ;
	7'h59 :
		TR_14 = RG_rl_185 ;
	7'h5a :
		TR_14 = RG_rl_185 ;
	7'h5b :
		TR_14 = RG_rl_185 ;
	7'h5c :
		TR_14 = RG_rl_185 ;
	7'h5d :
		TR_14 = RG_rl_185 ;
	7'h5e :
		TR_14 = RG_rl_185 ;
	7'h5f :
		TR_14 = RG_rl_185 ;
	7'h60 :
		TR_14 = RG_rl_185 ;
	7'h61 :
		TR_14 = RG_rl_185 ;
	7'h62 :
		TR_14 = RG_rl_185 ;
	7'h63 :
		TR_14 = RG_rl_185 ;
	7'h64 :
		TR_14 = RG_rl_185 ;
	7'h65 :
		TR_14 = RG_rl_185 ;
	7'h66 :
		TR_14 = RG_rl_185 ;
	7'h67 :
		TR_14 = RG_rl_185 ;
	7'h68 :
		TR_14 = RG_rl_185 ;
	7'h69 :
		TR_14 = RG_rl_185 ;
	7'h6a :
		TR_14 = RG_rl_185 ;
	7'h6b :
		TR_14 = RG_rl_185 ;
	7'h6c :
		TR_14 = RG_rl_185 ;
	7'h6d :
		TR_14 = RG_rl_185 ;
	7'h6e :
		TR_14 = RG_rl_185 ;
	7'h6f :
		TR_14 = RG_rl_185 ;
	7'h70 :
		TR_14 = RG_rl_185 ;
	7'h71 :
		TR_14 = RG_rl_185 ;
	7'h72 :
		TR_14 = RG_rl_185 ;
	7'h73 :
		TR_14 = RG_rl_185 ;
	7'h74 :
		TR_14 = RG_rl_185 ;
	7'h75 :
		TR_14 = RG_rl_185 ;
	7'h76 :
		TR_14 = RG_rl_185 ;
	7'h77 :
		TR_14 = RG_rl_185 ;
	7'h78 :
		TR_14 = RG_rl_185 ;
	7'h79 :
		TR_14 = RG_rl_185 ;
	7'h7a :
		TR_14 = RG_rl_185 ;
	7'h7b :
		TR_14 = RG_rl_185 ;
	7'h7c :
		TR_14 = RG_rl_185 ;
	7'h7d :
		TR_14 = RG_rl_185 ;
	7'h7e :
		TR_14 = RG_rl_185 ;
	7'h7f :
		TR_14 = RG_rl_185 ;
	default :
		TR_14 = 9'hx ;
	endcase
always @ ( RG_rl_186 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_15 = RG_rl_186 ;
	7'h01 :
		TR_15 = RG_rl_186 ;
	7'h02 :
		TR_15 = RG_rl_186 ;
	7'h03 :
		TR_15 = 9'h000 ;	// line#=../rle.cpp:68
	7'h04 :
		TR_15 = RG_rl_186 ;
	7'h05 :
		TR_15 = RG_rl_186 ;
	7'h06 :
		TR_15 = RG_rl_186 ;
	7'h07 :
		TR_15 = RG_rl_186 ;
	7'h08 :
		TR_15 = RG_rl_186 ;
	7'h09 :
		TR_15 = RG_rl_186 ;
	7'h0a :
		TR_15 = RG_rl_186 ;
	7'h0b :
		TR_15 = RG_rl_186 ;
	7'h0c :
		TR_15 = RG_rl_186 ;
	7'h0d :
		TR_15 = RG_rl_186 ;
	7'h0e :
		TR_15 = RG_rl_186 ;
	7'h0f :
		TR_15 = RG_rl_186 ;
	7'h10 :
		TR_15 = RG_rl_186 ;
	7'h11 :
		TR_15 = RG_rl_186 ;
	7'h12 :
		TR_15 = RG_rl_186 ;
	7'h13 :
		TR_15 = RG_rl_186 ;
	7'h14 :
		TR_15 = RG_rl_186 ;
	7'h15 :
		TR_15 = RG_rl_186 ;
	7'h16 :
		TR_15 = RG_rl_186 ;
	7'h17 :
		TR_15 = RG_rl_186 ;
	7'h18 :
		TR_15 = RG_rl_186 ;
	7'h19 :
		TR_15 = RG_rl_186 ;
	7'h1a :
		TR_15 = RG_rl_186 ;
	7'h1b :
		TR_15 = RG_rl_186 ;
	7'h1c :
		TR_15 = RG_rl_186 ;
	7'h1d :
		TR_15 = RG_rl_186 ;
	7'h1e :
		TR_15 = RG_rl_186 ;
	7'h1f :
		TR_15 = RG_rl_186 ;
	7'h20 :
		TR_15 = RG_rl_186 ;
	7'h21 :
		TR_15 = RG_rl_186 ;
	7'h22 :
		TR_15 = RG_rl_186 ;
	7'h23 :
		TR_15 = RG_rl_186 ;
	7'h24 :
		TR_15 = RG_rl_186 ;
	7'h25 :
		TR_15 = RG_rl_186 ;
	7'h26 :
		TR_15 = RG_rl_186 ;
	7'h27 :
		TR_15 = RG_rl_186 ;
	7'h28 :
		TR_15 = RG_rl_186 ;
	7'h29 :
		TR_15 = RG_rl_186 ;
	7'h2a :
		TR_15 = RG_rl_186 ;
	7'h2b :
		TR_15 = RG_rl_186 ;
	7'h2c :
		TR_15 = RG_rl_186 ;
	7'h2d :
		TR_15 = RG_rl_186 ;
	7'h2e :
		TR_15 = RG_rl_186 ;
	7'h2f :
		TR_15 = RG_rl_186 ;
	7'h30 :
		TR_15 = RG_rl_186 ;
	7'h31 :
		TR_15 = RG_rl_186 ;
	7'h32 :
		TR_15 = RG_rl_186 ;
	7'h33 :
		TR_15 = RG_rl_186 ;
	7'h34 :
		TR_15 = RG_rl_186 ;
	7'h35 :
		TR_15 = RG_rl_186 ;
	7'h36 :
		TR_15 = RG_rl_186 ;
	7'h37 :
		TR_15 = RG_rl_186 ;
	7'h38 :
		TR_15 = RG_rl_186 ;
	7'h39 :
		TR_15 = RG_rl_186 ;
	7'h3a :
		TR_15 = RG_rl_186 ;
	7'h3b :
		TR_15 = RG_rl_186 ;
	7'h3c :
		TR_15 = RG_rl_186 ;
	7'h3d :
		TR_15 = RG_rl_186 ;
	7'h3e :
		TR_15 = RG_rl_186 ;
	7'h3f :
		TR_15 = RG_rl_186 ;
	7'h40 :
		TR_15 = RG_rl_186 ;
	7'h41 :
		TR_15 = RG_rl_186 ;
	7'h42 :
		TR_15 = RG_rl_186 ;
	7'h43 :
		TR_15 = RG_rl_186 ;
	7'h44 :
		TR_15 = RG_rl_186 ;
	7'h45 :
		TR_15 = RG_rl_186 ;
	7'h46 :
		TR_15 = RG_rl_186 ;
	7'h47 :
		TR_15 = RG_rl_186 ;
	7'h48 :
		TR_15 = RG_rl_186 ;
	7'h49 :
		TR_15 = RG_rl_186 ;
	7'h4a :
		TR_15 = RG_rl_186 ;
	7'h4b :
		TR_15 = RG_rl_186 ;
	7'h4c :
		TR_15 = RG_rl_186 ;
	7'h4d :
		TR_15 = RG_rl_186 ;
	7'h4e :
		TR_15 = RG_rl_186 ;
	7'h4f :
		TR_15 = RG_rl_186 ;
	7'h50 :
		TR_15 = RG_rl_186 ;
	7'h51 :
		TR_15 = RG_rl_186 ;
	7'h52 :
		TR_15 = RG_rl_186 ;
	7'h53 :
		TR_15 = RG_rl_186 ;
	7'h54 :
		TR_15 = RG_rl_186 ;
	7'h55 :
		TR_15 = RG_rl_186 ;
	7'h56 :
		TR_15 = RG_rl_186 ;
	7'h57 :
		TR_15 = RG_rl_186 ;
	7'h58 :
		TR_15 = RG_rl_186 ;
	7'h59 :
		TR_15 = RG_rl_186 ;
	7'h5a :
		TR_15 = RG_rl_186 ;
	7'h5b :
		TR_15 = RG_rl_186 ;
	7'h5c :
		TR_15 = RG_rl_186 ;
	7'h5d :
		TR_15 = RG_rl_186 ;
	7'h5e :
		TR_15 = RG_rl_186 ;
	7'h5f :
		TR_15 = RG_rl_186 ;
	7'h60 :
		TR_15 = RG_rl_186 ;
	7'h61 :
		TR_15 = RG_rl_186 ;
	7'h62 :
		TR_15 = RG_rl_186 ;
	7'h63 :
		TR_15 = RG_rl_186 ;
	7'h64 :
		TR_15 = RG_rl_186 ;
	7'h65 :
		TR_15 = RG_rl_186 ;
	7'h66 :
		TR_15 = RG_rl_186 ;
	7'h67 :
		TR_15 = RG_rl_186 ;
	7'h68 :
		TR_15 = RG_rl_186 ;
	7'h69 :
		TR_15 = RG_rl_186 ;
	7'h6a :
		TR_15 = RG_rl_186 ;
	7'h6b :
		TR_15 = RG_rl_186 ;
	7'h6c :
		TR_15 = RG_rl_186 ;
	7'h6d :
		TR_15 = RG_rl_186 ;
	7'h6e :
		TR_15 = RG_rl_186 ;
	7'h6f :
		TR_15 = RG_rl_186 ;
	7'h70 :
		TR_15 = RG_rl_186 ;
	7'h71 :
		TR_15 = RG_rl_186 ;
	7'h72 :
		TR_15 = RG_rl_186 ;
	7'h73 :
		TR_15 = RG_rl_186 ;
	7'h74 :
		TR_15 = RG_rl_186 ;
	7'h75 :
		TR_15 = RG_rl_186 ;
	7'h76 :
		TR_15 = RG_rl_186 ;
	7'h77 :
		TR_15 = RG_rl_186 ;
	7'h78 :
		TR_15 = RG_rl_186 ;
	7'h79 :
		TR_15 = RG_rl_186 ;
	7'h7a :
		TR_15 = RG_rl_186 ;
	7'h7b :
		TR_15 = RG_rl_186 ;
	7'h7c :
		TR_15 = RG_rl_186 ;
	7'h7d :
		TR_15 = RG_rl_186 ;
	7'h7e :
		TR_15 = RG_rl_186 ;
	7'h7f :
		TR_15 = RG_rl_186 ;
	default :
		TR_15 = 9'hx ;
	endcase
always @ ( RG_rl_187 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_16 = RG_rl_187 ;
	7'h01 :
		TR_16 = RG_rl_187 ;
	7'h02 :
		TR_16 = RG_rl_187 ;
	7'h03 :
		TR_16 = RG_rl_187 ;
	7'h04 :
		TR_16 = 9'h000 ;	// line#=../rle.cpp:68
	7'h05 :
		TR_16 = RG_rl_187 ;
	7'h06 :
		TR_16 = RG_rl_187 ;
	7'h07 :
		TR_16 = RG_rl_187 ;
	7'h08 :
		TR_16 = RG_rl_187 ;
	7'h09 :
		TR_16 = RG_rl_187 ;
	7'h0a :
		TR_16 = RG_rl_187 ;
	7'h0b :
		TR_16 = RG_rl_187 ;
	7'h0c :
		TR_16 = RG_rl_187 ;
	7'h0d :
		TR_16 = RG_rl_187 ;
	7'h0e :
		TR_16 = RG_rl_187 ;
	7'h0f :
		TR_16 = RG_rl_187 ;
	7'h10 :
		TR_16 = RG_rl_187 ;
	7'h11 :
		TR_16 = RG_rl_187 ;
	7'h12 :
		TR_16 = RG_rl_187 ;
	7'h13 :
		TR_16 = RG_rl_187 ;
	7'h14 :
		TR_16 = RG_rl_187 ;
	7'h15 :
		TR_16 = RG_rl_187 ;
	7'h16 :
		TR_16 = RG_rl_187 ;
	7'h17 :
		TR_16 = RG_rl_187 ;
	7'h18 :
		TR_16 = RG_rl_187 ;
	7'h19 :
		TR_16 = RG_rl_187 ;
	7'h1a :
		TR_16 = RG_rl_187 ;
	7'h1b :
		TR_16 = RG_rl_187 ;
	7'h1c :
		TR_16 = RG_rl_187 ;
	7'h1d :
		TR_16 = RG_rl_187 ;
	7'h1e :
		TR_16 = RG_rl_187 ;
	7'h1f :
		TR_16 = RG_rl_187 ;
	7'h20 :
		TR_16 = RG_rl_187 ;
	7'h21 :
		TR_16 = RG_rl_187 ;
	7'h22 :
		TR_16 = RG_rl_187 ;
	7'h23 :
		TR_16 = RG_rl_187 ;
	7'h24 :
		TR_16 = RG_rl_187 ;
	7'h25 :
		TR_16 = RG_rl_187 ;
	7'h26 :
		TR_16 = RG_rl_187 ;
	7'h27 :
		TR_16 = RG_rl_187 ;
	7'h28 :
		TR_16 = RG_rl_187 ;
	7'h29 :
		TR_16 = RG_rl_187 ;
	7'h2a :
		TR_16 = RG_rl_187 ;
	7'h2b :
		TR_16 = RG_rl_187 ;
	7'h2c :
		TR_16 = RG_rl_187 ;
	7'h2d :
		TR_16 = RG_rl_187 ;
	7'h2e :
		TR_16 = RG_rl_187 ;
	7'h2f :
		TR_16 = RG_rl_187 ;
	7'h30 :
		TR_16 = RG_rl_187 ;
	7'h31 :
		TR_16 = RG_rl_187 ;
	7'h32 :
		TR_16 = RG_rl_187 ;
	7'h33 :
		TR_16 = RG_rl_187 ;
	7'h34 :
		TR_16 = RG_rl_187 ;
	7'h35 :
		TR_16 = RG_rl_187 ;
	7'h36 :
		TR_16 = RG_rl_187 ;
	7'h37 :
		TR_16 = RG_rl_187 ;
	7'h38 :
		TR_16 = RG_rl_187 ;
	7'h39 :
		TR_16 = RG_rl_187 ;
	7'h3a :
		TR_16 = RG_rl_187 ;
	7'h3b :
		TR_16 = RG_rl_187 ;
	7'h3c :
		TR_16 = RG_rl_187 ;
	7'h3d :
		TR_16 = RG_rl_187 ;
	7'h3e :
		TR_16 = RG_rl_187 ;
	7'h3f :
		TR_16 = RG_rl_187 ;
	7'h40 :
		TR_16 = RG_rl_187 ;
	7'h41 :
		TR_16 = RG_rl_187 ;
	7'h42 :
		TR_16 = RG_rl_187 ;
	7'h43 :
		TR_16 = RG_rl_187 ;
	7'h44 :
		TR_16 = RG_rl_187 ;
	7'h45 :
		TR_16 = RG_rl_187 ;
	7'h46 :
		TR_16 = RG_rl_187 ;
	7'h47 :
		TR_16 = RG_rl_187 ;
	7'h48 :
		TR_16 = RG_rl_187 ;
	7'h49 :
		TR_16 = RG_rl_187 ;
	7'h4a :
		TR_16 = RG_rl_187 ;
	7'h4b :
		TR_16 = RG_rl_187 ;
	7'h4c :
		TR_16 = RG_rl_187 ;
	7'h4d :
		TR_16 = RG_rl_187 ;
	7'h4e :
		TR_16 = RG_rl_187 ;
	7'h4f :
		TR_16 = RG_rl_187 ;
	7'h50 :
		TR_16 = RG_rl_187 ;
	7'h51 :
		TR_16 = RG_rl_187 ;
	7'h52 :
		TR_16 = RG_rl_187 ;
	7'h53 :
		TR_16 = RG_rl_187 ;
	7'h54 :
		TR_16 = RG_rl_187 ;
	7'h55 :
		TR_16 = RG_rl_187 ;
	7'h56 :
		TR_16 = RG_rl_187 ;
	7'h57 :
		TR_16 = RG_rl_187 ;
	7'h58 :
		TR_16 = RG_rl_187 ;
	7'h59 :
		TR_16 = RG_rl_187 ;
	7'h5a :
		TR_16 = RG_rl_187 ;
	7'h5b :
		TR_16 = RG_rl_187 ;
	7'h5c :
		TR_16 = RG_rl_187 ;
	7'h5d :
		TR_16 = RG_rl_187 ;
	7'h5e :
		TR_16 = RG_rl_187 ;
	7'h5f :
		TR_16 = RG_rl_187 ;
	7'h60 :
		TR_16 = RG_rl_187 ;
	7'h61 :
		TR_16 = RG_rl_187 ;
	7'h62 :
		TR_16 = RG_rl_187 ;
	7'h63 :
		TR_16 = RG_rl_187 ;
	7'h64 :
		TR_16 = RG_rl_187 ;
	7'h65 :
		TR_16 = RG_rl_187 ;
	7'h66 :
		TR_16 = RG_rl_187 ;
	7'h67 :
		TR_16 = RG_rl_187 ;
	7'h68 :
		TR_16 = RG_rl_187 ;
	7'h69 :
		TR_16 = RG_rl_187 ;
	7'h6a :
		TR_16 = RG_rl_187 ;
	7'h6b :
		TR_16 = RG_rl_187 ;
	7'h6c :
		TR_16 = RG_rl_187 ;
	7'h6d :
		TR_16 = RG_rl_187 ;
	7'h6e :
		TR_16 = RG_rl_187 ;
	7'h6f :
		TR_16 = RG_rl_187 ;
	7'h70 :
		TR_16 = RG_rl_187 ;
	7'h71 :
		TR_16 = RG_rl_187 ;
	7'h72 :
		TR_16 = RG_rl_187 ;
	7'h73 :
		TR_16 = RG_rl_187 ;
	7'h74 :
		TR_16 = RG_rl_187 ;
	7'h75 :
		TR_16 = RG_rl_187 ;
	7'h76 :
		TR_16 = RG_rl_187 ;
	7'h77 :
		TR_16 = RG_rl_187 ;
	7'h78 :
		TR_16 = RG_rl_187 ;
	7'h79 :
		TR_16 = RG_rl_187 ;
	7'h7a :
		TR_16 = RG_rl_187 ;
	7'h7b :
		TR_16 = RG_rl_187 ;
	7'h7c :
		TR_16 = RG_rl_187 ;
	7'h7d :
		TR_16 = RG_rl_187 ;
	7'h7e :
		TR_16 = RG_rl_187 ;
	7'h7f :
		TR_16 = RG_rl_187 ;
	default :
		TR_16 = 9'hx ;
	endcase
always @ ( RG_rl_188 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_17 = RG_rl_188 ;
	7'h01 :
		TR_17 = RG_rl_188 ;
	7'h02 :
		TR_17 = RG_rl_188 ;
	7'h03 :
		TR_17 = RG_rl_188 ;
	7'h04 :
		TR_17 = RG_rl_188 ;
	7'h05 :
		TR_17 = 9'h000 ;	// line#=../rle.cpp:68
	7'h06 :
		TR_17 = RG_rl_188 ;
	7'h07 :
		TR_17 = RG_rl_188 ;
	7'h08 :
		TR_17 = RG_rl_188 ;
	7'h09 :
		TR_17 = RG_rl_188 ;
	7'h0a :
		TR_17 = RG_rl_188 ;
	7'h0b :
		TR_17 = RG_rl_188 ;
	7'h0c :
		TR_17 = RG_rl_188 ;
	7'h0d :
		TR_17 = RG_rl_188 ;
	7'h0e :
		TR_17 = RG_rl_188 ;
	7'h0f :
		TR_17 = RG_rl_188 ;
	7'h10 :
		TR_17 = RG_rl_188 ;
	7'h11 :
		TR_17 = RG_rl_188 ;
	7'h12 :
		TR_17 = RG_rl_188 ;
	7'h13 :
		TR_17 = RG_rl_188 ;
	7'h14 :
		TR_17 = RG_rl_188 ;
	7'h15 :
		TR_17 = RG_rl_188 ;
	7'h16 :
		TR_17 = RG_rl_188 ;
	7'h17 :
		TR_17 = RG_rl_188 ;
	7'h18 :
		TR_17 = RG_rl_188 ;
	7'h19 :
		TR_17 = RG_rl_188 ;
	7'h1a :
		TR_17 = RG_rl_188 ;
	7'h1b :
		TR_17 = RG_rl_188 ;
	7'h1c :
		TR_17 = RG_rl_188 ;
	7'h1d :
		TR_17 = RG_rl_188 ;
	7'h1e :
		TR_17 = RG_rl_188 ;
	7'h1f :
		TR_17 = RG_rl_188 ;
	7'h20 :
		TR_17 = RG_rl_188 ;
	7'h21 :
		TR_17 = RG_rl_188 ;
	7'h22 :
		TR_17 = RG_rl_188 ;
	7'h23 :
		TR_17 = RG_rl_188 ;
	7'h24 :
		TR_17 = RG_rl_188 ;
	7'h25 :
		TR_17 = RG_rl_188 ;
	7'h26 :
		TR_17 = RG_rl_188 ;
	7'h27 :
		TR_17 = RG_rl_188 ;
	7'h28 :
		TR_17 = RG_rl_188 ;
	7'h29 :
		TR_17 = RG_rl_188 ;
	7'h2a :
		TR_17 = RG_rl_188 ;
	7'h2b :
		TR_17 = RG_rl_188 ;
	7'h2c :
		TR_17 = RG_rl_188 ;
	7'h2d :
		TR_17 = RG_rl_188 ;
	7'h2e :
		TR_17 = RG_rl_188 ;
	7'h2f :
		TR_17 = RG_rl_188 ;
	7'h30 :
		TR_17 = RG_rl_188 ;
	7'h31 :
		TR_17 = RG_rl_188 ;
	7'h32 :
		TR_17 = RG_rl_188 ;
	7'h33 :
		TR_17 = RG_rl_188 ;
	7'h34 :
		TR_17 = RG_rl_188 ;
	7'h35 :
		TR_17 = RG_rl_188 ;
	7'h36 :
		TR_17 = RG_rl_188 ;
	7'h37 :
		TR_17 = RG_rl_188 ;
	7'h38 :
		TR_17 = RG_rl_188 ;
	7'h39 :
		TR_17 = RG_rl_188 ;
	7'h3a :
		TR_17 = RG_rl_188 ;
	7'h3b :
		TR_17 = RG_rl_188 ;
	7'h3c :
		TR_17 = RG_rl_188 ;
	7'h3d :
		TR_17 = RG_rl_188 ;
	7'h3e :
		TR_17 = RG_rl_188 ;
	7'h3f :
		TR_17 = RG_rl_188 ;
	7'h40 :
		TR_17 = RG_rl_188 ;
	7'h41 :
		TR_17 = RG_rl_188 ;
	7'h42 :
		TR_17 = RG_rl_188 ;
	7'h43 :
		TR_17 = RG_rl_188 ;
	7'h44 :
		TR_17 = RG_rl_188 ;
	7'h45 :
		TR_17 = RG_rl_188 ;
	7'h46 :
		TR_17 = RG_rl_188 ;
	7'h47 :
		TR_17 = RG_rl_188 ;
	7'h48 :
		TR_17 = RG_rl_188 ;
	7'h49 :
		TR_17 = RG_rl_188 ;
	7'h4a :
		TR_17 = RG_rl_188 ;
	7'h4b :
		TR_17 = RG_rl_188 ;
	7'h4c :
		TR_17 = RG_rl_188 ;
	7'h4d :
		TR_17 = RG_rl_188 ;
	7'h4e :
		TR_17 = RG_rl_188 ;
	7'h4f :
		TR_17 = RG_rl_188 ;
	7'h50 :
		TR_17 = RG_rl_188 ;
	7'h51 :
		TR_17 = RG_rl_188 ;
	7'h52 :
		TR_17 = RG_rl_188 ;
	7'h53 :
		TR_17 = RG_rl_188 ;
	7'h54 :
		TR_17 = RG_rl_188 ;
	7'h55 :
		TR_17 = RG_rl_188 ;
	7'h56 :
		TR_17 = RG_rl_188 ;
	7'h57 :
		TR_17 = RG_rl_188 ;
	7'h58 :
		TR_17 = RG_rl_188 ;
	7'h59 :
		TR_17 = RG_rl_188 ;
	7'h5a :
		TR_17 = RG_rl_188 ;
	7'h5b :
		TR_17 = RG_rl_188 ;
	7'h5c :
		TR_17 = RG_rl_188 ;
	7'h5d :
		TR_17 = RG_rl_188 ;
	7'h5e :
		TR_17 = RG_rl_188 ;
	7'h5f :
		TR_17 = RG_rl_188 ;
	7'h60 :
		TR_17 = RG_rl_188 ;
	7'h61 :
		TR_17 = RG_rl_188 ;
	7'h62 :
		TR_17 = RG_rl_188 ;
	7'h63 :
		TR_17 = RG_rl_188 ;
	7'h64 :
		TR_17 = RG_rl_188 ;
	7'h65 :
		TR_17 = RG_rl_188 ;
	7'h66 :
		TR_17 = RG_rl_188 ;
	7'h67 :
		TR_17 = RG_rl_188 ;
	7'h68 :
		TR_17 = RG_rl_188 ;
	7'h69 :
		TR_17 = RG_rl_188 ;
	7'h6a :
		TR_17 = RG_rl_188 ;
	7'h6b :
		TR_17 = RG_rl_188 ;
	7'h6c :
		TR_17 = RG_rl_188 ;
	7'h6d :
		TR_17 = RG_rl_188 ;
	7'h6e :
		TR_17 = RG_rl_188 ;
	7'h6f :
		TR_17 = RG_rl_188 ;
	7'h70 :
		TR_17 = RG_rl_188 ;
	7'h71 :
		TR_17 = RG_rl_188 ;
	7'h72 :
		TR_17 = RG_rl_188 ;
	7'h73 :
		TR_17 = RG_rl_188 ;
	7'h74 :
		TR_17 = RG_rl_188 ;
	7'h75 :
		TR_17 = RG_rl_188 ;
	7'h76 :
		TR_17 = RG_rl_188 ;
	7'h77 :
		TR_17 = RG_rl_188 ;
	7'h78 :
		TR_17 = RG_rl_188 ;
	7'h79 :
		TR_17 = RG_rl_188 ;
	7'h7a :
		TR_17 = RG_rl_188 ;
	7'h7b :
		TR_17 = RG_rl_188 ;
	7'h7c :
		TR_17 = RG_rl_188 ;
	7'h7d :
		TR_17 = RG_rl_188 ;
	7'h7e :
		TR_17 = RG_rl_188 ;
	7'h7f :
		TR_17 = RG_rl_188 ;
	default :
		TR_17 = 9'hx ;
	endcase
always @ ( RG_rl_189 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_18 = RG_rl_189 ;
	7'h01 :
		TR_18 = RG_rl_189 ;
	7'h02 :
		TR_18 = RG_rl_189 ;
	7'h03 :
		TR_18 = RG_rl_189 ;
	7'h04 :
		TR_18 = RG_rl_189 ;
	7'h05 :
		TR_18 = RG_rl_189 ;
	7'h06 :
		TR_18 = 9'h000 ;	// line#=../rle.cpp:68
	7'h07 :
		TR_18 = RG_rl_189 ;
	7'h08 :
		TR_18 = RG_rl_189 ;
	7'h09 :
		TR_18 = RG_rl_189 ;
	7'h0a :
		TR_18 = RG_rl_189 ;
	7'h0b :
		TR_18 = RG_rl_189 ;
	7'h0c :
		TR_18 = RG_rl_189 ;
	7'h0d :
		TR_18 = RG_rl_189 ;
	7'h0e :
		TR_18 = RG_rl_189 ;
	7'h0f :
		TR_18 = RG_rl_189 ;
	7'h10 :
		TR_18 = RG_rl_189 ;
	7'h11 :
		TR_18 = RG_rl_189 ;
	7'h12 :
		TR_18 = RG_rl_189 ;
	7'h13 :
		TR_18 = RG_rl_189 ;
	7'h14 :
		TR_18 = RG_rl_189 ;
	7'h15 :
		TR_18 = RG_rl_189 ;
	7'h16 :
		TR_18 = RG_rl_189 ;
	7'h17 :
		TR_18 = RG_rl_189 ;
	7'h18 :
		TR_18 = RG_rl_189 ;
	7'h19 :
		TR_18 = RG_rl_189 ;
	7'h1a :
		TR_18 = RG_rl_189 ;
	7'h1b :
		TR_18 = RG_rl_189 ;
	7'h1c :
		TR_18 = RG_rl_189 ;
	7'h1d :
		TR_18 = RG_rl_189 ;
	7'h1e :
		TR_18 = RG_rl_189 ;
	7'h1f :
		TR_18 = RG_rl_189 ;
	7'h20 :
		TR_18 = RG_rl_189 ;
	7'h21 :
		TR_18 = RG_rl_189 ;
	7'h22 :
		TR_18 = RG_rl_189 ;
	7'h23 :
		TR_18 = RG_rl_189 ;
	7'h24 :
		TR_18 = RG_rl_189 ;
	7'h25 :
		TR_18 = RG_rl_189 ;
	7'h26 :
		TR_18 = RG_rl_189 ;
	7'h27 :
		TR_18 = RG_rl_189 ;
	7'h28 :
		TR_18 = RG_rl_189 ;
	7'h29 :
		TR_18 = RG_rl_189 ;
	7'h2a :
		TR_18 = RG_rl_189 ;
	7'h2b :
		TR_18 = RG_rl_189 ;
	7'h2c :
		TR_18 = RG_rl_189 ;
	7'h2d :
		TR_18 = RG_rl_189 ;
	7'h2e :
		TR_18 = RG_rl_189 ;
	7'h2f :
		TR_18 = RG_rl_189 ;
	7'h30 :
		TR_18 = RG_rl_189 ;
	7'h31 :
		TR_18 = RG_rl_189 ;
	7'h32 :
		TR_18 = RG_rl_189 ;
	7'h33 :
		TR_18 = RG_rl_189 ;
	7'h34 :
		TR_18 = RG_rl_189 ;
	7'h35 :
		TR_18 = RG_rl_189 ;
	7'h36 :
		TR_18 = RG_rl_189 ;
	7'h37 :
		TR_18 = RG_rl_189 ;
	7'h38 :
		TR_18 = RG_rl_189 ;
	7'h39 :
		TR_18 = RG_rl_189 ;
	7'h3a :
		TR_18 = RG_rl_189 ;
	7'h3b :
		TR_18 = RG_rl_189 ;
	7'h3c :
		TR_18 = RG_rl_189 ;
	7'h3d :
		TR_18 = RG_rl_189 ;
	7'h3e :
		TR_18 = RG_rl_189 ;
	7'h3f :
		TR_18 = RG_rl_189 ;
	7'h40 :
		TR_18 = RG_rl_189 ;
	7'h41 :
		TR_18 = RG_rl_189 ;
	7'h42 :
		TR_18 = RG_rl_189 ;
	7'h43 :
		TR_18 = RG_rl_189 ;
	7'h44 :
		TR_18 = RG_rl_189 ;
	7'h45 :
		TR_18 = RG_rl_189 ;
	7'h46 :
		TR_18 = RG_rl_189 ;
	7'h47 :
		TR_18 = RG_rl_189 ;
	7'h48 :
		TR_18 = RG_rl_189 ;
	7'h49 :
		TR_18 = RG_rl_189 ;
	7'h4a :
		TR_18 = RG_rl_189 ;
	7'h4b :
		TR_18 = RG_rl_189 ;
	7'h4c :
		TR_18 = RG_rl_189 ;
	7'h4d :
		TR_18 = RG_rl_189 ;
	7'h4e :
		TR_18 = RG_rl_189 ;
	7'h4f :
		TR_18 = RG_rl_189 ;
	7'h50 :
		TR_18 = RG_rl_189 ;
	7'h51 :
		TR_18 = RG_rl_189 ;
	7'h52 :
		TR_18 = RG_rl_189 ;
	7'h53 :
		TR_18 = RG_rl_189 ;
	7'h54 :
		TR_18 = RG_rl_189 ;
	7'h55 :
		TR_18 = RG_rl_189 ;
	7'h56 :
		TR_18 = RG_rl_189 ;
	7'h57 :
		TR_18 = RG_rl_189 ;
	7'h58 :
		TR_18 = RG_rl_189 ;
	7'h59 :
		TR_18 = RG_rl_189 ;
	7'h5a :
		TR_18 = RG_rl_189 ;
	7'h5b :
		TR_18 = RG_rl_189 ;
	7'h5c :
		TR_18 = RG_rl_189 ;
	7'h5d :
		TR_18 = RG_rl_189 ;
	7'h5e :
		TR_18 = RG_rl_189 ;
	7'h5f :
		TR_18 = RG_rl_189 ;
	7'h60 :
		TR_18 = RG_rl_189 ;
	7'h61 :
		TR_18 = RG_rl_189 ;
	7'h62 :
		TR_18 = RG_rl_189 ;
	7'h63 :
		TR_18 = RG_rl_189 ;
	7'h64 :
		TR_18 = RG_rl_189 ;
	7'h65 :
		TR_18 = RG_rl_189 ;
	7'h66 :
		TR_18 = RG_rl_189 ;
	7'h67 :
		TR_18 = RG_rl_189 ;
	7'h68 :
		TR_18 = RG_rl_189 ;
	7'h69 :
		TR_18 = RG_rl_189 ;
	7'h6a :
		TR_18 = RG_rl_189 ;
	7'h6b :
		TR_18 = RG_rl_189 ;
	7'h6c :
		TR_18 = RG_rl_189 ;
	7'h6d :
		TR_18 = RG_rl_189 ;
	7'h6e :
		TR_18 = RG_rl_189 ;
	7'h6f :
		TR_18 = RG_rl_189 ;
	7'h70 :
		TR_18 = RG_rl_189 ;
	7'h71 :
		TR_18 = RG_rl_189 ;
	7'h72 :
		TR_18 = RG_rl_189 ;
	7'h73 :
		TR_18 = RG_rl_189 ;
	7'h74 :
		TR_18 = RG_rl_189 ;
	7'h75 :
		TR_18 = RG_rl_189 ;
	7'h76 :
		TR_18 = RG_rl_189 ;
	7'h77 :
		TR_18 = RG_rl_189 ;
	7'h78 :
		TR_18 = RG_rl_189 ;
	7'h79 :
		TR_18 = RG_rl_189 ;
	7'h7a :
		TR_18 = RG_rl_189 ;
	7'h7b :
		TR_18 = RG_rl_189 ;
	7'h7c :
		TR_18 = RG_rl_189 ;
	7'h7d :
		TR_18 = RG_rl_189 ;
	7'h7e :
		TR_18 = RG_rl_189 ;
	7'h7f :
		TR_18 = RG_rl_189 ;
	default :
		TR_18 = 9'hx ;
	endcase
always @ ( RG_rl_190 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_19 = RG_rl_190 ;
	7'h01 :
		TR_19 = RG_rl_190 ;
	7'h02 :
		TR_19 = RG_rl_190 ;
	7'h03 :
		TR_19 = RG_rl_190 ;
	7'h04 :
		TR_19 = RG_rl_190 ;
	7'h05 :
		TR_19 = RG_rl_190 ;
	7'h06 :
		TR_19 = RG_rl_190 ;
	7'h07 :
		TR_19 = 9'h000 ;	// line#=../rle.cpp:68
	7'h08 :
		TR_19 = RG_rl_190 ;
	7'h09 :
		TR_19 = RG_rl_190 ;
	7'h0a :
		TR_19 = RG_rl_190 ;
	7'h0b :
		TR_19 = RG_rl_190 ;
	7'h0c :
		TR_19 = RG_rl_190 ;
	7'h0d :
		TR_19 = RG_rl_190 ;
	7'h0e :
		TR_19 = RG_rl_190 ;
	7'h0f :
		TR_19 = RG_rl_190 ;
	7'h10 :
		TR_19 = RG_rl_190 ;
	7'h11 :
		TR_19 = RG_rl_190 ;
	7'h12 :
		TR_19 = RG_rl_190 ;
	7'h13 :
		TR_19 = RG_rl_190 ;
	7'h14 :
		TR_19 = RG_rl_190 ;
	7'h15 :
		TR_19 = RG_rl_190 ;
	7'h16 :
		TR_19 = RG_rl_190 ;
	7'h17 :
		TR_19 = RG_rl_190 ;
	7'h18 :
		TR_19 = RG_rl_190 ;
	7'h19 :
		TR_19 = RG_rl_190 ;
	7'h1a :
		TR_19 = RG_rl_190 ;
	7'h1b :
		TR_19 = RG_rl_190 ;
	7'h1c :
		TR_19 = RG_rl_190 ;
	7'h1d :
		TR_19 = RG_rl_190 ;
	7'h1e :
		TR_19 = RG_rl_190 ;
	7'h1f :
		TR_19 = RG_rl_190 ;
	7'h20 :
		TR_19 = RG_rl_190 ;
	7'h21 :
		TR_19 = RG_rl_190 ;
	7'h22 :
		TR_19 = RG_rl_190 ;
	7'h23 :
		TR_19 = RG_rl_190 ;
	7'h24 :
		TR_19 = RG_rl_190 ;
	7'h25 :
		TR_19 = RG_rl_190 ;
	7'h26 :
		TR_19 = RG_rl_190 ;
	7'h27 :
		TR_19 = RG_rl_190 ;
	7'h28 :
		TR_19 = RG_rl_190 ;
	7'h29 :
		TR_19 = RG_rl_190 ;
	7'h2a :
		TR_19 = RG_rl_190 ;
	7'h2b :
		TR_19 = RG_rl_190 ;
	7'h2c :
		TR_19 = RG_rl_190 ;
	7'h2d :
		TR_19 = RG_rl_190 ;
	7'h2e :
		TR_19 = RG_rl_190 ;
	7'h2f :
		TR_19 = RG_rl_190 ;
	7'h30 :
		TR_19 = RG_rl_190 ;
	7'h31 :
		TR_19 = RG_rl_190 ;
	7'h32 :
		TR_19 = RG_rl_190 ;
	7'h33 :
		TR_19 = RG_rl_190 ;
	7'h34 :
		TR_19 = RG_rl_190 ;
	7'h35 :
		TR_19 = RG_rl_190 ;
	7'h36 :
		TR_19 = RG_rl_190 ;
	7'h37 :
		TR_19 = RG_rl_190 ;
	7'h38 :
		TR_19 = RG_rl_190 ;
	7'h39 :
		TR_19 = RG_rl_190 ;
	7'h3a :
		TR_19 = RG_rl_190 ;
	7'h3b :
		TR_19 = RG_rl_190 ;
	7'h3c :
		TR_19 = RG_rl_190 ;
	7'h3d :
		TR_19 = RG_rl_190 ;
	7'h3e :
		TR_19 = RG_rl_190 ;
	7'h3f :
		TR_19 = RG_rl_190 ;
	7'h40 :
		TR_19 = RG_rl_190 ;
	7'h41 :
		TR_19 = RG_rl_190 ;
	7'h42 :
		TR_19 = RG_rl_190 ;
	7'h43 :
		TR_19 = RG_rl_190 ;
	7'h44 :
		TR_19 = RG_rl_190 ;
	7'h45 :
		TR_19 = RG_rl_190 ;
	7'h46 :
		TR_19 = RG_rl_190 ;
	7'h47 :
		TR_19 = RG_rl_190 ;
	7'h48 :
		TR_19 = RG_rl_190 ;
	7'h49 :
		TR_19 = RG_rl_190 ;
	7'h4a :
		TR_19 = RG_rl_190 ;
	7'h4b :
		TR_19 = RG_rl_190 ;
	7'h4c :
		TR_19 = RG_rl_190 ;
	7'h4d :
		TR_19 = RG_rl_190 ;
	7'h4e :
		TR_19 = RG_rl_190 ;
	7'h4f :
		TR_19 = RG_rl_190 ;
	7'h50 :
		TR_19 = RG_rl_190 ;
	7'h51 :
		TR_19 = RG_rl_190 ;
	7'h52 :
		TR_19 = RG_rl_190 ;
	7'h53 :
		TR_19 = RG_rl_190 ;
	7'h54 :
		TR_19 = RG_rl_190 ;
	7'h55 :
		TR_19 = RG_rl_190 ;
	7'h56 :
		TR_19 = RG_rl_190 ;
	7'h57 :
		TR_19 = RG_rl_190 ;
	7'h58 :
		TR_19 = RG_rl_190 ;
	7'h59 :
		TR_19 = RG_rl_190 ;
	7'h5a :
		TR_19 = RG_rl_190 ;
	7'h5b :
		TR_19 = RG_rl_190 ;
	7'h5c :
		TR_19 = RG_rl_190 ;
	7'h5d :
		TR_19 = RG_rl_190 ;
	7'h5e :
		TR_19 = RG_rl_190 ;
	7'h5f :
		TR_19 = RG_rl_190 ;
	7'h60 :
		TR_19 = RG_rl_190 ;
	7'h61 :
		TR_19 = RG_rl_190 ;
	7'h62 :
		TR_19 = RG_rl_190 ;
	7'h63 :
		TR_19 = RG_rl_190 ;
	7'h64 :
		TR_19 = RG_rl_190 ;
	7'h65 :
		TR_19 = RG_rl_190 ;
	7'h66 :
		TR_19 = RG_rl_190 ;
	7'h67 :
		TR_19 = RG_rl_190 ;
	7'h68 :
		TR_19 = RG_rl_190 ;
	7'h69 :
		TR_19 = RG_rl_190 ;
	7'h6a :
		TR_19 = RG_rl_190 ;
	7'h6b :
		TR_19 = RG_rl_190 ;
	7'h6c :
		TR_19 = RG_rl_190 ;
	7'h6d :
		TR_19 = RG_rl_190 ;
	7'h6e :
		TR_19 = RG_rl_190 ;
	7'h6f :
		TR_19 = RG_rl_190 ;
	7'h70 :
		TR_19 = RG_rl_190 ;
	7'h71 :
		TR_19 = RG_rl_190 ;
	7'h72 :
		TR_19 = RG_rl_190 ;
	7'h73 :
		TR_19 = RG_rl_190 ;
	7'h74 :
		TR_19 = RG_rl_190 ;
	7'h75 :
		TR_19 = RG_rl_190 ;
	7'h76 :
		TR_19 = RG_rl_190 ;
	7'h77 :
		TR_19 = RG_rl_190 ;
	7'h78 :
		TR_19 = RG_rl_190 ;
	7'h79 :
		TR_19 = RG_rl_190 ;
	7'h7a :
		TR_19 = RG_rl_190 ;
	7'h7b :
		TR_19 = RG_rl_190 ;
	7'h7c :
		TR_19 = RG_rl_190 ;
	7'h7d :
		TR_19 = RG_rl_190 ;
	7'h7e :
		TR_19 = RG_rl_190 ;
	7'h7f :
		TR_19 = RG_rl_190 ;
	default :
		TR_19 = 9'hx ;
	endcase
always @ ( RG_rl_191 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_20 = RG_rl_191 ;
	7'h01 :
		TR_20 = RG_rl_191 ;
	7'h02 :
		TR_20 = RG_rl_191 ;
	7'h03 :
		TR_20 = RG_rl_191 ;
	7'h04 :
		TR_20 = RG_rl_191 ;
	7'h05 :
		TR_20 = RG_rl_191 ;
	7'h06 :
		TR_20 = RG_rl_191 ;
	7'h07 :
		TR_20 = RG_rl_191 ;
	7'h08 :
		TR_20 = 9'h000 ;	// line#=../rle.cpp:68
	7'h09 :
		TR_20 = RG_rl_191 ;
	7'h0a :
		TR_20 = RG_rl_191 ;
	7'h0b :
		TR_20 = RG_rl_191 ;
	7'h0c :
		TR_20 = RG_rl_191 ;
	7'h0d :
		TR_20 = RG_rl_191 ;
	7'h0e :
		TR_20 = RG_rl_191 ;
	7'h0f :
		TR_20 = RG_rl_191 ;
	7'h10 :
		TR_20 = RG_rl_191 ;
	7'h11 :
		TR_20 = RG_rl_191 ;
	7'h12 :
		TR_20 = RG_rl_191 ;
	7'h13 :
		TR_20 = RG_rl_191 ;
	7'h14 :
		TR_20 = RG_rl_191 ;
	7'h15 :
		TR_20 = RG_rl_191 ;
	7'h16 :
		TR_20 = RG_rl_191 ;
	7'h17 :
		TR_20 = RG_rl_191 ;
	7'h18 :
		TR_20 = RG_rl_191 ;
	7'h19 :
		TR_20 = RG_rl_191 ;
	7'h1a :
		TR_20 = RG_rl_191 ;
	7'h1b :
		TR_20 = RG_rl_191 ;
	7'h1c :
		TR_20 = RG_rl_191 ;
	7'h1d :
		TR_20 = RG_rl_191 ;
	7'h1e :
		TR_20 = RG_rl_191 ;
	7'h1f :
		TR_20 = RG_rl_191 ;
	7'h20 :
		TR_20 = RG_rl_191 ;
	7'h21 :
		TR_20 = RG_rl_191 ;
	7'h22 :
		TR_20 = RG_rl_191 ;
	7'h23 :
		TR_20 = RG_rl_191 ;
	7'h24 :
		TR_20 = RG_rl_191 ;
	7'h25 :
		TR_20 = RG_rl_191 ;
	7'h26 :
		TR_20 = RG_rl_191 ;
	7'h27 :
		TR_20 = RG_rl_191 ;
	7'h28 :
		TR_20 = RG_rl_191 ;
	7'h29 :
		TR_20 = RG_rl_191 ;
	7'h2a :
		TR_20 = RG_rl_191 ;
	7'h2b :
		TR_20 = RG_rl_191 ;
	7'h2c :
		TR_20 = RG_rl_191 ;
	7'h2d :
		TR_20 = RG_rl_191 ;
	7'h2e :
		TR_20 = RG_rl_191 ;
	7'h2f :
		TR_20 = RG_rl_191 ;
	7'h30 :
		TR_20 = RG_rl_191 ;
	7'h31 :
		TR_20 = RG_rl_191 ;
	7'h32 :
		TR_20 = RG_rl_191 ;
	7'h33 :
		TR_20 = RG_rl_191 ;
	7'h34 :
		TR_20 = RG_rl_191 ;
	7'h35 :
		TR_20 = RG_rl_191 ;
	7'h36 :
		TR_20 = RG_rl_191 ;
	7'h37 :
		TR_20 = RG_rl_191 ;
	7'h38 :
		TR_20 = RG_rl_191 ;
	7'h39 :
		TR_20 = RG_rl_191 ;
	7'h3a :
		TR_20 = RG_rl_191 ;
	7'h3b :
		TR_20 = RG_rl_191 ;
	7'h3c :
		TR_20 = RG_rl_191 ;
	7'h3d :
		TR_20 = RG_rl_191 ;
	7'h3e :
		TR_20 = RG_rl_191 ;
	7'h3f :
		TR_20 = RG_rl_191 ;
	7'h40 :
		TR_20 = RG_rl_191 ;
	7'h41 :
		TR_20 = RG_rl_191 ;
	7'h42 :
		TR_20 = RG_rl_191 ;
	7'h43 :
		TR_20 = RG_rl_191 ;
	7'h44 :
		TR_20 = RG_rl_191 ;
	7'h45 :
		TR_20 = RG_rl_191 ;
	7'h46 :
		TR_20 = RG_rl_191 ;
	7'h47 :
		TR_20 = RG_rl_191 ;
	7'h48 :
		TR_20 = RG_rl_191 ;
	7'h49 :
		TR_20 = RG_rl_191 ;
	7'h4a :
		TR_20 = RG_rl_191 ;
	7'h4b :
		TR_20 = RG_rl_191 ;
	7'h4c :
		TR_20 = RG_rl_191 ;
	7'h4d :
		TR_20 = RG_rl_191 ;
	7'h4e :
		TR_20 = RG_rl_191 ;
	7'h4f :
		TR_20 = RG_rl_191 ;
	7'h50 :
		TR_20 = RG_rl_191 ;
	7'h51 :
		TR_20 = RG_rl_191 ;
	7'h52 :
		TR_20 = RG_rl_191 ;
	7'h53 :
		TR_20 = RG_rl_191 ;
	7'h54 :
		TR_20 = RG_rl_191 ;
	7'h55 :
		TR_20 = RG_rl_191 ;
	7'h56 :
		TR_20 = RG_rl_191 ;
	7'h57 :
		TR_20 = RG_rl_191 ;
	7'h58 :
		TR_20 = RG_rl_191 ;
	7'h59 :
		TR_20 = RG_rl_191 ;
	7'h5a :
		TR_20 = RG_rl_191 ;
	7'h5b :
		TR_20 = RG_rl_191 ;
	7'h5c :
		TR_20 = RG_rl_191 ;
	7'h5d :
		TR_20 = RG_rl_191 ;
	7'h5e :
		TR_20 = RG_rl_191 ;
	7'h5f :
		TR_20 = RG_rl_191 ;
	7'h60 :
		TR_20 = RG_rl_191 ;
	7'h61 :
		TR_20 = RG_rl_191 ;
	7'h62 :
		TR_20 = RG_rl_191 ;
	7'h63 :
		TR_20 = RG_rl_191 ;
	7'h64 :
		TR_20 = RG_rl_191 ;
	7'h65 :
		TR_20 = RG_rl_191 ;
	7'h66 :
		TR_20 = RG_rl_191 ;
	7'h67 :
		TR_20 = RG_rl_191 ;
	7'h68 :
		TR_20 = RG_rl_191 ;
	7'h69 :
		TR_20 = RG_rl_191 ;
	7'h6a :
		TR_20 = RG_rl_191 ;
	7'h6b :
		TR_20 = RG_rl_191 ;
	7'h6c :
		TR_20 = RG_rl_191 ;
	7'h6d :
		TR_20 = RG_rl_191 ;
	7'h6e :
		TR_20 = RG_rl_191 ;
	7'h6f :
		TR_20 = RG_rl_191 ;
	7'h70 :
		TR_20 = RG_rl_191 ;
	7'h71 :
		TR_20 = RG_rl_191 ;
	7'h72 :
		TR_20 = RG_rl_191 ;
	7'h73 :
		TR_20 = RG_rl_191 ;
	7'h74 :
		TR_20 = RG_rl_191 ;
	7'h75 :
		TR_20 = RG_rl_191 ;
	7'h76 :
		TR_20 = RG_rl_191 ;
	7'h77 :
		TR_20 = RG_rl_191 ;
	7'h78 :
		TR_20 = RG_rl_191 ;
	7'h79 :
		TR_20 = RG_rl_191 ;
	7'h7a :
		TR_20 = RG_rl_191 ;
	7'h7b :
		TR_20 = RG_rl_191 ;
	7'h7c :
		TR_20 = RG_rl_191 ;
	7'h7d :
		TR_20 = RG_rl_191 ;
	7'h7e :
		TR_20 = RG_rl_191 ;
	7'h7f :
		TR_20 = RG_rl_191 ;
	default :
		TR_20 = 9'hx ;
	endcase
always @ ( RG_rl_192 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_21 = RG_rl_192 ;
	7'h01 :
		TR_21 = RG_rl_192 ;
	7'h02 :
		TR_21 = RG_rl_192 ;
	7'h03 :
		TR_21 = RG_rl_192 ;
	7'h04 :
		TR_21 = RG_rl_192 ;
	7'h05 :
		TR_21 = RG_rl_192 ;
	7'h06 :
		TR_21 = RG_rl_192 ;
	7'h07 :
		TR_21 = RG_rl_192 ;
	7'h08 :
		TR_21 = RG_rl_192 ;
	7'h09 :
		TR_21 = 9'h000 ;	// line#=../rle.cpp:68
	7'h0a :
		TR_21 = RG_rl_192 ;
	7'h0b :
		TR_21 = RG_rl_192 ;
	7'h0c :
		TR_21 = RG_rl_192 ;
	7'h0d :
		TR_21 = RG_rl_192 ;
	7'h0e :
		TR_21 = RG_rl_192 ;
	7'h0f :
		TR_21 = RG_rl_192 ;
	7'h10 :
		TR_21 = RG_rl_192 ;
	7'h11 :
		TR_21 = RG_rl_192 ;
	7'h12 :
		TR_21 = RG_rl_192 ;
	7'h13 :
		TR_21 = RG_rl_192 ;
	7'h14 :
		TR_21 = RG_rl_192 ;
	7'h15 :
		TR_21 = RG_rl_192 ;
	7'h16 :
		TR_21 = RG_rl_192 ;
	7'h17 :
		TR_21 = RG_rl_192 ;
	7'h18 :
		TR_21 = RG_rl_192 ;
	7'h19 :
		TR_21 = RG_rl_192 ;
	7'h1a :
		TR_21 = RG_rl_192 ;
	7'h1b :
		TR_21 = RG_rl_192 ;
	7'h1c :
		TR_21 = RG_rl_192 ;
	7'h1d :
		TR_21 = RG_rl_192 ;
	7'h1e :
		TR_21 = RG_rl_192 ;
	7'h1f :
		TR_21 = RG_rl_192 ;
	7'h20 :
		TR_21 = RG_rl_192 ;
	7'h21 :
		TR_21 = RG_rl_192 ;
	7'h22 :
		TR_21 = RG_rl_192 ;
	7'h23 :
		TR_21 = RG_rl_192 ;
	7'h24 :
		TR_21 = RG_rl_192 ;
	7'h25 :
		TR_21 = RG_rl_192 ;
	7'h26 :
		TR_21 = RG_rl_192 ;
	7'h27 :
		TR_21 = RG_rl_192 ;
	7'h28 :
		TR_21 = RG_rl_192 ;
	7'h29 :
		TR_21 = RG_rl_192 ;
	7'h2a :
		TR_21 = RG_rl_192 ;
	7'h2b :
		TR_21 = RG_rl_192 ;
	7'h2c :
		TR_21 = RG_rl_192 ;
	7'h2d :
		TR_21 = RG_rl_192 ;
	7'h2e :
		TR_21 = RG_rl_192 ;
	7'h2f :
		TR_21 = RG_rl_192 ;
	7'h30 :
		TR_21 = RG_rl_192 ;
	7'h31 :
		TR_21 = RG_rl_192 ;
	7'h32 :
		TR_21 = RG_rl_192 ;
	7'h33 :
		TR_21 = RG_rl_192 ;
	7'h34 :
		TR_21 = RG_rl_192 ;
	7'h35 :
		TR_21 = RG_rl_192 ;
	7'h36 :
		TR_21 = RG_rl_192 ;
	7'h37 :
		TR_21 = RG_rl_192 ;
	7'h38 :
		TR_21 = RG_rl_192 ;
	7'h39 :
		TR_21 = RG_rl_192 ;
	7'h3a :
		TR_21 = RG_rl_192 ;
	7'h3b :
		TR_21 = RG_rl_192 ;
	7'h3c :
		TR_21 = RG_rl_192 ;
	7'h3d :
		TR_21 = RG_rl_192 ;
	7'h3e :
		TR_21 = RG_rl_192 ;
	7'h3f :
		TR_21 = RG_rl_192 ;
	7'h40 :
		TR_21 = RG_rl_192 ;
	7'h41 :
		TR_21 = RG_rl_192 ;
	7'h42 :
		TR_21 = RG_rl_192 ;
	7'h43 :
		TR_21 = RG_rl_192 ;
	7'h44 :
		TR_21 = RG_rl_192 ;
	7'h45 :
		TR_21 = RG_rl_192 ;
	7'h46 :
		TR_21 = RG_rl_192 ;
	7'h47 :
		TR_21 = RG_rl_192 ;
	7'h48 :
		TR_21 = RG_rl_192 ;
	7'h49 :
		TR_21 = RG_rl_192 ;
	7'h4a :
		TR_21 = RG_rl_192 ;
	7'h4b :
		TR_21 = RG_rl_192 ;
	7'h4c :
		TR_21 = RG_rl_192 ;
	7'h4d :
		TR_21 = RG_rl_192 ;
	7'h4e :
		TR_21 = RG_rl_192 ;
	7'h4f :
		TR_21 = RG_rl_192 ;
	7'h50 :
		TR_21 = RG_rl_192 ;
	7'h51 :
		TR_21 = RG_rl_192 ;
	7'h52 :
		TR_21 = RG_rl_192 ;
	7'h53 :
		TR_21 = RG_rl_192 ;
	7'h54 :
		TR_21 = RG_rl_192 ;
	7'h55 :
		TR_21 = RG_rl_192 ;
	7'h56 :
		TR_21 = RG_rl_192 ;
	7'h57 :
		TR_21 = RG_rl_192 ;
	7'h58 :
		TR_21 = RG_rl_192 ;
	7'h59 :
		TR_21 = RG_rl_192 ;
	7'h5a :
		TR_21 = RG_rl_192 ;
	7'h5b :
		TR_21 = RG_rl_192 ;
	7'h5c :
		TR_21 = RG_rl_192 ;
	7'h5d :
		TR_21 = RG_rl_192 ;
	7'h5e :
		TR_21 = RG_rl_192 ;
	7'h5f :
		TR_21 = RG_rl_192 ;
	7'h60 :
		TR_21 = RG_rl_192 ;
	7'h61 :
		TR_21 = RG_rl_192 ;
	7'h62 :
		TR_21 = RG_rl_192 ;
	7'h63 :
		TR_21 = RG_rl_192 ;
	7'h64 :
		TR_21 = RG_rl_192 ;
	7'h65 :
		TR_21 = RG_rl_192 ;
	7'h66 :
		TR_21 = RG_rl_192 ;
	7'h67 :
		TR_21 = RG_rl_192 ;
	7'h68 :
		TR_21 = RG_rl_192 ;
	7'h69 :
		TR_21 = RG_rl_192 ;
	7'h6a :
		TR_21 = RG_rl_192 ;
	7'h6b :
		TR_21 = RG_rl_192 ;
	7'h6c :
		TR_21 = RG_rl_192 ;
	7'h6d :
		TR_21 = RG_rl_192 ;
	7'h6e :
		TR_21 = RG_rl_192 ;
	7'h6f :
		TR_21 = RG_rl_192 ;
	7'h70 :
		TR_21 = RG_rl_192 ;
	7'h71 :
		TR_21 = RG_rl_192 ;
	7'h72 :
		TR_21 = RG_rl_192 ;
	7'h73 :
		TR_21 = RG_rl_192 ;
	7'h74 :
		TR_21 = RG_rl_192 ;
	7'h75 :
		TR_21 = RG_rl_192 ;
	7'h76 :
		TR_21 = RG_rl_192 ;
	7'h77 :
		TR_21 = RG_rl_192 ;
	7'h78 :
		TR_21 = RG_rl_192 ;
	7'h79 :
		TR_21 = RG_rl_192 ;
	7'h7a :
		TR_21 = RG_rl_192 ;
	7'h7b :
		TR_21 = RG_rl_192 ;
	7'h7c :
		TR_21 = RG_rl_192 ;
	7'h7d :
		TR_21 = RG_rl_192 ;
	7'h7e :
		TR_21 = RG_rl_192 ;
	7'h7f :
		TR_21 = RG_rl_192 ;
	default :
		TR_21 = 9'hx ;
	endcase
always @ ( RG_rl_193 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_22 = RG_rl_193 ;
	7'h01 :
		TR_22 = RG_rl_193 ;
	7'h02 :
		TR_22 = RG_rl_193 ;
	7'h03 :
		TR_22 = RG_rl_193 ;
	7'h04 :
		TR_22 = RG_rl_193 ;
	7'h05 :
		TR_22 = RG_rl_193 ;
	7'h06 :
		TR_22 = RG_rl_193 ;
	7'h07 :
		TR_22 = RG_rl_193 ;
	7'h08 :
		TR_22 = RG_rl_193 ;
	7'h09 :
		TR_22 = RG_rl_193 ;
	7'h0a :
		TR_22 = 9'h000 ;	// line#=../rle.cpp:68
	7'h0b :
		TR_22 = RG_rl_193 ;
	7'h0c :
		TR_22 = RG_rl_193 ;
	7'h0d :
		TR_22 = RG_rl_193 ;
	7'h0e :
		TR_22 = RG_rl_193 ;
	7'h0f :
		TR_22 = RG_rl_193 ;
	7'h10 :
		TR_22 = RG_rl_193 ;
	7'h11 :
		TR_22 = RG_rl_193 ;
	7'h12 :
		TR_22 = RG_rl_193 ;
	7'h13 :
		TR_22 = RG_rl_193 ;
	7'h14 :
		TR_22 = RG_rl_193 ;
	7'h15 :
		TR_22 = RG_rl_193 ;
	7'h16 :
		TR_22 = RG_rl_193 ;
	7'h17 :
		TR_22 = RG_rl_193 ;
	7'h18 :
		TR_22 = RG_rl_193 ;
	7'h19 :
		TR_22 = RG_rl_193 ;
	7'h1a :
		TR_22 = RG_rl_193 ;
	7'h1b :
		TR_22 = RG_rl_193 ;
	7'h1c :
		TR_22 = RG_rl_193 ;
	7'h1d :
		TR_22 = RG_rl_193 ;
	7'h1e :
		TR_22 = RG_rl_193 ;
	7'h1f :
		TR_22 = RG_rl_193 ;
	7'h20 :
		TR_22 = RG_rl_193 ;
	7'h21 :
		TR_22 = RG_rl_193 ;
	7'h22 :
		TR_22 = RG_rl_193 ;
	7'h23 :
		TR_22 = RG_rl_193 ;
	7'h24 :
		TR_22 = RG_rl_193 ;
	7'h25 :
		TR_22 = RG_rl_193 ;
	7'h26 :
		TR_22 = RG_rl_193 ;
	7'h27 :
		TR_22 = RG_rl_193 ;
	7'h28 :
		TR_22 = RG_rl_193 ;
	7'h29 :
		TR_22 = RG_rl_193 ;
	7'h2a :
		TR_22 = RG_rl_193 ;
	7'h2b :
		TR_22 = RG_rl_193 ;
	7'h2c :
		TR_22 = RG_rl_193 ;
	7'h2d :
		TR_22 = RG_rl_193 ;
	7'h2e :
		TR_22 = RG_rl_193 ;
	7'h2f :
		TR_22 = RG_rl_193 ;
	7'h30 :
		TR_22 = RG_rl_193 ;
	7'h31 :
		TR_22 = RG_rl_193 ;
	7'h32 :
		TR_22 = RG_rl_193 ;
	7'h33 :
		TR_22 = RG_rl_193 ;
	7'h34 :
		TR_22 = RG_rl_193 ;
	7'h35 :
		TR_22 = RG_rl_193 ;
	7'h36 :
		TR_22 = RG_rl_193 ;
	7'h37 :
		TR_22 = RG_rl_193 ;
	7'h38 :
		TR_22 = RG_rl_193 ;
	7'h39 :
		TR_22 = RG_rl_193 ;
	7'h3a :
		TR_22 = RG_rl_193 ;
	7'h3b :
		TR_22 = RG_rl_193 ;
	7'h3c :
		TR_22 = RG_rl_193 ;
	7'h3d :
		TR_22 = RG_rl_193 ;
	7'h3e :
		TR_22 = RG_rl_193 ;
	7'h3f :
		TR_22 = RG_rl_193 ;
	7'h40 :
		TR_22 = RG_rl_193 ;
	7'h41 :
		TR_22 = RG_rl_193 ;
	7'h42 :
		TR_22 = RG_rl_193 ;
	7'h43 :
		TR_22 = RG_rl_193 ;
	7'h44 :
		TR_22 = RG_rl_193 ;
	7'h45 :
		TR_22 = RG_rl_193 ;
	7'h46 :
		TR_22 = RG_rl_193 ;
	7'h47 :
		TR_22 = RG_rl_193 ;
	7'h48 :
		TR_22 = RG_rl_193 ;
	7'h49 :
		TR_22 = RG_rl_193 ;
	7'h4a :
		TR_22 = RG_rl_193 ;
	7'h4b :
		TR_22 = RG_rl_193 ;
	7'h4c :
		TR_22 = RG_rl_193 ;
	7'h4d :
		TR_22 = RG_rl_193 ;
	7'h4e :
		TR_22 = RG_rl_193 ;
	7'h4f :
		TR_22 = RG_rl_193 ;
	7'h50 :
		TR_22 = RG_rl_193 ;
	7'h51 :
		TR_22 = RG_rl_193 ;
	7'h52 :
		TR_22 = RG_rl_193 ;
	7'h53 :
		TR_22 = RG_rl_193 ;
	7'h54 :
		TR_22 = RG_rl_193 ;
	7'h55 :
		TR_22 = RG_rl_193 ;
	7'h56 :
		TR_22 = RG_rl_193 ;
	7'h57 :
		TR_22 = RG_rl_193 ;
	7'h58 :
		TR_22 = RG_rl_193 ;
	7'h59 :
		TR_22 = RG_rl_193 ;
	7'h5a :
		TR_22 = RG_rl_193 ;
	7'h5b :
		TR_22 = RG_rl_193 ;
	7'h5c :
		TR_22 = RG_rl_193 ;
	7'h5d :
		TR_22 = RG_rl_193 ;
	7'h5e :
		TR_22 = RG_rl_193 ;
	7'h5f :
		TR_22 = RG_rl_193 ;
	7'h60 :
		TR_22 = RG_rl_193 ;
	7'h61 :
		TR_22 = RG_rl_193 ;
	7'h62 :
		TR_22 = RG_rl_193 ;
	7'h63 :
		TR_22 = RG_rl_193 ;
	7'h64 :
		TR_22 = RG_rl_193 ;
	7'h65 :
		TR_22 = RG_rl_193 ;
	7'h66 :
		TR_22 = RG_rl_193 ;
	7'h67 :
		TR_22 = RG_rl_193 ;
	7'h68 :
		TR_22 = RG_rl_193 ;
	7'h69 :
		TR_22 = RG_rl_193 ;
	7'h6a :
		TR_22 = RG_rl_193 ;
	7'h6b :
		TR_22 = RG_rl_193 ;
	7'h6c :
		TR_22 = RG_rl_193 ;
	7'h6d :
		TR_22 = RG_rl_193 ;
	7'h6e :
		TR_22 = RG_rl_193 ;
	7'h6f :
		TR_22 = RG_rl_193 ;
	7'h70 :
		TR_22 = RG_rl_193 ;
	7'h71 :
		TR_22 = RG_rl_193 ;
	7'h72 :
		TR_22 = RG_rl_193 ;
	7'h73 :
		TR_22 = RG_rl_193 ;
	7'h74 :
		TR_22 = RG_rl_193 ;
	7'h75 :
		TR_22 = RG_rl_193 ;
	7'h76 :
		TR_22 = RG_rl_193 ;
	7'h77 :
		TR_22 = RG_rl_193 ;
	7'h78 :
		TR_22 = RG_rl_193 ;
	7'h79 :
		TR_22 = RG_rl_193 ;
	7'h7a :
		TR_22 = RG_rl_193 ;
	7'h7b :
		TR_22 = RG_rl_193 ;
	7'h7c :
		TR_22 = RG_rl_193 ;
	7'h7d :
		TR_22 = RG_rl_193 ;
	7'h7e :
		TR_22 = RG_rl_193 ;
	7'h7f :
		TR_22 = RG_rl_193 ;
	default :
		TR_22 = 9'hx ;
	endcase
always @ ( RG_rl_194 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_23 = RG_rl_194 ;
	7'h01 :
		TR_23 = RG_rl_194 ;
	7'h02 :
		TR_23 = RG_rl_194 ;
	7'h03 :
		TR_23 = RG_rl_194 ;
	7'h04 :
		TR_23 = RG_rl_194 ;
	7'h05 :
		TR_23 = RG_rl_194 ;
	7'h06 :
		TR_23 = RG_rl_194 ;
	7'h07 :
		TR_23 = RG_rl_194 ;
	7'h08 :
		TR_23 = RG_rl_194 ;
	7'h09 :
		TR_23 = RG_rl_194 ;
	7'h0a :
		TR_23 = RG_rl_194 ;
	7'h0b :
		TR_23 = 9'h000 ;	// line#=../rle.cpp:68
	7'h0c :
		TR_23 = RG_rl_194 ;
	7'h0d :
		TR_23 = RG_rl_194 ;
	7'h0e :
		TR_23 = RG_rl_194 ;
	7'h0f :
		TR_23 = RG_rl_194 ;
	7'h10 :
		TR_23 = RG_rl_194 ;
	7'h11 :
		TR_23 = RG_rl_194 ;
	7'h12 :
		TR_23 = RG_rl_194 ;
	7'h13 :
		TR_23 = RG_rl_194 ;
	7'h14 :
		TR_23 = RG_rl_194 ;
	7'h15 :
		TR_23 = RG_rl_194 ;
	7'h16 :
		TR_23 = RG_rl_194 ;
	7'h17 :
		TR_23 = RG_rl_194 ;
	7'h18 :
		TR_23 = RG_rl_194 ;
	7'h19 :
		TR_23 = RG_rl_194 ;
	7'h1a :
		TR_23 = RG_rl_194 ;
	7'h1b :
		TR_23 = RG_rl_194 ;
	7'h1c :
		TR_23 = RG_rl_194 ;
	7'h1d :
		TR_23 = RG_rl_194 ;
	7'h1e :
		TR_23 = RG_rl_194 ;
	7'h1f :
		TR_23 = RG_rl_194 ;
	7'h20 :
		TR_23 = RG_rl_194 ;
	7'h21 :
		TR_23 = RG_rl_194 ;
	7'h22 :
		TR_23 = RG_rl_194 ;
	7'h23 :
		TR_23 = RG_rl_194 ;
	7'h24 :
		TR_23 = RG_rl_194 ;
	7'h25 :
		TR_23 = RG_rl_194 ;
	7'h26 :
		TR_23 = RG_rl_194 ;
	7'h27 :
		TR_23 = RG_rl_194 ;
	7'h28 :
		TR_23 = RG_rl_194 ;
	7'h29 :
		TR_23 = RG_rl_194 ;
	7'h2a :
		TR_23 = RG_rl_194 ;
	7'h2b :
		TR_23 = RG_rl_194 ;
	7'h2c :
		TR_23 = RG_rl_194 ;
	7'h2d :
		TR_23 = RG_rl_194 ;
	7'h2e :
		TR_23 = RG_rl_194 ;
	7'h2f :
		TR_23 = RG_rl_194 ;
	7'h30 :
		TR_23 = RG_rl_194 ;
	7'h31 :
		TR_23 = RG_rl_194 ;
	7'h32 :
		TR_23 = RG_rl_194 ;
	7'h33 :
		TR_23 = RG_rl_194 ;
	7'h34 :
		TR_23 = RG_rl_194 ;
	7'h35 :
		TR_23 = RG_rl_194 ;
	7'h36 :
		TR_23 = RG_rl_194 ;
	7'h37 :
		TR_23 = RG_rl_194 ;
	7'h38 :
		TR_23 = RG_rl_194 ;
	7'h39 :
		TR_23 = RG_rl_194 ;
	7'h3a :
		TR_23 = RG_rl_194 ;
	7'h3b :
		TR_23 = RG_rl_194 ;
	7'h3c :
		TR_23 = RG_rl_194 ;
	7'h3d :
		TR_23 = RG_rl_194 ;
	7'h3e :
		TR_23 = RG_rl_194 ;
	7'h3f :
		TR_23 = RG_rl_194 ;
	7'h40 :
		TR_23 = RG_rl_194 ;
	7'h41 :
		TR_23 = RG_rl_194 ;
	7'h42 :
		TR_23 = RG_rl_194 ;
	7'h43 :
		TR_23 = RG_rl_194 ;
	7'h44 :
		TR_23 = RG_rl_194 ;
	7'h45 :
		TR_23 = RG_rl_194 ;
	7'h46 :
		TR_23 = RG_rl_194 ;
	7'h47 :
		TR_23 = RG_rl_194 ;
	7'h48 :
		TR_23 = RG_rl_194 ;
	7'h49 :
		TR_23 = RG_rl_194 ;
	7'h4a :
		TR_23 = RG_rl_194 ;
	7'h4b :
		TR_23 = RG_rl_194 ;
	7'h4c :
		TR_23 = RG_rl_194 ;
	7'h4d :
		TR_23 = RG_rl_194 ;
	7'h4e :
		TR_23 = RG_rl_194 ;
	7'h4f :
		TR_23 = RG_rl_194 ;
	7'h50 :
		TR_23 = RG_rl_194 ;
	7'h51 :
		TR_23 = RG_rl_194 ;
	7'h52 :
		TR_23 = RG_rl_194 ;
	7'h53 :
		TR_23 = RG_rl_194 ;
	7'h54 :
		TR_23 = RG_rl_194 ;
	7'h55 :
		TR_23 = RG_rl_194 ;
	7'h56 :
		TR_23 = RG_rl_194 ;
	7'h57 :
		TR_23 = RG_rl_194 ;
	7'h58 :
		TR_23 = RG_rl_194 ;
	7'h59 :
		TR_23 = RG_rl_194 ;
	7'h5a :
		TR_23 = RG_rl_194 ;
	7'h5b :
		TR_23 = RG_rl_194 ;
	7'h5c :
		TR_23 = RG_rl_194 ;
	7'h5d :
		TR_23 = RG_rl_194 ;
	7'h5e :
		TR_23 = RG_rl_194 ;
	7'h5f :
		TR_23 = RG_rl_194 ;
	7'h60 :
		TR_23 = RG_rl_194 ;
	7'h61 :
		TR_23 = RG_rl_194 ;
	7'h62 :
		TR_23 = RG_rl_194 ;
	7'h63 :
		TR_23 = RG_rl_194 ;
	7'h64 :
		TR_23 = RG_rl_194 ;
	7'h65 :
		TR_23 = RG_rl_194 ;
	7'h66 :
		TR_23 = RG_rl_194 ;
	7'h67 :
		TR_23 = RG_rl_194 ;
	7'h68 :
		TR_23 = RG_rl_194 ;
	7'h69 :
		TR_23 = RG_rl_194 ;
	7'h6a :
		TR_23 = RG_rl_194 ;
	7'h6b :
		TR_23 = RG_rl_194 ;
	7'h6c :
		TR_23 = RG_rl_194 ;
	7'h6d :
		TR_23 = RG_rl_194 ;
	7'h6e :
		TR_23 = RG_rl_194 ;
	7'h6f :
		TR_23 = RG_rl_194 ;
	7'h70 :
		TR_23 = RG_rl_194 ;
	7'h71 :
		TR_23 = RG_rl_194 ;
	7'h72 :
		TR_23 = RG_rl_194 ;
	7'h73 :
		TR_23 = RG_rl_194 ;
	7'h74 :
		TR_23 = RG_rl_194 ;
	7'h75 :
		TR_23 = RG_rl_194 ;
	7'h76 :
		TR_23 = RG_rl_194 ;
	7'h77 :
		TR_23 = RG_rl_194 ;
	7'h78 :
		TR_23 = RG_rl_194 ;
	7'h79 :
		TR_23 = RG_rl_194 ;
	7'h7a :
		TR_23 = RG_rl_194 ;
	7'h7b :
		TR_23 = RG_rl_194 ;
	7'h7c :
		TR_23 = RG_rl_194 ;
	7'h7d :
		TR_23 = RG_rl_194 ;
	7'h7e :
		TR_23 = RG_rl_194 ;
	7'h7f :
		TR_23 = RG_rl_194 ;
	default :
		TR_23 = 9'hx ;
	endcase
always @ ( RG_rl_195 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_24 = RG_rl_195 ;
	7'h01 :
		TR_24 = RG_rl_195 ;
	7'h02 :
		TR_24 = RG_rl_195 ;
	7'h03 :
		TR_24 = RG_rl_195 ;
	7'h04 :
		TR_24 = RG_rl_195 ;
	7'h05 :
		TR_24 = RG_rl_195 ;
	7'h06 :
		TR_24 = RG_rl_195 ;
	7'h07 :
		TR_24 = RG_rl_195 ;
	7'h08 :
		TR_24 = RG_rl_195 ;
	7'h09 :
		TR_24 = RG_rl_195 ;
	7'h0a :
		TR_24 = RG_rl_195 ;
	7'h0b :
		TR_24 = RG_rl_195 ;
	7'h0c :
		TR_24 = 9'h000 ;	// line#=../rle.cpp:68
	7'h0d :
		TR_24 = RG_rl_195 ;
	7'h0e :
		TR_24 = RG_rl_195 ;
	7'h0f :
		TR_24 = RG_rl_195 ;
	7'h10 :
		TR_24 = RG_rl_195 ;
	7'h11 :
		TR_24 = RG_rl_195 ;
	7'h12 :
		TR_24 = RG_rl_195 ;
	7'h13 :
		TR_24 = RG_rl_195 ;
	7'h14 :
		TR_24 = RG_rl_195 ;
	7'h15 :
		TR_24 = RG_rl_195 ;
	7'h16 :
		TR_24 = RG_rl_195 ;
	7'h17 :
		TR_24 = RG_rl_195 ;
	7'h18 :
		TR_24 = RG_rl_195 ;
	7'h19 :
		TR_24 = RG_rl_195 ;
	7'h1a :
		TR_24 = RG_rl_195 ;
	7'h1b :
		TR_24 = RG_rl_195 ;
	7'h1c :
		TR_24 = RG_rl_195 ;
	7'h1d :
		TR_24 = RG_rl_195 ;
	7'h1e :
		TR_24 = RG_rl_195 ;
	7'h1f :
		TR_24 = RG_rl_195 ;
	7'h20 :
		TR_24 = RG_rl_195 ;
	7'h21 :
		TR_24 = RG_rl_195 ;
	7'h22 :
		TR_24 = RG_rl_195 ;
	7'h23 :
		TR_24 = RG_rl_195 ;
	7'h24 :
		TR_24 = RG_rl_195 ;
	7'h25 :
		TR_24 = RG_rl_195 ;
	7'h26 :
		TR_24 = RG_rl_195 ;
	7'h27 :
		TR_24 = RG_rl_195 ;
	7'h28 :
		TR_24 = RG_rl_195 ;
	7'h29 :
		TR_24 = RG_rl_195 ;
	7'h2a :
		TR_24 = RG_rl_195 ;
	7'h2b :
		TR_24 = RG_rl_195 ;
	7'h2c :
		TR_24 = RG_rl_195 ;
	7'h2d :
		TR_24 = RG_rl_195 ;
	7'h2e :
		TR_24 = RG_rl_195 ;
	7'h2f :
		TR_24 = RG_rl_195 ;
	7'h30 :
		TR_24 = RG_rl_195 ;
	7'h31 :
		TR_24 = RG_rl_195 ;
	7'h32 :
		TR_24 = RG_rl_195 ;
	7'h33 :
		TR_24 = RG_rl_195 ;
	7'h34 :
		TR_24 = RG_rl_195 ;
	7'h35 :
		TR_24 = RG_rl_195 ;
	7'h36 :
		TR_24 = RG_rl_195 ;
	7'h37 :
		TR_24 = RG_rl_195 ;
	7'h38 :
		TR_24 = RG_rl_195 ;
	7'h39 :
		TR_24 = RG_rl_195 ;
	7'h3a :
		TR_24 = RG_rl_195 ;
	7'h3b :
		TR_24 = RG_rl_195 ;
	7'h3c :
		TR_24 = RG_rl_195 ;
	7'h3d :
		TR_24 = RG_rl_195 ;
	7'h3e :
		TR_24 = RG_rl_195 ;
	7'h3f :
		TR_24 = RG_rl_195 ;
	7'h40 :
		TR_24 = RG_rl_195 ;
	7'h41 :
		TR_24 = RG_rl_195 ;
	7'h42 :
		TR_24 = RG_rl_195 ;
	7'h43 :
		TR_24 = RG_rl_195 ;
	7'h44 :
		TR_24 = RG_rl_195 ;
	7'h45 :
		TR_24 = RG_rl_195 ;
	7'h46 :
		TR_24 = RG_rl_195 ;
	7'h47 :
		TR_24 = RG_rl_195 ;
	7'h48 :
		TR_24 = RG_rl_195 ;
	7'h49 :
		TR_24 = RG_rl_195 ;
	7'h4a :
		TR_24 = RG_rl_195 ;
	7'h4b :
		TR_24 = RG_rl_195 ;
	7'h4c :
		TR_24 = RG_rl_195 ;
	7'h4d :
		TR_24 = RG_rl_195 ;
	7'h4e :
		TR_24 = RG_rl_195 ;
	7'h4f :
		TR_24 = RG_rl_195 ;
	7'h50 :
		TR_24 = RG_rl_195 ;
	7'h51 :
		TR_24 = RG_rl_195 ;
	7'h52 :
		TR_24 = RG_rl_195 ;
	7'h53 :
		TR_24 = RG_rl_195 ;
	7'h54 :
		TR_24 = RG_rl_195 ;
	7'h55 :
		TR_24 = RG_rl_195 ;
	7'h56 :
		TR_24 = RG_rl_195 ;
	7'h57 :
		TR_24 = RG_rl_195 ;
	7'h58 :
		TR_24 = RG_rl_195 ;
	7'h59 :
		TR_24 = RG_rl_195 ;
	7'h5a :
		TR_24 = RG_rl_195 ;
	7'h5b :
		TR_24 = RG_rl_195 ;
	7'h5c :
		TR_24 = RG_rl_195 ;
	7'h5d :
		TR_24 = RG_rl_195 ;
	7'h5e :
		TR_24 = RG_rl_195 ;
	7'h5f :
		TR_24 = RG_rl_195 ;
	7'h60 :
		TR_24 = RG_rl_195 ;
	7'h61 :
		TR_24 = RG_rl_195 ;
	7'h62 :
		TR_24 = RG_rl_195 ;
	7'h63 :
		TR_24 = RG_rl_195 ;
	7'h64 :
		TR_24 = RG_rl_195 ;
	7'h65 :
		TR_24 = RG_rl_195 ;
	7'h66 :
		TR_24 = RG_rl_195 ;
	7'h67 :
		TR_24 = RG_rl_195 ;
	7'h68 :
		TR_24 = RG_rl_195 ;
	7'h69 :
		TR_24 = RG_rl_195 ;
	7'h6a :
		TR_24 = RG_rl_195 ;
	7'h6b :
		TR_24 = RG_rl_195 ;
	7'h6c :
		TR_24 = RG_rl_195 ;
	7'h6d :
		TR_24 = RG_rl_195 ;
	7'h6e :
		TR_24 = RG_rl_195 ;
	7'h6f :
		TR_24 = RG_rl_195 ;
	7'h70 :
		TR_24 = RG_rl_195 ;
	7'h71 :
		TR_24 = RG_rl_195 ;
	7'h72 :
		TR_24 = RG_rl_195 ;
	7'h73 :
		TR_24 = RG_rl_195 ;
	7'h74 :
		TR_24 = RG_rl_195 ;
	7'h75 :
		TR_24 = RG_rl_195 ;
	7'h76 :
		TR_24 = RG_rl_195 ;
	7'h77 :
		TR_24 = RG_rl_195 ;
	7'h78 :
		TR_24 = RG_rl_195 ;
	7'h79 :
		TR_24 = RG_rl_195 ;
	7'h7a :
		TR_24 = RG_rl_195 ;
	7'h7b :
		TR_24 = RG_rl_195 ;
	7'h7c :
		TR_24 = RG_rl_195 ;
	7'h7d :
		TR_24 = RG_rl_195 ;
	7'h7e :
		TR_24 = RG_rl_195 ;
	7'h7f :
		TR_24 = RG_rl_195 ;
	default :
		TR_24 = 9'hx ;
	endcase
always @ ( RG_rl_196 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_25 = RG_rl_196 ;
	7'h01 :
		TR_25 = RG_rl_196 ;
	7'h02 :
		TR_25 = RG_rl_196 ;
	7'h03 :
		TR_25 = RG_rl_196 ;
	7'h04 :
		TR_25 = RG_rl_196 ;
	7'h05 :
		TR_25 = RG_rl_196 ;
	7'h06 :
		TR_25 = RG_rl_196 ;
	7'h07 :
		TR_25 = RG_rl_196 ;
	7'h08 :
		TR_25 = RG_rl_196 ;
	7'h09 :
		TR_25 = RG_rl_196 ;
	7'h0a :
		TR_25 = RG_rl_196 ;
	7'h0b :
		TR_25 = RG_rl_196 ;
	7'h0c :
		TR_25 = RG_rl_196 ;
	7'h0d :
		TR_25 = 9'h000 ;	// line#=../rle.cpp:68
	7'h0e :
		TR_25 = RG_rl_196 ;
	7'h0f :
		TR_25 = RG_rl_196 ;
	7'h10 :
		TR_25 = RG_rl_196 ;
	7'h11 :
		TR_25 = RG_rl_196 ;
	7'h12 :
		TR_25 = RG_rl_196 ;
	7'h13 :
		TR_25 = RG_rl_196 ;
	7'h14 :
		TR_25 = RG_rl_196 ;
	7'h15 :
		TR_25 = RG_rl_196 ;
	7'h16 :
		TR_25 = RG_rl_196 ;
	7'h17 :
		TR_25 = RG_rl_196 ;
	7'h18 :
		TR_25 = RG_rl_196 ;
	7'h19 :
		TR_25 = RG_rl_196 ;
	7'h1a :
		TR_25 = RG_rl_196 ;
	7'h1b :
		TR_25 = RG_rl_196 ;
	7'h1c :
		TR_25 = RG_rl_196 ;
	7'h1d :
		TR_25 = RG_rl_196 ;
	7'h1e :
		TR_25 = RG_rl_196 ;
	7'h1f :
		TR_25 = RG_rl_196 ;
	7'h20 :
		TR_25 = RG_rl_196 ;
	7'h21 :
		TR_25 = RG_rl_196 ;
	7'h22 :
		TR_25 = RG_rl_196 ;
	7'h23 :
		TR_25 = RG_rl_196 ;
	7'h24 :
		TR_25 = RG_rl_196 ;
	7'h25 :
		TR_25 = RG_rl_196 ;
	7'h26 :
		TR_25 = RG_rl_196 ;
	7'h27 :
		TR_25 = RG_rl_196 ;
	7'h28 :
		TR_25 = RG_rl_196 ;
	7'h29 :
		TR_25 = RG_rl_196 ;
	7'h2a :
		TR_25 = RG_rl_196 ;
	7'h2b :
		TR_25 = RG_rl_196 ;
	7'h2c :
		TR_25 = RG_rl_196 ;
	7'h2d :
		TR_25 = RG_rl_196 ;
	7'h2e :
		TR_25 = RG_rl_196 ;
	7'h2f :
		TR_25 = RG_rl_196 ;
	7'h30 :
		TR_25 = RG_rl_196 ;
	7'h31 :
		TR_25 = RG_rl_196 ;
	7'h32 :
		TR_25 = RG_rl_196 ;
	7'h33 :
		TR_25 = RG_rl_196 ;
	7'h34 :
		TR_25 = RG_rl_196 ;
	7'h35 :
		TR_25 = RG_rl_196 ;
	7'h36 :
		TR_25 = RG_rl_196 ;
	7'h37 :
		TR_25 = RG_rl_196 ;
	7'h38 :
		TR_25 = RG_rl_196 ;
	7'h39 :
		TR_25 = RG_rl_196 ;
	7'h3a :
		TR_25 = RG_rl_196 ;
	7'h3b :
		TR_25 = RG_rl_196 ;
	7'h3c :
		TR_25 = RG_rl_196 ;
	7'h3d :
		TR_25 = RG_rl_196 ;
	7'h3e :
		TR_25 = RG_rl_196 ;
	7'h3f :
		TR_25 = RG_rl_196 ;
	7'h40 :
		TR_25 = RG_rl_196 ;
	7'h41 :
		TR_25 = RG_rl_196 ;
	7'h42 :
		TR_25 = RG_rl_196 ;
	7'h43 :
		TR_25 = RG_rl_196 ;
	7'h44 :
		TR_25 = RG_rl_196 ;
	7'h45 :
		TR_25 = RG_rl_196 ;
	7'h46 :
		TR_25 = RG_rl_196 ;
	7'h47 :
		TR_25 = RG_rl_196 ;
	7'h48 :
		TR_25 = RG_rl_196 ;
	7'h49 :
		TR_25 = RG_rl_196 ;
	7'h4a :
		TR_25 = RG_rl_196 ;
	7'h4b :
		TR_25 = RG_rl_196 ;
	7'h4c :
		TR_25 = RG_rl_196 ;
	7'h4d :
		TR_25 = RG_rl_196 ;
	7'h4e :
		TR_25 = RG_rl_196 ;
	7'h4f :
		TR_25 = RG_rl_196 ;
	7'h50 :
		TR_25 = RG_rl_196 ;
	7'h51 :
		TR_25 = RG_rl_196 ;
	7'h52 :
		TR_25 = RG_rl_196 ;
	7'h53 :
		TR_25 = RG_rl_196 ;
	7'h54 :
		TR_25 = RG_rl_196 ;
	7'h55 :
		TR_25 = RG_rl_196 ;
	7'h56 :
		TR_25 = RG_rl_196 ;
	7'h57 :
		TR_25 = RG_rl_196 ;
	7'h58 :
		TR_25 = RG_rl_196 ;
	7'h59 :
		TR_25 = RG_rl_196 ;
	7'h5a :
		TR_25 = RG_rl_196 ;
	7'h5b :
		TR_25 = RG_rl_196 ;
	7'h5c :
		TR_25 = RG_rl_196 ;
	7'h5d :
		TR_25 = RG_rl_196 ;
	7'h5e :
		TR_25 = RG_rl_196 ;
	7'h5f :
		TR_25 = RG_rl_196 ;
	7'h60 :
		TR_25 = RG_rl_196 ;
	7'h61 :
		TR_25 = RG_rl_196 ;
	7'h62 :
		TR_25 = RG_rl_196 ;
	7'h63 :
		TR_25 = RG_rl_196 ;
	7'h64 :
		TR_25 = RG_rl_196 ;
	7'h65 :
		TR_25 = RG_rl_196 ;
	7'h66 :
		TR_25 = RG_rl_196 ;
	7'h67 :
		TR_25 = RG_rl_196 ;
	7'h68 :
		TR_25 = RG_rl_196 ;
	7'h69 :
		TR_25 = RG_rl_196 ;
	7'h6a :
		TR_25 = RG_rl_196 ;
	7'h6b :
		TR_25 = RG_rl_196 ;
	7'h6c :
		TR_25 = RG_rl_196 ;
	7'h6d :
		TR_25 = RG_rl_196 ;
	7'h6e :
		TR_25 = RG_rl_196 ;
	7'h6f :
		TR_25 = RG_rl_196 ;
	7'h70 :
		TR_25 = RG_rl_196 ;
	7'h71 :
		TR_25 = RG_rl_196 ;
	7'h72 :
		TR_25 = RG_rl_196 ;
	7'h73 :
		TR_25 = RG_rl_196 ;
	7'h74 :
		TR_25 = RG_rl_196 ;
	7'h75 :
		TR_25 = RG_rl_196 ;
	7'h76 :
		TR_25 = RG_rl_196 ;
	7'h77 :
		TR_25 = RG_rl_196 ;
	7'h78 :
		TR_25 = RG_rl_196 ;
	7'h79 :
		TR_25 = RG_rl_196 ;
	7'h7a :
		TR_25 = RG_rl_196 ;
	7'h7b :
		TR_25 = RG_rl_196 ;
	7'h7c :
		TR_25 = RG_rl_196 ;
	7'h7d :
		TR_25 = RG_rl_196 ;
	7'h7e :
		TR_25 = RG_rl_196 ;
	7'h7f :
		TR_25 = RG_rl_196 ;
	default :
		TR_25 = 9'hx ;
	endcase
always @ ( RG_rl_197 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_26 = RG_rl_197 ;
	7'h01 :
		TR_26 = RG_rl_197 ;
	7'h02 :
		TR_26 = RG_rl_197 ;
	7'h03 :
		TR_26 = RG_rl_197 ;
	7'h04 :
		TR_26 = RG_rl_197 ;
	7'h05 :
		TR_26 = RG_rl_197 ;
	7'h06 :
		TR_26 = RG_rl_197 ;
	7'h07 :
		TR_26 = RG_rl_197 ;
	7'h08 :
		TR_26 = RG_rl_197 ;
	7'h09 :
		TR_26 = RG_rl_197 ;
	7'h0a :
		TR_26 = RG_rl_197 ;
	7'h0b :
		TR_26 = RG_rl_197 ;
	7'h0c :
		TR_26 = RG_rl_197 ;
	7'h0d :
		TR_26 = RG_rl_197 ;
	7'h0e :
		TR_26 = 9'h000 ;	// line#=../rle.cpp:68
	7'h0f :
		TR_26 = RG_rl_197 ;
	7'h10 :
		TR_26 = RG_rl_197 ;
	7'h11 :
		TR_26 = RG_rl_197 ;
	7'h12 :
		TR_26 = RG_rl_197 ;
	7'h13 :
		TR_26 = RG_rl_197 ;
	7'h14 :
		TR_26 = RG_rl_197 ;
	7'h15 :
		TR_26 = RG_rl_197 ;
	7'h16 :
		TR_26 = RG_rl_197 ;
	7'h17 :
		TR_26 = RG_rl_197 ;
	7'h18 :
		TR_26 = RG_rl_197 ;
	7'h19 :
		TR_26 = RG_rl_197 ;
	7'h1a :
		TR_26 = RG_rl_197 ;
	7'h1b :
		TR_26 = RG_rl_197 ;
	7'h1c :
		TR_26 = RG_rl_197 ;
	7'h1d :
		TR_26 = RG_rl_197 ;
	7'h1e :
		TR_26 = RG_rl_197 ;
	7'h1f :
		TR_26 = RG_rl_197 ;
	7'h20 :
		TR_26 = RG_rl_197 ;
	7'h21 :
		TR_26 = RG_rl_197 ;
	7'h22 :
		TR_26 = RG_rl_197 ;
	7'h23 :
		TR_26 = RG_rl_197 ;
	7'h24 :
		TR_26 = RG_rl_197 ;
	7'h25 :
		TR_26 = RG_rl_197 ;
	7'h26 :
		TR_26 = RG_rl_197 ;
	7'h27 :
		TR_26 = RG_rl_197 ;
	7'h28 :
		TR_26 = RG_rl_197 ;
	7'h29 :
		TR_26 = RG_rl_197 ;
	7'h2a :
		TR_26 = RG_rl_197 ;
	7'h2b :
		TR_26 = RG_rl_197 ;
	7'h2c :
		TR_26 = RG_rl_197 ;
	7'h2d :
		TR_26 = RG_rl_197 ;
	7'h2e :
		TR_26 = RG_rl_197 ;
	7'h2f :
		TR_26 = RG_rl_197 ;
	7'h30 :
		TR_26 = RG_rl_197 ;
	7'h31 :
		TR_26 = RG_rl_197 ;
	7'h32 :
		TR_26 = RG_rl_197 ;
	7'h33 :
		TR_26 = RG_rl_197 ;
	7'h34 :
		TR_26 = RG_rl_197 ;
	7'h35 :
		TR_26 = RG_rl_197 ;
	7'h36 :
		TR_26 = RG_rl_197 ;
	7'h37 :
		TR_26 = RG_rl_197 ;
	7'h38 :
		TR_26 = RG_rl_197 ;
	7'h39 :
		TR_26 = RG_rl_197 ;
	7'h3a :
		TR_26 = RG_rl_197 ;
	7'h3b :
		TR_26 = RG_rl_197 ;
	7'h3c :
		TR_26 = RG_rl_197 ;
	7'h3d :
		TR_26 = RG_rl_197 ;
	7'h3e :
		TR_26 = RG_rl_197 ;
	7'h3f :
		TR_26 = RG_rl_197 ;
	7'h40 :
		TR_26 = RG_rl_197 ;
	7'h41 :
		TR_26 = RG_rl_197 ;
	7'h42 :
		TR_26 = RG_rl_197 ;
	7'h43 :
		TR_26 = RG_rl_197 ;
	7'h44 :
		TR_26 = RG_rl_197 ;
	7'h45 :
		TR_26 = RG_rl_197 ;
	7'h46 :
		TR_26 = RG_rl_197 ;
	7'h47 :
		TR_26 = RG_rl_197 ;
	7'h48 :
		TR_26 = RG_rl_197 ;
	7'h49 :
		TR_26 = RG_rl_197 ;
	7'h4a :
		TR_26 = RG_rl_197 ;
	7'h4b :
		TR_26 = RG_rl_197 ;
	7'h4c :
		TR_26 = RG_rl_197 ;
	7'h4d :
		TR_26 = RG_rl_197 ;
	7'h4e :
		TR_26 = RG_rl_197 ;
	7'h4f :
		TR_26 = RG_rl_197 ;
	7'h50 :
		TR_26 = RG_rl_197 ;
	7'h51 :
		TR_26 = RG_rl_197 ;
	7'h52 :
		TR_26 = RG_rl_197 ;
	7'h53 :
		TR_26 = RG_rl_197 ;
	7'h54 :
		TR_26 = RG_rl_197 ;
	7'h55 :
		TR_26 = RG_rl_197 ;
	7'h56 :
		TR_26 = RG_rl_197 ;
	7'h57 :
		TR_26 = RG_rl_197 ;
	7'h58 :
		TR_26 = RG_rl_197 ;
	7'h59 :
		TR_26 = RG_rl_197 ;
	7'h5a :
		TR_26 = RG_rl_197 ;
	7'h5b :
		TR_26 = RG_rl_197 ;
	7'h5c :
		TR_26 = RG_rl_197 ;
	7'h5d :
		TR_26 = RG_rl_197 ;
	7'h5e :
		TR_26 = RG_rl_197 ;
	7'h5f :
		TR_26 = RG_rl_197 ;
	7'h60 :
		TR_26 = RG_rl_197 ;
	7'h61 :
		TR_26 = RG_rl_197 ;
	7'h62 :
		TR_26 = RG_rl_197 ;
	7'h63 :
		TR_26 = RG_rl_197 ;
	7'h64 :
		TR_26 = RG_rl_197 ;
	7'h65 :
		TR_26 = RG_rl_197 ;
	7'h66 :
		TR_26 = RG_rl_197 ;
	7'h67 :
		TR_26 = RG_rl_197 ;
	7'h68 :
		TR_26 = RG_rl_197 ;
	7'h69 :
		TR_26 = RG_rl_197 ;
	7'h6a :
		TR_26 = RG_rl_197 ;
	7'h6b :
		TR_26 = RG_rl_197 ;
	7'h6c :
		TR_26 = RG_rl_197 ;
	7'h6d :
		TR_26 = RG_rl_197 ;
	7'h6e :
		TR_26 = RG_rl_197 ;
	7'h6f :
		TR_26 = RG_rl_197 ;
	7'h70 :
		TR_26 = RG_rl_197 ;
	7'h71 :
		TR_26 = RG_rl_197 ;
	7'h72 :
		TR_26 = RG_rl_197 ;
	7'h73 :
		TR_26 = RG_rl_197 ;
	7'h74 :
		TR_26 = RG_rl_197 ;
	7'h75 :
		TR_26 = RG_rl_197 ;
	7'h76 :
		TR_26 = RG_rl_197 ;
	7'h77 :
		TR_26 = RG_rl_197 ;
	7'h78 :
		TR_26 = RG_rl_197 ;
	7'h79 :
		TR_26 = RG_rl_197 ;
	7'h7a :
		TR_26 = RG_rl_197 ;
	7'h7b :
		TR_26 = RG_rl_197 ;
	7'h7c :
		TR_26 = RG_rl_197 ;
	7'h7d :
		TR_26 = RG_rl_197 ;
	7'h7e :
		TR_26 = RG_rl_197 ;
	7'h7f :
		TR_26 = RG_rl_197 ;
	default :
		TR_26 = 9'hx ;
	endcase
always @ ( RG_rl_198 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_27 = RG_rl_198 ;
	7'h01 :
		TR_27 = RG_rl_198 ;
	7'h02 :
		TR_27 = RG_rl_198 ;
	7'h03 :
		TR_27 = RG_rl_198 ;
	7'h04 :
		TR_27 = RG_rl_198 ;
	7'h05 :
		TR_27 = RG_rl_198 ;
	7'h06 :
		TR_27 = RG_rl_198 ;
	7'h07 :
		TR_27 = RG_rl_198 ;
	7'h08 :
		TR_27 = RG_rl_198 ;
	7'h09 :
		TR_27 = RG_rl_198 ;
	7'h0a :
		TR_27 = RG_rl_198 ;
	7'h0b :
		TR_27 = RG_rl_198 ;
	7'h0c :
		TR_27 = RG_rl_198 ;
	7'h0d :
		TR_27 = RG_rl_198 ;
	7'h0e :
		TR_27 = RG_rl_198 ;
	7'h0f :
		TR_27 = 9'h000 ;	// line#=../rle.cpp:68
	7'h10 :
		TR_27 = RG_rl_198 ;
	7'h11 :
		TR_27 = RG_rl_198 ;
	7'h12 :
		TR_27 = RG_rl_198 ;
	7'h13 :
		TR_27 = RG_rl_198 ;
	7'h14 :
		TR_27 = RG_rl_198 ;
	7'h15 :
		TR_27 = RG_rl_198 ;
	7'h16 :
		TR_27 = RG_rl_198 ;
	7'h17 :
		TR_27 = RG_rl_198 ;
	7'h18 :
		TR_27 = RG_rl_198 ;
	7'h19 :
		TR_27 = RG_rl_198 ;
	7'h1a :
		TR_27 = RG_rl_198 ;
	7'h1b :
		TR_27 = RG_rl_198 ;
	7'h1c :
		TR_27 = RG_rl_198 ;
	7'h1d :
		TR_27 = RG_rl_198 ;
	7'h1e :
		TR_27 = RG_rl_198 ;
	7'h1f :
		TR_27 = RG_rl_198 ;
	7'h20 :
		TR_27 = RG_rl_198 ;
	7'h21 :
		TR_27 = RG_rl_198 ;
	7'h22 :
		TR_27 = RG_rl_198 ;
	7'h23 :
		TR_27 = RG_rl_198 ;
	7'h24 :
		TR_27 = RG_rl_198 ;
	7'h25 :
		TR_27 = RG_rl_198 ;
	7'h26 :
		TR_27 = RG_rl_198 ;
	7'h27 :
		TR_27 = RG_rl_198 ;
	7'h28 :
		TR_27 = RG_rl_198 ;
	7'h29 :
		TR_27 = RG_rl_198 ;
	7'h2a :
		TR_27 = RG_rl_198 ;
	7'h2b :
		TR_27 = RG_rl_198 ;
	7'h2c :
		TR_27 = RG_rl_198 ;
	7'h2d :
		TR_27 = RG_rl_198 ;
	7'h2e :
		TR_27 = RG_rl_198 ;
	7'h2f :
		TR_27 = RG_rl_198 ;
	7'h30 :
		TR_27 = RG_rl_198 ;
	7'h31 :
		TR_27 = RG_rl_198 ;
	7'h32 :
		TR_27 = RG_rl_198 ;
	7'h33 :
		TR_27 = RG_rl_198 ;
	7'h34 :
		TR_27 = RG_rl_198 ;
	7'h35 :
		TR_27 = RG_rl_198 ;
	7'h36 :
		TR_27 = RG_rl_198 ;
	7'h37 :
		TR_27 = RG_rl_198 ;
	7'h38 :
		TR_27 = RG_rl_198 ;
	7'h39 :
		TR_27 = RG_rl_198 ;
	7'h3a :
		TR_27 = RG_rl_198 ;
	7'h3b :
		TR_27 = RG_rl_198 ;
	7'h3c :
		TR_27 = RG_rl_198 ;
	7'h3d :
		TR_27 = RG_rl_198 ;
	7'h3e :
		TR_27 = RG_rl_198 ;
	7'h3f :
		TR_27 = RG_rl_198 ;
	7'h40 :
		TR_27 = RG_rl_198 ;
	7'h41 :
		TR_27 = RG_rl_198 ;
	7'h42 :
		TR_27 = RG_rl_198 ;
	7'h43 :
		TR_27 = RG_rl_198 ;
	7'h44 :
		TR_27 = RG_rl_198 ;
	7'h45 :
		TR_27 = RG_rl_198 ;
	7'h46 :
		TR_27 = RG_rl_198 ;
	7'h47 :
		TR_27 = RG_rl_198 ;
	7'h48 :
		TR_27 = RG_rl_198 ;
	7'h49 :
		TR_27 = RG_rl_198 ;
	7'h4a :
		TR_27 = RG_rl_198 ;
	7'h4b :
		TR_27 = RG_rl_198 ;
	7'h4c :
		TR_27 = RG_rl_198 ;
	7'h4d :
		TR_27 = RG_rl_198 ;
	7'h4e :
		TR_27 = RG_rl_198 ;
	7'h4f :
		TR_27 = RG_rl_198 ;
	7'h50 :
		TR_27 = RG_rl_198 ;
	7'h51 :
		TR_27 = RG_rl_198 ;
	7'h52 :
		TR_27 = RG_rl_198 ;
	7'h53 :
		TR_27 = RG_rl_198 ;
	7'h54 :
		TR_27 = RG_rl_198 ;
	7'h55 :
		TR_27 = RG_rl_198 ;
	7'h56 :
		TR_27 = RG_rl_198 ;
	7'h57 :
		TR_27 = RG_rl_198 ;
	7'h58 :
		TR_27 = RG_rl_198 ;
	7'h59 :
		TR_27 = RG_rl_198 ;
	7'h5a :
		TR_27 = RG_rl_198 ;
	7'h5b :
		TR_27 = RG_rl_198 ;
	7'h5c :
		TR_27 = RG_rl_198 ;
	7'h5d :
		TR_27 = RG_rl_198 ;
	7'h5e :
		TR_27 = RG_rl_198 ;
	7'h5f :
		TR_27 = RG_rl_198 ;
	7'h60 :
		TR_27 = RG_rl_198 ;
	7'h61 :
		TR_27 = RG_rl_198 ;
	7'h62 :
		TR_27 = RG_rl_198 ;
	7'h63 :
		TR_27 = RG_rl_198 ;
	7'h64 :
		TR_27 = RG_rl_198 ;
	7'h65 :
		TR_27 = RG_rl_198 ;
	7'h66 :
		TR_27 = RG_rl_198 ;
	7'h67 :
		TR_27 = RG_rl_198 ;
	7'h68 :
		TR_27 = RG_rl_198 ;
	7'h69 :
		TR_27 = RG_rl_198 ;
	7'h6a :
		TR_27 = RG_rl_198 ;
	7'h6b :
		TR_27 = RG_rl_198 ;
	7'h6c :
		TR_27 = RG_rl_198 ;
	7'h6d :
		TR_27 = RG_rl_198 ;
	7'h6e :
		TR_27 = RG_rl_198 ;
	7'h6f :
		TR_27 = RG_rl_198 ;
	7'h70 :
		TR_27 = RG_rl_198 ;
	7'h71 :
		TR_27 = RG_rl_198 ;
	7'h72 :
		TR_27 = RG_rl_198 ;
	7'h73 :
		TR_27 = RG_rl_198 ;
	7'h74 :
		TR_27 = RG_rl_198 ;
	7'h75 :
		TR_27 = RG_rl_198 ;
	7'h76 :
		TR_27 = RG_rl_198 ;
	7'h77 :
		TR_27 = RG_rl_198 ;
	7'h78 :
		TR_27 = RG_rl_198 ;
	7'h79 :
		TR_27 = RG_rl_198 ;
	7'h7a :
		TR_27 = RG_rl_198 ;
	7'h7b :
		TR_27 = RG_rl_198 ;
	7'h7c :
		TR_27 = RG_rl_198 ;
	7'h7d :
		TR_27 = RG_rl_198 ;
	7'h7e :
		TR_27 = RG_rl_198 ;
	7'h7f :
		TR_27 = RG_rl_198 ;
	default :
		TR_27 = 9'hx ;
	endcase
always @ ( RG_rl_199 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_28 = RG_rl_199 ;
	7'h01 :
		TR_28 = RG_rl_199 ;
	7'h02 :
		TR_28 = RG_rl_199 ;
	7'h03 :
		TR_28 = RG_rl_199 ;
	7'h04 :
		TR_28 = RG_rl_199 ;
	7'h05 :
		TR_28 = RG_rl_199 ;
	7'h06 :
		TR_28 = RG_rl_199 ;
	7'h07 :
		TR_28 = RG_rl_199 ;
	7'h08 :
		TR_28 = RG_rl_199 ;
	7'h09 :
		TR_28 = RG_rl_199 ;
	7'h0a :
		TR_28 = RG_rl_199 ;
	7'h0b :
		TR_28 = RG_rl_199 ;
	7'h0c :
		TR_28 = RG_rl_199 ;
	7'h0d :
		TR_28 = RG_rl_199 ;
	7'h0e :
		TR_28 = RG_rl_199 ;
	7'h0f :
		TR_28 = RG_rl_199 ;
	7'h10 :
		TR_28 = 9'h000 ;	// line#=../rle.cpp:68
	7'h11 :
		TR_28 = RG_rl_199 ;
	7'h12 :
		TR_28 = RG_rl_199 ;
	7'h13 :
		TR_28 = RG_rl_199 ;
	7'h14 :
		TR_28 = RG_rl_199 ;
	7'h15 :
		TR_28 = RG_rl_199 ;
	7'h16 :
		TR_28 = RG_rl_199 ;
	7'h17 :
		TR_28 = RG_rl_199 ;
	7'h18 :
		TR_28 = RG_rl_199 ;
	7'h19 :
		TR_28 = RG_rl_199 ;
	7'h1a :
		TR_28 = RG_rl_199 ;
	7'h1b :
		TR_28 = RG_rl_199 ;
	7'h1c :
		TR_28 = RG_rl_199 ;
	7'h1d :
		TR_28 = RG_rl_199 ;
	7'h1e :
		TR_28 = RG_rl_199 ;
	7'h1f :
		TR_28 = RG_rl_199 ;
	7'h20 :
		TR_28 = RG_rl_199 ;
	7'h21 :
		TR_28 = RG_rl_199 ;
	7'h22 :
		TR_28 = RG_rl_199 ;
	7'h23 :
		TR_28 = RG_rl_199 ;
	7'h24 :
		TR_28 = RG_rl_199 ;
	7'h25 :
		TR_28 = RG_rl_199 ;
	7'h26 :
		TR_28 = RG_rl_199 ;
	7'h27 :
		TR_28 = RG_rl_199 ;
	7'h28 :
		TR_28 = RG_rl_199 ;
	7'h29 :
		TR_28 = RG_rl_199 ;
	7'h2a :
		TR_28 = RG_rl_199 ;
	7'h2b :
		TR_28 = RG_rl_199 ;
	7'h2c :
		TR_28 = RG_rl_199 ;
	7'h2d :
		TR_28 = RG_rl_199 ;
	7'h2e :
		TR_28 = RG_rl_199 ;
	7'h2f :
		TR_28 = RG_rl_199 ;
	7'h30 :
		TR_28 = RG_rl_199 ;
	7'h31 :
		TR_28 = RG_rl_199 ;
	7'h32 :
		TR_28 = RG_rl_199 ;
	7'h33 :
		TR_28 = RG_rl_199 ;
	7'h34 :
		TR_28 = RG_rl_199 ;
	7'h35 :
		TR_28 = RG_rl_199 ;
	7'h36 :
		TR_28 = RG_rl_199 ;
	7'h37 :
		TR_28 = RG_rl_199 ;
	7'h38 :
		TR_28 = RG_rl_199 ;
	7'h39 :
		TR_28 = RG_rl_199 ;
	7'h3a :
		TR_28 = RG_rl_199 ;
	7'h3b :
		TR_28 = RG_rl_199 ;
	7'h3c :
		TR_28 = RG_rl_199 ;
	7'h3d :
		TR_28 = RG_rl_199 ;
	7'h3e :
		TR_28 = RG_rl_199 ;
	7'h3f :
		TR_28 = RG_rl_199 ;
	7'h40 :
		TR_28 = RG_rl_199 ;
	7'h41 :
		TR_28 = RG_rl_199 ;
	7'h42 :
		TR_28 = RG_rl_199 ;
	7'h43 :
		TR_28 = RG_rl_199 ;
	7'h44 :
		TR_28 = RG_rl_199 ;
	7'h45 :
		TR_28 = RG_rl_199 ;
	7'h46 :
		TR_28 = RG_rl_199 ;
	7'h47 :
		TR_28 = RG_rl_199 ;
	7'h48 :
		TR_28 = RG_rl_199 ;
	7'h49 :
		TR_28 = RG_rl_199 ;
	7'h4a :
		TR_28 = RG_rl_199 ;
	7'h4b :
		TR_28 = RG_rl_199 ;
	7'h4c :
		TR_28 = RG_rl_199 ;
	7'h4d :
		TR_28 = RG_rl_199 ;
	7'h4e :
		TR_28 = RG_rl_199 ;
	7'h4f :
		TR_28 = RG_rl_199 ;
	7'h50 :
		TR_28 = RG_rl_199 ;
	7'h51 :
		TR_28 = RG_rl_199 ;
	7'h52 :
		TR_28 = RG_rl_199 ;
	7'h53 :
		TR_28 = RG_rl_199 ;
	7'h54 :
		TR_28 = RG_rl_199 ;
	7'h55 :
		TR_28 = RG_rl_199 ;
	7'h56 :
		TR_28 = RG_rl_199 ;
	7'h57 :
		TR_28 = RG_rl_199 ;
	7'h58 :
		TR_28 = RG_rl_199 ;
	7'h59 :
		TR_28 = RG_rl_199 ;
	7'h5a :
		TR_28 = RG_rl_199 ;
	7'h5b :
		TR_28 = RG_rl_199 ;
	7'h5c :
		TR_28 = RG_rl_199 ;
	7'h5d :
		TR_28 = RG_rl_199 ;
	7'h5e :
		TR_28 = RG_rl_199 ;
	7'h5f :
		TR_28 = RG_rl_199 ;
	7'h60 :
		TR_28 = RG_rl_199 ;
	7'h61 :
		TR_28 = RG_rl_199 ;
	7'h62 :
		TR_28 = RG_rl_199 ;
	7'h63 :
		TR_28 = RG_rl_199 ;
	7'h64 :
		TR_28 = RG_rl_199 ;
	7'h65 :
		TR_28 = RG_rl_199 ;
	7'h66 :
		TR_28 = RG_rl_199 ;
	7'h67 :
		TR_28 = RG_rl_199 ;
	7'h68 :
		TR_28 = RG_rl_199 ;
	7'h69 :
		TR_28 = RG_rl_199 ;
	7'h6a :
		TR_28 = RG_rl_199 ;
	7'h6b :
		TR_28 = RG_rl_199 ;
	7'h6c :
		TR_28 = RG_rl_199 ;
	7'h6d :
		TR_28 = RG_rl_199 ;
	7'h6e :
		TR_28 = RG_rl_199 ;
	7'h6f :
		TR_28 = RG_rl_199 ;
	7'h70 :
		TR_28 = RG_rl_199 ;
	7'h71 :
		TR_28 = RG_rl_199 ;
	7'h72 :
		TR_28 = RG_rl_199 ;
	7'h73 :
		TR_28 = RG_rl_199 ;
	7'h74 :
		TR_28 = RG_rl_199 ;
	7'h75 :
		TR_28 = RG_rl_199 ;
	7'h76 :
		TR_28 = RG_rl_199 ;
	7'h77 :
		TR_28 = RG_rl_199 ;
	7'h78 :
		TR_28 = RG_rl_199 ;
	7'h79 :
		TR_28 = RG_rl_199 ;
	7'h7a :
		TR_28 = RG_rl_199 ;
	7'h7b :
		TR_28 = RG_rl_199 ;
	7'h7c :
		TR_28 = RG_rl_199 ;
	7'h7d :
		TR_28 = RG_rl_199 ;
	7'h7e :
		TR_28 = RG_rl_199 ;
	7'h7f :
		TR_28 = RG_rl_199 ;
	default :
		TR_28 = 9'hx ;
	endcase
always @ ( RG_rl_200 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_29 = RG_rl_200 ;
	7'h01 :
		TR_29 = RG_rl_200 ;
	7'h02 :
		TR_29 = RG_rl_200 ;
	7'h03 :
		TR_29 = RG_rl_200 ;
	7'h04 :
		TR_29 = RG_rl_200 ;
	7'h05 :
		TR_29 = RG_rl_200 ;
	7'h06 :
		TR_29 = RG_rl_200 ;
	7'h07 :
		TR_29 = RG_rl_200 ;
	7'h08 :
		TR_29 = RG_rl_200 ;
	7'h09 :
		TR_29 = RG_rl_200 ;
	7'h0a :
		TR_29 = RG_rl_200 ;
	7'h0b :
		TR_29 = RG_rl_200 ;
	7'h0c :
		TR_29 = RG_rl_200 ;
	7'h0d :
		TR_29 = RG_rl_200 ;
	7'h0e :
		TR_29 = RG_rl_200 ;
	7'h0f :
		TR_29 = RG_rl_200 ;
	7'h10 :
		TR_29 = RG_rl_200 ;
	7'h11 :
		TR_29 = 9'h000 ;	// line#=../rle.cpp:68
	7'h12 :
		TR_29 = RG_rl_200 ;
	7'h13 :
		TR_29 = RG_rl_200 ;
	7'h14 :
		TR_29 = RG_rl_200 ;
	7'h15 :
		TR_29 = RG_rl_200 ;
	7'h16 :
		TR_29 = RG_rl_200 ;
	7'h17 :
		TR_29 = RG_rl_200 ;
	7'h18 :
		TR_29 = RG_rl_200 ;
	7'h19 :
		TR_29 = RG_rl_200 ;
	7'h1a :
		TR_29 = RG_rl_200 ;
	7'h1b :
		TR_29 = RG_rl_200 ;
	7'h1c :
		TR_29 = RG_rl_200 ;
	7'h1d :
		TR_29 = RG_rl_200 ;
	7'h1e :
		TR_29 = RG_rl_200 ;
	7'h1f :
		TR_29 = RG_rl_200 ;
	7'h20 :
		TR_29 = RG_rl_200 ;
	7'h21 :
		TR_29 = RG_rl_200 ;
	7'h22 :
		TR_29 = RG_rl_200 ;
	7'h23 :
		TR_29 = RG_rl_200 ;
	7'h24 :
		TR_29 = RG_rl_200 ;
	7'h25 :
		TR_29 = RG_rl_200 ;
	7'h26 :
		TR_29 = RG_rl_200 ;
	7'h27 :
		TR_29 = RG_rl_200 ;
	7'h28 :
		TR_29 = RG_rl_200 ;
	7'h29 :
		TR_29 = RG_rl_200 ;
	7'h2a :
		TR_29 = RG_rl_200 ;
	7'h2b :
		TR_29 = RG_rl_200 ;
	7'h2c :
		TR_29 = RG_rl_200 ;
	7'h2d :
		TR_29 = RG_rl_200 ;
	7'h2e :
		TR_29 = RG_rl_200 ;
	7'h2f :
		TR_29 = RG_rl_200 ;
	7'h30 :
		TR_29 = RG_rl_200 ;
	7'h31 :
		TR_29 = RG_rl_200 ;
	7'h32 :
		TR_29 = RG_rl_200 ;
	7'h33 :
		TR_29 = RG_rl_200 ;
	7'h34 :
		TR_29 = RG_rl_200 ;
	7'h35 :
		TR_29 = RG_rl_200 ;
	7'h36 :
		TR_29 = RG_rl_200 ;
	7'h37 :
		TR_29 = RG_rl_200 ;
	7'h38 :
		TR_29 = RG_rl_200 ;
	7'h39 :
		TR_29 = RG_rl_200 ;
	7'h3a :
		TR_29 = RG_rl_200 ;
	7'h3b :
		TR_29 = RG_rl_200 ;
	7'h3c :
		TR_29 = RG_rl_200 ;
	7'h3d :
		TR_29 = RG_rl_200 ;
	7'h3e :
		TR_29 = RG_rl_200 ;
	7'h3f :
		TR_29 = RG_rl_200 ;
	7'h40 :
		TR_29 = RG_rl_200 ;
	7'h41 :
		TR_29 = RG_rl_200 ;
	7'h42 :
		TR_29 = RG_rl_200 ;
	7'h43 :
		TR_29 = RG_rl_200 ;
	7'h44 :
		TR_29 = RG_rl_200 ;
	7'h45 :
		TR_29 = RG_rl_200 ;
	7'h46 :
		TR_29 = RG_rl_200 ;
	7'h47 :
		TR_29 = RG_rl_200 ;
	7'h48 :
		TR_29 = RG_rl_200 ;
	7'h49 :
		TR_29 = RG_rl_200 ;
	7'h4a :
		TR_29 = RG_rl_200 ;
	7'h4b :
		TR_29 = RG_rl_200 ;
	7'h4c :
		TR_29 = RG_rl_200 ;
	7'h4d :
		TR_29 = RG_rl_200 ;
	7'h4e :
		TR_29 = RG_rl_200 ;
	7'h4f :
		TR_29 = RG_rl_200 ;
	7'h50 :
		TR_29 = RG_rl_200 ;
	7'h51 :
		TR_29 = RG_rl_200 ;
	7'h52 :
		TR_29 = RG_rl_200 ;
	7'h53 :
		TR_29 = RG_rl_200 ;
	7'h54 :
		TR_29 = RG_rl_200 ;
	7'h55 :
		TR_29 = RG_rl_200 ;
	7'h56 :
		TR_29 = RG_rl_200 ;
	7'h57 :
		TR_29 = RG_rl_200 ;
	7'h58 :
		TR_29 = RG_rl_200 ;
	7'h59 :
		TR_29 = RG_rl_200 ;
	7'h5a :
		TR_29 = RG_rl_200 ;
	7'h5b :
		TR_29 = RG_rl_200 ;
	7'h5c :
		TR_29 = RG_rl_200 ;
	7'h5d :
		TR_29 = RG_rl_200 ;
	7'h5e :
		TR_29 = RG_rl_200 ;
	7'h5f :
		TR_29 = RG_rl_200 ;
	7'h60 :
		TR_29 = RG_rl_200 ;
	7'h61 :
		TR_29 = RG_rl_200 ;
	7'h62 :
		TR_29 = RG_rl_200 ;
	7'h63 :
		TR_29 = RG_rl_200 ;
	7'h64 :
		TR_29 = RG_rl_200 ;
	7'h65 :
		TR_29 = RG_rl_200 ;
	7'h66 :
		TR_29 = RG_rl_200 ;
	7'h67 :
		TR_29 = RG_rl_200 ;
	7'h68 :
		TR_29 = RG_rl_200 ;
	7'h69 :
		TR_29 = RG_rl_200 ;
	7'h6a :
		TR_29 = RG_rl_200 ;
	7'h6b :
		TR_29 = RG_rl_200 ;
	7'h6c :
		TR_29 = RG_rl_200 ;
	7'h6d :
		TR_29 = RG_rl_200 ;
	7'h6e :
		TR_29 = RG_rl_200 ;
	7'h6f :
		TR_29 = RG_rl_200 ;
	7'h70 :
		TR_29 = RG_rl_200 ;
	7'h71 :
		TR_29 = RG_rl_200 ;
	7'h72 :
		TR_29 = RG_rl_200 ;
	7'h73 :
		TR_29 = RG_rl_200 ;
	7'h74 :
		TR_29 = RG_rl_200 ;
	7'h75 :
		TR_29 = RG_rl_200 ;
	7'h76 :
		TR_29 = RG_rl_200 ;
	7'h77 :
		TR_29 = RG_rl_200 ;
	7'h78 :
		TR_29 = RG_rl_200 ;
	7'h79 :
		TR_29 = RG_rl_200 ;
	7'h7a :
		TR_29 = RG_rl_200 ;
	7'h7b :
		TR_29 = RG_rl_200 ;
	7'h7c :
		TR_29 = RG_rl_200 ;
	7'h7d :
		TR_29 = RG_rl_200 ;
	7'h7e :
		TR_29 = RG_rl_200 ;
	7'h7f :
		TR_29 = RG_rl_200 ;
	default :
		TR_29 = 9'hx ;
	endcase
always @ ( RG_rl_201 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_30 = RG_rl_201 ;
	7'h01 :
		TR_30 = RG_rl_201 ;
	7'h02 :
		TR_30 = RG_rl_201 ;
	7'h03 :
		TR_30 = RG_rl_201 ;
	7'h04 :
		TR_30 = RG_rl_201 ;
	7'h05 :
		TR_30 = RG_rl_201 ;
	7'h06 :
		TR_30 = RG_rl_201 ;
	7'h07 :
		TR_30 = RG_rl_201 ;
	7'h08 :
		TR_30 = RG_rl_201 ;
	7'h09 :
		TR_30 = RG_rl_201 ;
	7'h0a :
		TR_30 = RG_rl_201 ;
	7'h0b :
		TR_30 = RG_rl_201 ;
	7'h0c :
		TR_30 = RG_rl_201 ;
	7'h0d :
		TR_30 = RG_rl_201 ;
	7'h0e :
		TR_30 = RG_rl_201 ;
	7'h0f :
		TR_30 = RG_rl_201 ;
	7'h10 :
		TR_30 = RG_rl_201 ;
	7'h11 :
		TR_30 = RG_rl_201 ;
	7'h12 :
		TR_30 = 9'h000 ;	// line#=../rle.cpp:68
	7'h13 :
		TR_30 = RG_rl_201 ;
	7'h14 :
		TR_30 = RG_rl_201 ;
	7'h15 :
		TR_30 = RG_rl_201 ;
	7'h16 :
		TR_30 = RG_rl_201 ;
	7'h17 :
		TR_30 = RG_rl_201 ;
	7'h18 :
		TR_30 = RG_rl_201 ;
	7'h19 :
		TR_30 = RG_rl_201 ;
	7'h1a :
		TR_30 = RG_rl_201 ;
	7'h1b :
		TR_30 = RG_rl_201 ;
	7'h1c :
		TR_30 = RG_rl_201 ;
	7'h1d :
		TR_30 = RG_rl_201 ;
	7'h1e :
		TR_30 = RG_rl_201 ;
	7'h1f :
		TR_30 = RG_rl_201 ;
	7'h20 :
		TR_30 = RG_rl_201 ;
	7'h21 :
		TR_30 = RG_rl_201 ;
	7'h22 :
		TR_30 = RG_rl_201 ;
	7'h23 :
		TR_30 = RG_rl_201 ;
	7'h24 :
		TR_30 = RG_rl_201 ;
	7'h25 :
		TR_30 = RG_rl_201 ;
	7'h26 :
		TR_30 = RG_rl_201 ;
	7'h27 :
		TR_30 = RG_rl_201 ;
	7'h28 :
		TR_30 = RG_rl_201 ;
	7'h29 :
		TR_30 = RG_rl_201 ;
	7'h2a :
		TR_30 = RG_rl_201 ;
	7'h2b :
		TR_30 = RG_rl_201 ;
	7'h2c :
		TR_30 = RG_rl_201 ;
	7'h2d :
		TR_30 = RG_rl_201 ;
	7'h2e :
		TR_30 = RG_rl_201 ;
	7'h2f :
		TR_30 = RG_rl_201 ;
	7'h30 :
		TR_30 = RG_rl_201 ;
	7'h31 :
		TR_30 = RG_rl_201 ;
	7'h32 :
		TR_30 = RG_rl_201 ;
	7'h33 :
		TR_30 = RG_rl_201 ;
	7'h34 :
		TR_30 = RG_rl_201 ;
	7'h35 :
		TR_30 = RG_rl_201 ;
	7'h36 :
		TR_30 = RG_rl_201 ;
	7'h37 :
		TR_30 = RG_rl_201 ;
	7'h38 :
		TR_30 = RG_rl_201 ;
	7'h39 :
		TR_30 = RG_rl_201 ;
	7'h3a :
		TR_30 = RG_rl_201 ;
	7'h3b :
		TR_30 = RG_rl_201 ;
	7'h3c :
		TR_30 = RG_rl_201 ;
	7'h3d :
		TR_30 = RG_rl_201 ;
	7'h3e :
		TR_30 = RG_rl_201 ;
	7'h3f :
		TR_30 = RG_rl_201 ;
	7'h40 :
		TR_30 = RG_rl_201 ;
	7'h41 :
		TR_30 = RG_rl_201 ;
	7'h42 :
		TR_30 = RG_rl_201 ;
	7'h43 :
		TR_30 = RG_rl_201 ;
	7'h44 :
		TR_30 = RG_rl_201 ;
	7'h45 :
		TR_30 = RG_rl_201 ;
	7'h46 :
		TR_30 = RG_rl_201 ;
	7'h47 :
		TR_30 = RG_rl_201 ;
	7'h48 :
		TR_30 = RG_rl_201 ;
	7'h49 :
		TR_30 = RG_rl_201 ;
	7'h4a :
		TR_30 = RG_rl_201 ;
	7'h4b :
		TR_30 = RG_rl_201 ;
	7'h4c :
		TR_30 = RG_rl_201 ;
	7'h4d :
		TR_30 = RG_rl_201 ;
	7'h4e :
		TR_30 = RG_rl_201 ;
	7'h4f :
		TR_30 = RG_rl_201 ;
	7'h50 :
		TR_30 = RG_rl_201 ;
	7'h51 :
		TR_30 = RG_rl_201 ;
	7'h52 :
		TR_30 = RG_rl_201 ;
	7'h53 :
		TR_30 = RG_rl_201 ;
	7'h54 :
		TR_30 = RG_rl_201 ;
	7'h55 :
		TR_30 = RG_rl_201 ;
	7'h56 :
		TR_30 = RG_rl_201 ;
	7'h57 :
		TR_30 = RG_rl_201 ;
	7'h58 :
		TR_30 = RG_rl_201 ;
	7'h59 :
		TR_30 = RG_rl_201 ;
	7'h5a :
		TR_30 = RG_rl_201 ;
	7'h5b :
		TR_30 = RG_rl_201 ;
	7'h5c :
		TR_30 = RG_rl_201 ;
	7'h5d :
		TR_30 = RG_rl_201 ;
	7'h5e :
		TR_30 = RG_rl_201 ;
	7'h5f :
		TR_30 = RG_rl_201 ;
	7'h60 :
		TR_30 = RG_rl_201 ;
	7'h61 :
		TR_30 = RG_rl_201 ;
	7'h62 :
		TR_30 = RG_rl_201 ;
	7'h63 :
		TR_30 = RG_rl_201 ;
	7'h64 :
		TR_30 = RG_rl_201 ;
	7'h65 :
		TR_30 = RG_rl_201 ;
	7'h66 :
		TR_30 = RG_rl_201 ;
	7'h67 :
		TR_30 = RG_rl_201 ;
	7'h68 :
		TR_30 = RG_rl_201 ;
	7'h69 :
		TR_30 = RG_rl_201 ;
	7'h6a :
		TR_30 = RG_rl_201 ;
	7'h6b :
		TR_30 = RG_rl_201 ;
	7'h6c :
		TR_30 = RG_rl_201 ;
	7'h6d :
		TR_30 = RG_rl_201 ;
	7'h6e :
		TR_30 = RG_rl_201 ;
	7'h6f :
		TR_30 = RG_rl_201 ;
	7'h70 :
		TR_30 = RG_rl_201 ;
	7'h71 :
		TR_30 = RG_rl_201 ;
	7'h72 :
		TR_30 = RG_rl_201 ;
	7'h73 :
		TR_30 = RG_rl_201 ;
	7'h74 :
		TR_30 = RG_rl_201 ;
	7'h75 :
		TR_30 = RG_rl_201 ;
	7'h76 :
		TR_30 = RG_rl_201 ;
	7'h77 :
		TR_30 = RG_rl_201 ;
	7'h78 :
		TR_30 = RG_rl_201 ;
	7'h79 :
		TR_30 = RG_rl_201 ;
	7'h7a :
		TR_30 = RG_rl_201 ;
	7'h7b :
		TR_30 = RG_rl_201 ;
	7'h7c :
		TR_30 = RG_rl_201 ;
	7'h7d :
		TR_30 = RG_rl_201 ;
	7'h7e :
		TR_30 = RG_rl_201 ;
	7'h7f :
		TR_30 = RG_rl_201 ;
	default :
		TR_30 = 9'hx ;
	endcase
always @ ( RG_rl_202 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_31 = RG_rl_202 ;
	7'h01 :
		TR_31 = RG_rl_202 ;
	7'h02 :
		TR_31 = RG_rl_202 ;
	7'h03 :
		TR_31 = RG_rl_202 ;
	7'h04 :
		TR_31 = RG_rl_202 ;
	7'h05 :
		TR_31 = RG_rl_202 ;
	7'h06 :
		TR_31 = RG_rl_202 ;
	7'h07 :
		TR_31 = RG_rl_202 ;
	7'h08 :
		TR_31 = RG_rl_202 ;
	7'h09 :
		TR_31 = RG_rl_202 ;
	7'h0a :
		TR_31 = RG_rl_202 ;
	7'h0b :
		TR_31 = RG_rl_202 ;
	7'h0c :
		TR_31 = RG_rl_202 ;
	7'h0d :
		TR_31 = RG_rl_202 ;
	7'h0e :
		TR_31 = RG_rl_202 ;
	7'h0f :
		TR_31 = RG_rl_202 ;
	7'h10 :
		TR_31 = RG_rl_202 ;
	7'h11 :
		TR_31 = RG_rl_202 ;
	7'h12 :
		TR_31 = RG_rl_202 ;
	7'h13 :
		TR_31 = 9'h000 ;	// line#=../rle.cpp:68
	7'h14 :
		TR_31 = RG_rl_202 ;
	7'h15 :
		TR_31 = RG_rl_202 ;
	7'h16 :
		TR_31 = RG_rl_202 ;
	7'h17 :
		TR_31 = RG_rl_202 ;
	7'h18 :
		TR_31 = RG_rl_202 ;
	7'h19 :
		TR_31 = RG_rl_202 ;
	7'h1a :
		TR_31 = RG_rl_202 ;
	7'h1b :
		TR_31 = RG_rl_202 ;
	7'h1c :
		TR_31 = RG_rl_202 ;
	7'h1d :
		TR_31 = RG_rl_202 ;
	7'h1e :
		TR_31 = RG_rl_202 ;
	7'h1f :
		TR_31 = RG_rl_202 ;
	7'h20 :
		TR_31 = RG_rl_202 ;
	7'h21 :
		TR_31 = RG_rl_202 ;
	7'h22 :
		TR_31 = RG_rl_202 ;
	7'h23 :
		TR_31 = RG_rl_202 ;
	7'h24 :
		TR_31 = RG_rl_202 ;
	7'h25 :
		TR_31 = RG_rl_202 ;
	7'h26 :
		TR_31 = RG_rl_202 ;
	7'h27 :
		TR_31 = RG_rl_202 ;
	7'h28 :
		TR_31 = RG_rl_202 ;
	7'h29 :
		TR_31 = RG_rl_202 ;
	7'h2a :
		TR_31 = RG_rl_202 ;
	7'h2b :
		TR_31 = RG_rl_202 ;
	7'h2c :
		TR_31 = RG_rl_202 ;
	7'h2d :
		TR_31 = RG_rl_202 ;
	7'h2e :
		TR_31 = RG_rl_202 ;
	7'h2f :
		TR_31 = RG_rl_202 ;
	7'h30 :
		TR_31 = RG_rl_202 ;
	7'h31 :
		TR_31 = RG_rl_202 ;
	7'h32 :
		TR_31 = RG_rl_202 ;
	7'h33 :
		TR_31 = RG_rl_202 ;
	7'h34 :
		TR_31 = RG_rl_202 ;
	7'h35 :
		TR_31 = RG_rl_202 ;
	7'h36 :
		TR_31 = RG_rl_202 ;
	7'h37 :
		TR_31 = RG_rl_202 ;
	7'h38 :
		TR_31 = RG_rl_202 ;
	7'h39 :
		TR_31 = RG_rl_202 ;
	7'h3a :
		TR_31 = RG_rl_202 ;
	7'h3b :
		TR_31 = RG_rl_202 ;
	7'h3c :
		TR_31 = RG_rl_202 ;
	7'h3d :
		TR_31 = RG_rl_202 ;
	7'h3e :
		TR_31 = RG_rl_202 ;
	7'h3f :
		TR_31 = RG_rl_202 ;
	7'h40 :
		TR_31 = RG_rl_202 ;
	7'h41 :
		TR_31 = RG_rl_202 ;
	7'h42 :
		TR_31 = RG_rl_202 ;
	7'h43 :
		TR_31 = RG_rl_202 ;
	7'h44 :
		TR_31 = RG_rl_202 ;
	7'h45 :
		TR_31 = RG_rl_202 ;
	7'h46 :
		TR_31 = RG_rl_202 ;
	7'h47 :
		TR_31 = RG_rl_202 ;
	7'h48 :
		TR_31 = RG_rl_202 ;
	7'h49 :
		TR_31 = RG_rl_202 ;
	7'h4a :
		TR_31 = RG_rl_202 ;
	7'h4b :
		TR_31 = RG_rl_202 ;
	7'h4c :
		TR_31 = RG_rl_202 ;
	7'h4d :
		TR_31 = RG_rl_202 ;
	7'h4e :
		TR_31 = RG_rl_202 ;
	7'h4f :
		TR_31 = RG_rl_202 ;
	7'h50 :
		TR_31 = RG_rl_202 ;
	7'h51 :
		TR_31 = RG_rl_202 ;
	7'h52 :
		TR_31 = RG_rl_202 ;
	7'h53 :
		TR_31 = RG_rl_202 ;
	7'h54 :
		TR_31 = RG_rl_202 ;
	7'h55 :
		TR_31 = RG_rl_202 ;
	7'h56 :
		TR_31 = RG_rl_202 ;
	7'h57 :
		TR_31 = RG_rl_202 ;
	7'h58 :
		TR_31 = RG_rl_202 ;
	7'h59 :
		TR_31 = RG_rl_202 ;
	7'h5a :
		TR_31 = RG_rl_202 ;
	7'h5b :
		TR_31 = RG_rl_202 ;
	7'h5c :
		TR_31 = RG_rl_202 ;
	7'h5d :
		TR_31 = RG_rl_202 ;
	7'h5e :
		TR_31 = RG_rl_202 ;
	7'h5f :
		TR_31 = RG_rl_202 ;
	7'h60 :
		TR_31 = RG_rl_202 ;
	7'h61 :
		TR_31 = RG_rl_202 ;
	7'h62 :
		TR_31 = RG_rl_202 ;
	7'h63 :
		TR_31 = RG_rl_202 ;
	7'h64 :
		TR_31 = RG_rl_202 ;
	7'h65 :
		TR_31 = RG_rl_202 ;
	7'h66 :
		TR_31 = RG_rl_202 ;
	7'h67 :
		TR_31 = RG_rl_202 ;
	7'h68 :
		TR_31 = RG_rl_202 ;
	7'h69 :
		TR_31 = RG_rl_202 ;
	7'h6a :
		TR_31 = RG_rl_202 ;
	7'h6b :
		TR_31 = RG_rl_202 ;
	7'h6c :
		TR_31 = RG_rl_202 ;
	7'h6d :
		TR_31 = RG_rl_202 ;
	7'h6e :
		TR_31 = RG_rl_202 ;
	7'h6f :
		TR_31 = RG_rl_202 ;
	7'h70 :
		TR_31 = RG_rl_202 ;
	7'h71 :
		TR_31 = RG_rl_202 ;
	7'h72 :
		TR_31 = RG_rl_202 ;
	7'h73 :
		TR_31 = RG_rl_202 ;
	7'h74 :
		TR_31 = RG_rl_202 ;
	7'h75 :
		TR_31 = RG_rl_202 ;
	7'h76 :
		TR_31 = RG_rl_202 ;
	7'h77 :
		TR_31 = RG_rl_202 ;
	7'h78 :
		TR_31 = RG_rl_202 ;
	7'h79 :
		TR_31 = RG_rl_202 ;
	7'h7a :
		TR_31 = RG_rl_202 ;
	7'h7b :
		TR_31 = RG_rl_202 ;
	7'h7c :
		TR_31 = RG_rl_202 ;
	7'h7d :
		TR_31 = RG_rl_202 ;
	7'h7e :
		TR_31 = RG_rl_202 ;
	7'h7f :
		TR_31 = RG_rl_202 ;
	default :
		TR_31 = 9'hx ;
	endcase
always @ ( RG_rl_203 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_32 = RG_rl_203 ;
	7'h01 :
		TR_32 = RG_rl_203 ;
	7'h02 :
		TR_32 = RG_rl_203 ;
	7'h03 :
		TR_32 = RG_rl_203 ;
	7'h04 :
		TR_32 = RG_rl_203 ;
	7'h05 :
		TR_32 = RG_rl_203 ;
	7'h06 :
		TR_32 = RG_rl_203 ;
	7'h07 :
		TR_32 = RG_rl_203 ;
	7'h08 :
		TR_32 = RG_rl_203 ;
	7'h09 :
		TR_32 = RG_rl_203 ;
	7'h0a :
		TR_32 = RG_rl_203 ;
	7'h0b :
		TR_32 = RG_rl_203 ;
	7'h0c :
		TR_32 = RG_rl_203 ;
	7'h0d :
		TR_32 = RG_rl_203 ;
	7'h0e :
		TR_32 = RG_rl_203 ;
	7'h0f :
		TR_32 = RG_rl_203 ;
	7'h10 :
		TR_32 = RG_rl_203 ;
	7'h11 :
		TR_32 = RG_rl_203 ;
	7'h12 :
		TR_32 = RG_rl_203 ;
	7'h13 :
		TR_32 = RG_rl_203 ;
	7'h14 :
		TR_32 = 9'h000 ;	// line#=../rle.cpp:68
	7'h15 :
		TR_32 = RG_rl_203 ;
	7'h16 :
		TR_32 = RG_rl_203 ;
	7'h17 :
		TR_32 = RG_rl_203 ;
	7'h18 :
		TR_32 = RG_rl_203 ;
	7'h19 :
		TR_32 = RG_rl_203 ;
	7'h1a :
		TR_32 = RG_rl_203 ;
	7'h1b :
		TR_32 = RG_rl_203 ;
	7'h1c :
		TR_32 = RG_rl_203 ;
	7'h1d :
		TR_32 = RG_rl_203 ;
	7'h1e :
		TR_32 = RG_rl_203 ;
	7'h1f :
		TR_32 = RG_rl_203 ;
	7'h20 :
		TR_32 = RG_rl_203 ;
	7'h21 :
		TR_32 = RG_rl_203 ;
	7'h22 :
		TR_32 = RG_rl_203 ;
	7'h23 :
		TR_32 = RG_rl_203 ;
	7'h24 :
		TR_32 = RG_rl_203 ;
	7'h25 :
		TR_32 = RG_rl_203 ;
	7'h26 :
		TR_32 = RG_rl_203 ;
	7'h27 :
		TR_32 = RG_rl_203 ;
	7'h28 :
		TR_32 = RG_rl_203 ;
	7'h29 :
		TR_32 = RG_rl_203 ;
	7'h2a :
		TR_32 = RG_rl_203 ;
	7'h2b :
		TR_32 = RG_rl_203 ;
	7'h2c :
		TR_32 = RG_rl_203 ;
	7'h2d :
		TR_32 = RG_rl_203 ;
	7'h2e :
		TR_32 = RG_rl_203 ;
	7'h2f :
		TR_32 = RG_rl_203 ;
	7'h30 :
		TR_32 = RG_rl_203 ;
	7'h31 :
		TR_32 = RG_rl_203 ;
	7'h32 :
		TR_32 = RG_rl_203 ;
	7'h33 :
		TR_32 = RG_rl_203 ;
	7'h34 :
		TR_32 = RG_rl_203 ;
	7'h35 :
		TR_32 = RG_rl_203 ;
	7'h36 :
		TR_32 = RG_rl_203 ;
	7'h37 :
		TR_32 = RG_rl_203 ;
	7'h38 :
		TR_32 = RG_rl_203 ;
	7'h39 :
		TR_32 = RG_rl_203 ;
	7'h3a :
		TR_32 = RG_rl_203 ;
	7'h3b :
		TR_32 = RG_rl_203 ;
	7'h3c :
		TR_32 = RG_rl_203 ;
	7'h3d :
		TR_32 = RG_rl_203 ;
	7'h3e :
		TR_32 = RG_rl_203 ;
	7'h3f :
		TR_32 = RG_rl_203 ;
	7'h40 :
		TR_32 = RG_rl_203 ;
	7'h41 :
		TR_32 = RG_rl_203 ;
	7'h42 :
		TR_32 = RG_rl_203 ;
	7'h43 :
		TR_32 = RG_rl_203 ;
	7'h44 :
		TR_32 = RG_rl_203 ;
	7'h45 :
		TR_32 = RG_rl_203 ;
	7'h46 :
		TR_32 = RG_rl_203 ;
	7'h47 :
		TR_32 = RG_rl_203 ;
	7'h48 :
		TR_32 = RG_rl_203 ;
	7'h49 :
		TR_32 = RG_rl_203 ;
	7'h4a :
		TR_32 = RG_rl_203 ;
	7'h4b :
		TR_32 = RG_rl_203 ;
	7'h4c :
		TR_32 = RG_rl_203 ;
	7'h4d :
		TR_32 = RG_rl_203 ;
	7'h4e :
		TR_32 = RG_rl_203 ;
	7'h4f :
		TR_32 = RG_rl_203 ;
	7'h50 :
		TR_32 = RG_rl_203 ;
	7'h51 :
		TR_32 = RG_rl_203 ;
	7'h52 :
		TR_32 = RG_rl_203 ;
	7'h53 :
		TR_32 = RG_rl_203 ;
	7'h54 :
		TR_32 = RG_rl_203 ;
	7'h55 :
		TR_32 = RG_rl_203 ;
	7'h56 :
		TR_32 = RG_rl_203 ;
	7'h57 :
		TR_32 = RG_rl_203 ;
	7'h58 :
		TR_32 = RG_rl_203 ;
	7'h59 :
		TR_32 = RG_rl_203 ;
	7'h5a :
		TR_32 = RG_rl_203 ;
	7'h5b :
		TR_32 = RG_rl_203 ;
	7'h5c :
		TR_32 = RG_rl_203 ;
	7'h5d :
		TR_32 = RG_rl_203 ;
	7'h5e :
		TR_32 = RG_rl_203 ;
	7'h5f :
		TR_32 = RG_rl_203 ;
	7'h60 :
		TR_32 = RG_rl_203 ;
	7'h61 :
		TR_32 = RG_rl_203 ;
	7'h62 :
		TR_32 = RG_rl_203 ;
	7'h63 :
		TR_32 = RG_rl_203 ;
	7'h64 :
		TR_32 = RG_rl_203 ;
	7'h65 :
		TR_32 = RG_rl_203 ;
	7'h66 :
		TR_32 = RG_rl_203 ;
	7'h67 :
		TR_32 = RG_rl_203 ;
	7'h68 :
		TR_32 = RG_rl_203 ;
	7'h69 :
		TR_32 = RG_rl_203 ;
	7'h6a :
		TR_32 = RG_rl_203 ;
	7'h6b :
		TR_32 = RG_rl_203 ;
	7'h6c :
		TR_32 = RG_rl_203 ;
	7'h6d :
		TR_32 = RG_rl_203 ;
	7'h6e :
		TR_32 = RG_rl_203 ;
	7'h6f :
		TR_32 = RG_rl_203 ;
	7'h70 :
		TR_32 = RG_rl_203 ;
	7'h71 :
		TR_32 = RG_rl_203 ;
	7'h72 :
		TR_32 = RG_rl_203 ;
	7'h73 :
		TR_32 = RG_rl_203 ;
	7'h74 :
		TR_32 = RG_rl_203 ;
	7'h75 :
		TR_32 = RG_rl_203 ;
	7'h76 :
		TR_32 = RG_rl_203 ;
	7'h77 :
		TR_32 = RG_rl_203 ;
	7'h78 :
		TR_32 = RG_rl_203 ;
	7'h79 :
		TR_32 = RG_rl_203 ;
	7'h7a :
		TR_32 = RG_rl_203 ;
	7'h7b :
		TR_32 = RG_rl_203 ;
	7'h7c :
		TR_32 = RG_rl_203 ;
	7'h7d :
		TR_32 = RG_rl_203 ;
	7'h7e :
		TR_32 = RG_rl_203 ;
	7'h7f :
		TR_32 = RG_rl_203 ;
	default :
		TR_32 = 9'hx ;
	endcase
always @ ( RG_rl_204 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_33 = RG_rl_204 ;
	7'h01 :
		TR_33 = RG_rl_204 ;
	7'h02 :
		TR_33 = RG_rl_204 ;
	7'h03 :
		TR_33 = RG_rl_204 ;
	7'h04 :
		TR_33 = RG_rl_204 ;
	7'h05 :
		TR_33 = RG_rl_204 ;
	7'h06 :
		TR_33 = RG_rl_204 ;
	7'h07 :
		TR_33 = RG_rl_204 ;
	7'h08 :
		TR_33 = RG_rl_204 ;
	7'h09 :
		TR_33 = RG_rl_204 ;
	7'h0a :
		TR_33 = RG_rl_204 ;
	7'h0b :
		TR_33 = RG_rl_204 ;
	7'h0c :
		TR_33 = RG_rl_204 ;
	7'h0d :
		TR_33 = RG_rl_204 ;
	7'h0e :
		TR_33 = RG_rl_204 ;
	7'h0f :
		TR_33 = RG_rl_204 ;
	7'h10 :
		TR_33 = RG_rl_204 ;
	7'h11 :
		TR_33 = RG_rl_204 ;
	7'h12 :
		TR_33 = RG_rl_204 ;
	7'h13 :
		TR_33 = RG_rl_204 ;
	7'h14 :
		TR_33 = RG_rl_204 ;
	7'h15 :
		TR_33 = 9'h000 ;	// line#=../rle.cpp:68
	7'h16 :
		TR_33 = RG_rl_204 ;
	7'h17 :
		TR_33 = RG_rl_204 ;
	7'h18 :
		TR_33 = RG_rl_204 ;
	7'h19 :
		TR_33 = RG_rl_204 ;
	7'h1a :
		TR_33 = RG_rl_204 ;
	7'h1b :
		TR_33 = RG_rl_204 ;
	7'h1c :
		TR_33 = RG_rl_204 ;
	7'h1d :
		TR_33 = RG_rl_204 ;
	7'h1e :
		TR_33 = RG_rl_204 ;
	7'h1f :
		TR_33 = RG_rl_204 ;
	7'h20 :
		TR_33 = RG_rl_204 ;
	7'h21 :
		TR_33 = RG_rl_204 ;
	7'h22 :
		TR_33 = RG_rl_204 ;
	7'h23 :
		TR_33 = RG_rl_204 ;
	7'h24 :
		TR_33 = RG_rl_204 ;
	7'h25 :
		TR_33 = RG_rl_204 ;
	7'h26 :
		TR_33 = RG_rl_204 ;
	7'h27 :
		TR_33 = RG_rl_204 ;
	7'h28 :
		TR_33 = RG_rl_204 ;
	7'h29 :
		TR_33 = RG_rl_204 ;
	7'h2a :
		TR_33 = RG_rl_204 ;
	7'h2b :
		TR_33 = RG_rl_204 ;
	7'h2c :
		TR_33 = RG_rl_204 ;
	7'h2d :
		TR_33 = RG_rl_204 ;
	7'h2e :
		TR_33 = RG_rl_204 ;
	7'h2f :
		TR_33 = RG_rl_204 ;
	7'h30 :
		TR_33 = RG_rl_204 ;
	7'h31 :
		TR_33 = RG_rl_204 ;
	7'h32 :
		TR_33 = RG_rl_204 ;
	7'h33 :
		TR_33 = RG_rl_204 ;
	7'h34 :
		TR_33 = RG_rl_204 ;
	7'h35 :
		TR_33 = RG_rl_204 ;
	7'h36 :
		TR_33 = RG_rl_204 ;
	7'h37 :
		TR_33 = RG_rl_204 ;
	7'h38 :
		TR_33 = RG_rl_204 ;
	7'h39 :
		TR_33 = RG_rl_204 ;
	7'h3a :
		TR_33 = RG_rl_204 ;
	7'h3b :
		TR_33 = RG_rl_204 ;
	7'h3c :
		TR_33 = RG_rl_204 ;
	7'h3d :
		TR_33 = RG_rl_204 ;
	7'h3e :
		TR_33 = RG_rl_204 ;
	7'h3f :
		TR_33 = RG_rl_204 ;
	7'h40 :
		TR_33 = RG_rl_204 ;
	7'h41 :
		TR_33 = RG_rl_204 ;
	7'h42 :
		TR_33 = RG_rl_204 ;
	7'h43 :
		TR_33 = RG_rl_204 ;
	7'h44 :
		TR_33 = RG_rl_204 ;
	7'h45 :
		TR_33 = RG_rl_204 ;
	7'h46 :
		TR_33 = RG_rl_204 ;
	7'h47 :
		TR_33 = RG_rl_204 ;
	7'h48 :
		TR_33 = RG_rl_204 ;
	7'h49 :
		TR_33 = RG_rl_204 ;
	7'h4a :
		TR_33 = RG_rl_204 ;
	7'h4b :
		TR_33 = RG_rl_204 ;
	7'h4c :
		TR_33 = RG_rl_204 ;
	7'h4d :
		TR_33 = RG_rl_204 ;
	7'h4e :
		TR_33 = RG_rl_204 ;
	7'h4f :
		TR_33 = RG_rl_204 ;
	7'h50 :
		TR_33 = RG_rl_204 ;
	7'h51 :
		TR_33 = RG_rl_204 ;
	7'h52 :
		TR_33 = RG_rl_204 ;
	7'h53 :
		TR_33 = RG_rl_204 ;
	7'h54 :
		TR_33 = RG_rl_204 ;
	7'h55 :
		TR_33 = RG_rl_204 ;
	7'h56 :
		TR_33 = RG_rl_204 ;
	7'h57 :
		TR_33 = RG_rl_204 ;
	7'h58 :
		TR_33 = RG_rl_204 ;
	7'h59 :
		TR_33 = RG_rl_204 ;
	7'h5a :
		TR_33 = RG_rl_204 ;
	7'h5b :
		TR_33 = RG_rl_204 ;
	7'h5c :
		TR_33 = RG_rl_204 ;
	7'h5d :
		TR_33 = RG_rl_204 ;
	7'h5e :
		TR_33 = RG_rl_204 ;
	7'h5f :
		TR_33 = RG_rl_204 ;
	7'h60 :
		TR_33 = RG_rl_204 ;
	7'h61 :
		TR_33 = RG_rl_204 ;
	7'h62 :
		TR_33 = RG_rl_204 ;
	7'h63 :
		TR_33 = RG_rl_204 ;
	7'h64 :
		TR_33 = RG_rl_204 ;
	7'h65 :
		TR_33 = RG_rl_204 ;
	7'h66 :
		TR_33 = RG_rl_204 ;
	7'h67 :
		TR_33 = RG_rl_204 ;
	7'h68 :
		TR_33 = RG_rl_204 ;
	7'h69 :
		TR_33 = RG_rl_204 ;
	7'h6a :
		TR_33 = RG_rl_204 ;
	7'h6b :
		TR_33 = RG_rl_204 ;
	7'h6c :
		TR_33 = RG_rl_204 ;
	7'h6d :
		TR_33 = RG_rl_204 ;
	7'h6e :
		TR_33 = RG_rl_204 ;
	7'h6f :
		TR_33 = RG_rl_204 ;
	7'h70 :
		TR_33 = RG_rl_204 ;
	7'h71 :
		TR_33 = RG_rl_204 ;
	7'h72 :
		TR_33 = RG_rl_204 ;
	7'h73 :
		TR_33 = RG_rl_204 ;
	7'h74 :
		TR_33 = RG_rl_204 ;
	7'h75 :
		TR_33 = RG_rl_204 ;
	7'h76 :
		TR_33 = RG_rl_204 ;
	7'h77 :
		TR_33 = RG_rl_204 ;
	7'h78 :
		TR_33 = RG_rl_204 ;
	7'h79 :
		TR_33 = RG_rl_204 ;
	7'h7a :
		TR_33 = RG_rl_204 ;
	7'h7b :
		TR_33 = RG_rl_204 ;
	7'h7c :
		TR_33 = RG_rl_204 ;
	7'h7d :
		TR_33 = RG_rl_204 ;
	7'h7e :
		TR_33 = RG_rl_204 ;
	7'h7f :
		TR_33 = RG_rl_204 ;
	default :
		TR_33 = 9'hx ;
	endcase
always @ ( RG_rl_205 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_34 = RG_rl_205 ;
	7'h01 :
		TR_34 = RG_rl_205 ;
	7'h02 :
		TR_34 = RG_rl_205 ;
	7'h03 :
		TR_34 = RG_rl_205 ;
	7'h04 :
		TR_34 = RG_rl_205 ;
	7'h05 :
		TR_34 = RG_rl_205 ;
	7'h06 :
		TR_34 = RG_rl_205 ;
	7'h07 :
		TR_34 = RG_rl_205 ;
	7'h08 :
		TR_34 = RG_rl_205 ;
	7'h09 :
		TR_34 = RG_rl_205 ;
	7'h0a :
		TR_34 = RG_rl_205 ;
	7'h0b :
		TR_34 = RG_rl_205 ;
	7'h0c :
		TR_34 = RG_rl_205 ;
	7'h0d :
		TR_34 = RG_rl_205 ;
	7'h0e :
		TR_34 = RG_rl_205 ;
	7'h0f :
		TR_34 = RG_rl_205 ;
	7'h10 :
		TR_34 = RG_rl_205 ;
	7'h11 :
		TR_34 = RG_rl_205 ;
	7'h12 :
		TR_34 = RG_rl_205 ;
	7'h13 :
		TR_34 = RG_rl_205 ;
	7'h14 :
		TR_34 = RG_rl_205 ;
	7'h15 :
		TR_34 = RG_rl_205 ;
	7'h16 :
		TR_34 = 9'h000 ;	// line#=../rle.cpp:68
	7'h17 :
		TR_34 = RG_rl_205 ;
	7'h18 :
		TR_34 = RG_rl_205 ;
	7'h19 :
		TR_34 = RG_rl_205 ;
	7'h1a :
		TR_34 = RG_rl_205 ;
	7'h1b :
		TR_34 = RG_rl_205 ;
	7'h1c :
		TR_34 = RG_rl_205 ;
	7'h1d :
		TR_34 = RG_rl_205 ;
	7'h1e :
		TR_34 = RG_rl_205 ;
	7'h1f :
		TR_34 = RG_rl_205 ;
	7'h20 :
		TR_34 = RG_rl_205 ;
	7'h21 :
		TR_34 = RG_rl_205 ;
	7'h22 :
		TR_34 = RG_rl_205 ;
	7'h23 :
		TR_34 = RG_rl_205 ;
	7'h24 :
		TR_34 = RG_rl_205 ;
	7'h25 :
		TR_34 = RG_rl_205 ;
	7'h26 :
		TR_34 = RG_rl_205 ;
	7'h27 :
		TR_34 = RG_rl_205 ;
	7'h28 :
		TR_34 = RG_rl_205 ;
	7'h29 :
		TR_34 = RG_rl_205 ;
	7'h2a :
		TR_34 = RG_rl_205 ;
	7'h2b :
		TR_34 = RG_rl_205 ;
	7'h2c :
		TR_34 = RG_rl_205 ;
	7'h2d :
		TR_34 = RG_rl_205 ;
	7'h2e :
		TR_34 = RG_rl_205 ;
	7'h2f :
		TR_34 = RG_rl_205 ;
	7'h30 :
		TR_34 = RG_rl_205 ;
	7'h31 :
		TR_34 = RG_rl_205 ;
	7'h32 :
		TR_34 = RG_rl_205 ;
	7'h33 :
		TR_34 = RG_rl_205 ;
	7'h34 :
		TR_34 = RG_rl_205 ;
	7'h35 :
		TR_34 = RG_rl_205 ;
	7'h36 :
		TR_34 = RG_rl_205 ;
	7'h37 :
		TR_34 = RG_rl_205 ;
	7'h38 :
		TR_34 = RG_rl_205 ;
	7'h39 :
		TR_34 = RG_rl_205 ;
	7'h3a :
		TR_34 = RG_rl_205 ;
	7'h3b :
		TR_34 = RG_rl_205 ;
	7'h3c :
		TR_34 = RG_rl_205 ;
	7'h3d :
		TR_34 = RG_rl_205 ;
	7'h3e :
		TR_34 = RG_rl_205 ;
	7'h3f :
		TR_34 = RG_rl_205 ;
	7'h40 :
		TR_34 = RG_rl_205 ;
	7'h41 :
		TR_34 = RG_rl_205 ;
	7'h42 :
		TR_34 = RG_rl_205 ;
	7'h43 :
		TR_34 = RG_rl_205 ;
	7'h44 :
		TR_34 = RG_rl_205 ;
	7'h45 :
		TR_34 = RG_rl_205 ;
	7'h46 :
		TR_34 = RG_rl_205 ;
	7'h47 :
		TR_34 = RG_rl_205 ;
	7'h48 :
		TR_34 = RG_rl_205 ;
	7'h49 :
		TR_34 = RG_rl_205 ;
	7'h4a :
		TR_34 = RG_rl_205 ;
	7'h4b :
		TR_34 = RG_rl_205 ;
	7'h4c :
		TR_34 = RG_rl_205 ;
	7'h4d :
		TR_34 = RG_rl_205 ;
	7'h4e :
		TR_34 = RG_rl_205 ;
	7'h4f :
		TR_34 = RG_rl_205 ;
	7'h50 :
		TR_34 = RG_rl_205 ;
	7'h51 :
		TR_34 = RG_rl_205 ;
	7'h52 :
		TR_34 = RG_rl_205 ;
	7'h53 :
		TR_34 = RG_rl_205 ;
	7'h54 :
		TR_34 = RG_rl_205 ;
	7'h55 :
		TR_34 = RG_rl_205 ;
	7'h56 :
		TR_34 = RG_rl_205 ;
	7'h57 :
		TR_34 = RG_rl_205 ;
	7'h58 :
		TR_34 = RG_rl_205 ;
	7'h59 :
		TR_34 = RG_rl_205 ;
	7'h5a :
		TR_34 = RG_rl_205 ;
	7'h5b :
		TR_34 = RG_rl_205 ;
	7'h5c :
		TR_34 = RG_rl_205 ;
	7'h5d :
		TR_34 = RG_rl_205 ;
	7'h5e :
		TR_34 = RG_rl_205 ;
	7'h5f :
		TR_34 = RG_rl_205 ;
	7'h60 :
		TR_34 = RG_rl_205 ;
	7'h61 :
		TR_34 = RG_rl_205 ;
	7'h62 :
		TR_34 = RG_rl_205 ;
	7'h63 :
		TR_34 = RG_rl_205 ;
	7'h64 :
		TR_34 = RG_rl_205 ;
	7'h65 :
		TR_34 = RG_rl_205 ;
	7'h66 :
		TR_34 = RG_rl_205 ;
	7'h67 :
		TR_34 = RG_rl_205 ;
	7'h68 :
		TR_34 = RG_rl_205 ;
	7'h69 :
		TR_34 = RG_rl_205 ;
	7'h6a :
		TR_34 = RG_rl_205 ;
	7'h6b :
		TR_34 = RG_rl_205 ;
	7'h6c :
		TR_34 = RG_rl_205 ;
	7'h6d :
		TR_34 = RG_rl_205 ;
	7'h6e :
		TR_34 = RG_rl_205 ;
	7'h6f :
		TR_34 = RG_rl_205 ;
	7'h70 :
		TR_34 = RG_rl_205 ;
	7'h71 :
		TR_34 = RG_rl_205 ;
	7'h72 :
		TR_34 = RG_rl_205 ;
	7'h73 :
		TR_34 = RG_rl_205 ;
	7'h74 :
		TR_34 = RG_rl_205 ;
	7'h75 :
		TR_34 = RG_rl_205 ;
	7'h76 :
		TR_34 = RG_rl_205 ;
	7'h77 :
		TR_34 = RG_rl_205 ;
	7'h78 :
		TR_34 = RG_rl_205 ;
	7'h79 :
		TR_34 = RG_rl_205 ;
	7'h7a :
		TR_34 = RG_rl_205 ;
	7'h7b :
		TR_34 = RG_rl_205 ;
	7'h7c :
		TR_34 = RG_rl_205 ;
	7'h7d :
		TR_34 = RG_rl_205 ;
	7'h7e :
		TR_34 = RG_rl_205 ;
	7'h7f :
		TR_34 = RG_rl_205 ;
	default :
		TR_34 = 9'hx ;
	endcase
always @ ( RG_rl_206 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_35 = RG_rl_206 ;
	7'h01 :
		TR_35 = RG_rl_206 ;
	7'h02 :
		TR_35 = RG_rl_206 ;
	7'h03 :
		TR_35 = RG_rl_206 ;
	7'h04 :
		TR_35 = RG_rl_206 ;
	7'h05 :
		TR_35 = RG_rl_206 ;
	7'h06 :
		TR_35 = RG_rl_206 ;
	7'h07 :
		TR_35 = RG_rl_206 ;
	7'h08 :
		TR_35 = RG_rl_206 ;
	7'h09 :
		TR_35 = RG_rl_206 ;
	7'h0a :
		TR_35 = RG_rl_206 ;
	7'h0b :
		TR_35 = RG_rl_206 ;
	7'h0c :
		TR_35 = RG_rl_206 ;
	7'h0d :
		TR_35 = RG_rl_206 ;
	7'h0e :
		TR_35 = RG_rl_206 ;
	7'h0f :
		TR_35 = RG_rl_206 ;
	7'h10 :
		TR_35 = RG_rl_206 ;
	7'h11 :
		TR_35 = RG_rl_206 ;
	7'h12 :
		TR_35 = RG_rl_206 ;
	7'h13 :
		TR_35 = RG_rl_206 ;
	7'h14 :
		TR_35 = RG_rl_206 ;
	7'h15 :
		TR_35 = RG_rl_206 ;
	7'h16 :
		TR_35 = RG_rl_206 ;
	7'h17 :
		TR_35 = 9'h000 ;	// line#=../rle.cpp:68
	7'h18 :
		TR_35 = RG_rl_206 ;
	7'h19 :
		TR_35 = RG_rl_206 ;
	7'h1a :
		TR_35 = RG_rl_206 ;
	7'h1b :
		TR_35 = RG_rl_206 ;
	7'h1c :
		TR_35 = RG_rl_206 ;
	7'h1d :
		TR_35 = RG_rl_206 ;
	7'h1e :
		TR_35 = RG_rl_206 ;
	7'h1f :
		TR_35 = RG_rl_206 ;
	7'h20 :
		TR_35 = RG_rl_206 ;
	7'h21 :
		TR_35 = RG_rl_206 ;
	7'h22 :
		TR_35 = RG_rl_206 ;
	7'h23 :
		TR_35 = RG_rl_206 ;
	7'h24 :
		TR_35 = RG_rl_206 ;
	7'h25 :
		TR_35 = RG_rl_206 ;
	7'h26 :
		TR_35 = RG_rl_206 ;
	7'h27 :
		TR_35 = RG_rl_206 ;
	7'h28 :
		TR_35 = RG_rl_206 ;
	7'h29 :
		TR_35 = RG_rl_206 ;
	7'h2a :
		TR_35 = RG_rl_206 ;
	7'h2b :
		TR_35 = RG_rl_206 ;
	7'h2c :
		TR_35 = RG_rl_206 ;
	7'h2d :
		TR_35 = RG_rl_206 ;
	7'h2e :
		TR_35 = RG_rl_206 ;
	7'h2f :
		TR_35 = RG_rl_206 ;
	7'h30 :
		TR_35 = RG_rl_206 ;
	7'h31 :
		TR_35 = RG_rl_206 ;
	7'h32 :
		TR_35 = RG_rl_206 ;
	7'h33 :
		TR_35 = RG_rl_206 ;
	7'h34 :
		TR_35 = RG_rl_206 ;
	7'h35 :
		TR_35 = RG_rl_206 ;
	7'h36 :
		TR_35 = RG_rl_206 ;
	7'h37 :
		TR_35 = RG_rl_206 ;
	7'h38 :
		TR_35 = RG_rl_206 ;
	7'h39 :
		TR_35 = RG_rl_206 ;
	7'h3a :
		TR_35 = RG_rl_206 ;
	7'h3b :
		TR_35 = RG_rl_206 ;
	7'h3c :
		TR_35 = RG_rl_206 ;
	7'h3d :
		TR_35 = RG_rl_206 ;
	7'h3e :
		TR_35 = RG_rl_206 ;
	7'h3f :
		TR_35 = RG_rl_206 ;
	7'h40 :
		TR_35 = RG_rl_206 ;
	7'h41 :
		TR_35 = RG_rl_206 ;
	7'h42 :
		TR_35 = RG_rl_206 ;
	7'h43 :
		TR_35 = RG_rl_206 ;
	7'h44 :
		TR_35 = RG_rl_206 ;
	7'h45 :
		TR_35 = RG_rl_206 ;
	7'h46 :
		TR_35 = RG_rl_206 ;
	7'h47 :
		TR_35 = RG_rl_206 ;
	7'h48 :
		TR_35 = RG_rl_206 ;
	7'h49 :
		TR_35 = RG_rl_206 ;
	7'h4a :
		TR_35 = RG_rl_206 ;
	7'h4b :
		TR_35 = RG_rl_206 ;
	7'h4c :
		TR_35 = RG_rl_206 ;
	7'h4d :
		TR_35 = RG_rl_206 ;
	7'h4e :
		TR_35 = RG_rl_206 ;
	7'h4f :
		TR_35 = RG_rl_206 ;
	7'h50 :
		TR_35 = RG_rl_206 ;
	7'h51 :
		TR_35 = RG_rl_206 ;
	7'h52 :
		TR_35 = RG_rl_206 ;
	7'h53 :
		TR_35 = RG_rl_206 ;
	7'h54 :
		TR_35 = RG_rl_206 ;
	7'h55 :
		TR_35 = RG_rl_206 ;
	7'h56 :
		TR_35 = RG_rl_206 ;
	7'h57 :
		TR_35 = RG_rl_206 ;
	7'h58 :
		TR_35 = RG_rl_206 ;
	7'h59 :
		TR_35 = RG_rl_206 ;
	7'h5a :
		TR_35 = RG_rl_206 ;
	7'h5b :
		TR_35 = RG_rl_206 ;
	7'h5c :
		TR_35 = RG_rl_206 ;
	7'h5d :
		TR_35 = RG_rl_206 ;
	7'h5e :
		TR_35 = RG_rl_206 ;
	7'h5f :
		TR_35 = RG_rl_206 ;
	7'h60 :
		TR_35 = RG_rl_206 ;
	7'h61 :
		TR_35 = RG_rl_206 ;
	7'h62 :
		TR_35 = RG_rl_206 ;
	7'h63 :
		TR_35 = RG_rl_206 ;
	7'h64 :
		TR_35 = RG_rl_206 ;
	7'h65 :
		TR_35 = RG_rl_206 ;
	7'h66 :
		TR_35 = RG_rl_206 ;
	7'h67 :
		TR_35 = RG_rl_206 ;
	7'h68 :
		TR_35 = RG_rl_206 ;
	7'h69 :
		TR_35 = RG_rl_206 ;
	7'h6a :
		TR_35 = RG_rl_206 ;
	7'h6b :
		TR_35 = RG_rl_206 ;
	7'h6c :
		TR_35 = RG_rl_206 ;
	7'h6d :
		TR_35 = RG_rl_206 ;
	7'h6e :
		TR_35 = RG_rl_206 ;
	7'h6f :
		TR_35 = RG_rl_206 ;
	7'h70 :
		TR_35 = RG_rl_206 ;
	7'h71 :
		TR_35 = RG_rl_206 ;
	7'h72 :
		TR_35 = RG_rl_206 ;
	7'h73 :
		TR_35 = RG_rl_206 ;
	7'h74 :
		TR_35 = RG_rl_206 ;
	7'h75 :
		TR_35 = RG_rl_206 ;
	7'h76 :
		TR_35 = RG_rl_206 ;
	7'h77 :
		TR_35 = RG_rl_206 ;
	7'h78 :
		TR_35 = RG_rl_206 ;
	7'h79 :
		TR_35 = RG_rl_206 ;
	7'h7a :
		TR_35 = RG_rl_206 ;
	7'h7b :
		TR_35 = RG_rl_206 ;
	7'h7c :
		TR_35 = RG_rl_206 ;
	7'h7d :
		TR_35 = RG_rl_206 ;
	7'h7e :
		TR_35 = RG_rl_206 ;
	7'h7f :
		TR_35 = RG_rl_206 ;
	default :
		TR_35 = 9'hx ;
	endcase
always @ ( RG_rl_207 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_36 = RG_rl_207 ;
	7'h01 :
		TR_36 = RG_rl_207 ;
	7'h02 :
		TR_36 = RG_rl_207 ;
	7'h03 :
		TR_36 = RG_rl_207 ;
	7'h04 :
		TR_36 = RG_rl_207 ;
	7'h05 :
		TR_36 = RG_rl_207 ;
	7'h06 :
		TR_36 = RG_rl_207 ;
	7'h07 :
		TR_36 = RG_rl_207 ;
	7'h08 :
		TR_36 = RG_rl_207 ;
	7'h09 :
		TR_36 = RG_rl_207 ;
	7'h0a :
		TR_36 = RG_rl_207 ;
	7'h0b :
		TR_36 = RG_rl_207 ;
	7'h0c :
		TR_36 = RG_rl_207 ;
	7'h0d :
		TR_36 = RG_rl_207 ;
	7'h0e :
		TR_36 = RG_rl_207 ;
	7'h0f :
		TR_36 = RG_rl_207 ;
	7'h10 :
		TR_36 = RG_rl_207 ;
	7'h11 :
		TR_36 = RG_rl_207 ;
	7'h12 :
		TR_36 = RG_rl_207 ;
	7'h13 :
		TR_36 = RG_rl_207 ;
	7'h14 :
		TR_36 = RG_rl_207 ;
	7'h15 :
		TR_36 = RG_rl_207 ;
	7'h16 :
		TR_36 = RG_rl_207 ;
	7'h17 :
		TR_36 = RG_rl_207 ;
	7'h18 :
		TR_36 = 9'h000 ;	// line#=../rle.cpp:68
	7'h19 :
		TR_36 = RG_rl_207 ;
	7'h1a :
		TR_36 = RG_rl_207 ;
	7'h1b :
		TR_36 = RG_rl_207 ;
	7'h1c :
		TR_36 = RG_rl_207 ;
	7'h1d :
		TR_36 = RG_rl_207 ;
	7'h1e :
		TR_36 = RG_rl_207 ;
	7'h1f :
		TR_36 = RG_rl_207 ;
	7'h20 :
		TR_36 = RG_rl_207 ;
	7'h21 :
		TR_36 = RG_rl_207 ;
	7'h22 :
		TR_36 = RG_rl_207 ;
	7'h23 :
		TR_36 = RG_rl_207 ;
	7'h24 :
		TR_36 = RG_rl_207 ;
	7'h25 :
		TR_36 = RG_rl_207 ;
	7'h26 :
		TR_36 = RG_rl_207 ;
	7'h27 :
		TR_36 = RG_rl_207 ;
	7'h28 :
		TR_36 = RG_rl_207 ;
	7'h29 :
		TR_36 = RG_rl_207 ;
	7'h2a :
		TR_36 = RG_rl_207 ;
	7'h2b :
		TR_36 = RG_rl_207 ;
	7'h2c :
		TR_36 = RG_rl_207 ;
	7'h2d :
		TR_36 = RG_rl_207 ;
	7'h2e :
		TR_36 = RG_rl_207 ;
	7'h2f :
		TR_36 = RG_rl_207 ;
	7'h30 :
		TR_36 = RG_rl_207 ;
	7'h31 :
		TR_36 = RG_rl_207 ;
	7'h32 :
		TR_36 = RG_rl_207 ;
	7'h33 :
		TR_36 = RG_rl_207 ;
	7'h34 :
		TR_36 = RG_rl_207 ;
	7'h35 :
		TR_36 = RG_rl_207 ;
	7'h36 :
		TR_36 = RG_rl_207 ;
	7'h37 :
		TR_36 = RG_rl_207 ;
	7'h38 :
		TR_36 = RG_rl_207 ;
	7'h39 :
		TR_36 = RG_rl_207 ;
	7'h3a :
		TR_36 = RG_rl_207 ;
	7'h3b :
		TR_36 = RG_rl_207 ;
	7'h3c :
		TR_36 = RG_rl_207 ;
	7'h3d :
		TR_36 = RG_rl_207 ;
	7'h3e :
		TR_36 = RG_rl_207 ;
	7'h3f :
		TR_36 = RG_rl_207 ;
	7'h40 :
		TR_36 = RG_rl_207 ;
	7'h41 :
		TR_36 = RG_rl_207 ;
	7'h42 :
		TR_36 = RG_rl_207 ;
	7'h43 :
		TR_36 = RG_rl_207 ;
	7'h44 :
		TR_36 = RG_rl_207 ;
	7'h45 :
		TR_36 = RG_rl_207 ;
	7'h46 :
		TR_36 = RG_rl_207 ;
	7'h47 :
		TR_36 = RG_rl_207 ;
	7'h48 :
		TR_36 = RG_rl_207 ;
	7'h49 :
		TR_36 = RG_rl_207 ;
	7'h4a :
		TR_36 = RG_rl_207 ;
	7'h4b :
		TR_36 = RG_rl_207 ;
	7'h4c :
		TR_36 = RG_rl_207 ;
	7'h4d :
		TR_36 = RG_rl_207 ;
	7'h4e :
		TR_36 = RG_rl_207 ;
	7'h4f :
		TR_36 = RG_rl_207 ;
	7'h50 :
		TR_36 = RG_rl_207 ;
	7'h51 :
		TR_36 = RG_rl_207 ;
	7'h52 :
		TR_36 = RG_rl_207 ;
	7'h53 :
		TR_36 = RG_rl_207 ;
	7'h54 :
		TR_36 = RG_rl_207 ;
	7'h55 :
		TR_36 = RG_rl_207 ;
	7'h56 :
		TR_36 = RG_rl_207 ;
	7'h57 :
		TR_36 = RG_rl_207 ;
	7'h58 :
		TR_36 = RG_rl_207 ;
	7'h59 :
		TR_36 = RG_rl_207 ;
	7'h5a :
		TR_36 = RG_rl_207 ;
	7'h5b :
		TR_36 = RG_rl_207 ;
	7'h5c :
		TR_36 = RG_rl_207 ;
	7'h5d :
		TR_36 = RG_rl_207 ;
	7'h5e :
		TR_36 = RG_rl_207 ;
	7'h5f :
		TR_36 = RG_rl_207 ;
	7'h60 :
		TR_36 = RG_rl_207 ;
	7'h61 :
		TR_36 = RG_rl_207 ;
	7'h62 :
		TR_36 = RG_rl_207 ;
	7'h63 :
		TR_36 = RG_rl_207 ;
	7'h64 :
		TR_36 = RG_rl_207 ;
	7'h65 :
		TR_36 = RG_rl_207 ;
	7'h66 :
		TR_36 = RG_rl_207 ;
	7'h67 :
		TR_36 = RG_rl_207 ;
	7'h68 :
		TR_36 = RG_rl_207 ;
	7'h69 :
		TR_36 = RG_rl_207 ;
	7'h6a :
		TR_36 = RG_rl_207 ;
	7'h6b :
		TR_36 = RG_rl_207 ;
	7'h6c :
		TR_36 = RG_rl_207 ;
	7'h6d :
		TR_36 = RG_rl_207 ;
	7'h6e :
		TR_36 = RG_rl_207 ;
	7'h6f :
		TR_36 = RG_rl_207 ;
	7'h70 :
		TR_36 = RG_rl_207 ;
	7'h71 :
		TR_36 = RG_rl_207 ;
	7'h72 :
		TR_36 = RG_rl_207 ;
	7'h73 :
		TR_36 = RG_rl_207 ;
	7'h74 :
		TR_36 = RG_rl_207 ;
	7'h75 :
		TR_36 = RG_rl_207 ;
	7'h76 :
		TR_36 = RG_rl_207 ;
	7'h77 :
		TR_36 = RG_rl_207 ;
	7'h78 :
		TR_36 = RG_rl_207 ;
	7'h79 :
		TR_36 = RG_rl_207 ;
	7'h7a :
		TR_36 = RG_rl_207 ;
	7'h7b :
		TR_36 = RG_rl_207 ;
	7'h7c :
		TR_36 = RG_rl_207 ;
	7'h7d :
		TR_36 = RG_rl_207 ;
	7'h7e :
		TR_36 = RG_rl_207 ;
	7'h7f :
		TR_36 = RG_rl_207 ;
	default :
		TR_36 = 9'hx ;
	endcase
always @ ( RG_rl_208 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_37 = RG_rl_208 ;
	7'h01 :
		TR_37 = RG_rl_208 ;
	7'h02 :
		TR_37 = RG_rl_208 ;
	7'h03 :
		TR_37 = RG_rl_208 ;
	7'h04 :
		TR_37 = RG_rl_208 ;
	7'h05 :
		TR_37 = RG_rl_208 ;
	7'h06 :
		TR_37 = RG_rl_208 ;
	7'h07 :
		TR_37 = RG_rl_208 ;
	7'h08 :
		TR_37 = RG_rl_208 ;
	7'h09 :
		TR_37 = RG_rl_208 ;
	7'h0a :
		TR_37 = RG_rl_208 ;
	7'h0b :
		TR_37 = RG_rl_208 ;
	7'h0c :
		TR_37 = RG_rl_208 ;
	7'h0d :
		TR_37 = RG_rl_208 ;
	7'h0e :
		TR_37 = RG_rl_208 ;
	7'h0f :
		TR_37 = RG_rl_208 ;
	7'h10 :
		TR_37 = RG_rl_208 ;
	7'h11 :
		TR_37 = RG_rl_208 ;
	7'h12 :
		TR_37 = RG_rl_208 ;
	7'h13 :
		TR_37 = RG_rl_208 ;
	7'h14 :
		TR_37 = RG_rl_208 ;
	7'h15 :
		TR_37 = RG_rl_208 ;
	7'h16 :
		TR_37 = RG_rl_208 ;
	7'h17 :
		TR_37 = RG_rl_208 ;
	7'h18 :
		TR_37 = RG_rl_208 ;
	7'h19 :
		TR_37 = 9'h000 ;	// line#=../rle.cpp:68
	7'h1a :
		TR_37 = RG_rl_208 ;
	7'h1b :
		TR_37 = RG_rl_208 ;
	7'h1c :
		TR_37 = RG_rl_208 ;
	7'h1d :
		TR_37 = RG_rl_208 ;
	7'h1e :
		TR_37 = RG_rl_208 ;
	7'h1f :
		TR_37 = RG_rl_208 ;
	7'h20 :
		TR_37 = RG_rl_208 ;
	7'h21 :
		TR_37 = RG_rl_208 ;
	7'h22 :
		TR_37 = RG_rl_208 ;
	7'h23 :
		TR_37 = RG_rl_208 ;
	7'h24 :
		TR_37 = RG_rl_208 ;
	7'h25 :
		TR_37 = RG_rl_208 ;
	7'h26 :
		TR_37 = RG_rl_208 ;
	7'h27 :
		TR_37 = RG_rl_208 ;
	7'h28 :
		TR_37 = RG_rl_208 ;
	7'h29 :
		TR_37 = RG_rl_208 ;
	7'h2a :
		TR_37 = RG_rl_208 ;
	7'h2b :
		TR_37 = RG_rl_208 ;
	7'h2c :
		TR_37 = RG_rl_208 ;
	7'h2d :
		TR_37 = RG_rl_208 ;
	7'h2e :
		TR_37 = RG_rl_208 ;
	7'h2f :
		TR_37 = RG_rl_208 ;
	7'h30 :
		TR_37 = RG_rl_208 ;
	7'h31 :
		TR_37 = RG_rl_208 ;
	7'h32 :
		TR_37 = RG_rl_208 ;
	7'h33 :
		TR_37 = RG_rl_208 ;
	7'h34 :
		TR_37 = RG_rl_208 ;
	7'h35 :
		TR_37 = RG_rl_208 ;
	7'h36 :
		TR_37 = RG_rl_208 ;
	7'h37 :
		TR_37 = RG_rl_208 ;
	7'h38 :
		TR_37 = RG_rl_208 ;
	7'h39 :
		TR_37 = RG_rl_208 ;
	7'h3a :
		TR_37 = RG_rl_208 ;
	7'h3b :
		TR_37 = RG_rl_208 ;
	7'h3c :
		TR_37 = RG_rl_208 ;
	7'h3d :
		TR_37 = RG_rl_208 ;
	7'h3e :
		TR_37 = RG_rl_208 ;
	7'h3f :
		TR_37 = RG_rl_208 ;
	7'h40 :
		TR_37 = RG_rl_208 ;
	7'h41 :
		TR_37 = RG_rl_208 ;
	7'h42 :
		TR_37 = RG_rl_208 ;
	7'h43 :
		TR_37 = RG_rl_208 ;
	7'h44 :
		TR_37 = RG_rl_208 ;
	7'h45 :
		TR_37 = RG_rl_208 ;
	7'h46 :
		TR_37 = RG_rl_208 ;
	7'h47 :
		TR_37 = RG_rl_208 ;
	7'h48 :
		TR_37 = RG_rl_208 ;
	7'h49 :
		TR_37 = RG_rl_208 ;
	7'h4a :
		TR_37 = RG_rl_208 ;
	7'h4b :
		TR_37 = RG_rl_208 ;
	7'h4c :
		TR_37 = RG_rl_208 ;
	7'h4d :
		TR_37 = RG_rl_208 ;
	7'h4e :
		TR_37 = RG_rl_208 ;
	7'h4f :
		TR_37 = RG_rl_208 ;
	7'h50 :
		TR_37 = RG_rl_208 ;
	7'h51 :
		TR_37 = RG_rl_208 ;
	7'h52 :
		TR_37 = RG_rl_208 ;
	7'h53 :
		TR_37 = RG_rl_208 ;
	7'h54 :
		TR_37 = RG_rl_208 ;
	7'h55 :
		TR_37 = RG_rl_208 ;
	7'h56 :
		TR_37 = RG_rl_208 ;
	7'h57 :
		TR_37 = RG_rl_208 ;
	7'h58 :
		TR_37 = RG_rl_208 ;
	7'h59 :
		TR_37 = RG_rl_208 ;
	7'h5a :
		TR_37 = RG_rl_208 ;
	7'h5b :
		TR_37 = RG_rl_208 ;
	7'h5c :
		TR_37 = RG_rl_208 ;
	7'h5d :
		TR_37 = RG_rl_208 ;
	7'h5e :
		TR_37 = RG_rl_208 ;
	7'h5f :
		TR_37 = RG_rl_208 ;
	7'h60 :
		TR_37 = RG_rl_208 ;
	7'h61 :
		TR_37 = RG_rl_208 ;
	7'h62 :
		TR_37 = RG_rl_208 ;
	7'h63 :
		TR_37 = RG_rl_208 ;
	7'h64 :
		TR_37 = RG_rl_208 ;
	7'h65 :
		TR_37 = RG_rl_208 ;
	7'h66 :
		TR_37 = RG_rl_208 ;
	7'h67 :
		TR_37 = RG_rl_208 ;
	7'h68 :
		TR_37 = RG_rl_208 ;
	7'h69 :
		TR_37 = RG_rl_208 ;
	7'h6a :
		TR_37 = RG_rl_208 ;
	7'h6b :
		TR_37 = RG_rl_208 ;
	7'h6c :
		TR_37 = RG_rl_208 ;
	7'h6d :
		TR_37 = RG_rl_208 ;
	7'h6e :
		TR_37 = RG_rl_208 ;
	7'h6f :
		TR_37 = RG_rl_208 ;
	7'h70 :
		TR_37 = RG_rl_208 ;
	7'h71 :
		TR_37 = RG_rl_208 ;
	7'h72 :
		TR_37 = RG_rl_208 ;
	7'h73 :
		TR_37 = RG_rl_208 ;
	7'h74 :
		TR_37 = RG_rl_208 ;
	7'h75 :
		TR_37 = RG_rl_208 ;
	7'h76 :
		TR_37 = RG_rl_208 ;
	7'h77 :
		TR_37 = RG_rl_208 ;
	7'h78 :
		TR_37 = RG_rl_208 ;
	7'h79 :
		TR_37 = RG_rl_208 ;
	7'h7a :
		TR_37 = RG_rl_208 ;
	7'h7b :
		TR_37 = RG_rl_208 ;
	7'h7c :
		TR_37 = RG_rl_208 ;
	7'h7d :
		TR_37 = RG_rl_208 ;
	7'h7e :
		TR_37 = RG_rl_208 ;
	7'h7f :
		TR_37 = RG_rl_208 ;
	default :
		TR_37 = 9'hx ;
	endcase
always @ ( RG_rl_209 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_38 = RG_rl_209 ;
	7'h01 :
		TR_38 = RG_rl_209 ;
	7'h02 :
		TR_38 = RG_rl_209 ;
	7'h03 :
		TR_38 = RG_rl_209 ;
	7'h04 :
		TR_38 = RG_rl_209 ;
	7'h05 :
		TR_38 = RG_rl_209 ;
	7'h06 :
		TR_38 = RG_rl_209 ;
	7'h07 :
		TR_38 = RG_rl_209 ;
	7'h08 :
		TR_38 = RG_rl_209 ;
	7'h09 :
		TR_38 = RG_rl_209 ;
	7'h0a :
		TR_38 = RG_rl_209 ;
	7'h0b :
		TR_38 = RG_rl_209 ;
	7'h0c :
		TR_38 = RG_rl_209 ;
	7'h0d :
		TR_38 = RG_rl_209 ;
	7'h0e :
		TR_38 = RG_rl_209 ;
	7'h0f :
		TR_38 = RG_rl_209 ;
	7'h10 :
		TR_38 = RG_rl_209 ;
	7'h11 :
		TR_38 = RG_rl_209 ;
	7'h12 :
		TR_38 = RG_rl_209 ;
	7'h13 :
		TR_38 = RG_rl_209 ;
	7'h14 :
		TR_38 = RG_rl_209 ;
	7'h15 :
		TR_38 = RG_rl_209 ;
	7'h16 :
		TR_38 = RG_rl_209 ;
	7'h17 :
		TR_38 = RG_rl_209 ;
	7'h18 :
		TR_38 = RG_rl_209 ;
	7'h19 :
		TR_38 = RG_rl_209 ;
	7'h1a :
		TR_38 = 9'h000 ;	// line#=../rle.cpp:68
	7'h1b :
		TR_38 = RG_rl_209 ;
	7'h1c :
		TR_38 = RG_rl_209 ;
	7'h1d :
		TR_38 = RG_rl_209 ;
	7'h1e :
		TR_38 = RG_rl_209 ;
	7'h1f :
		TR_38 = RG_rl_209 ;
	7'h20 :
		TR_38 = RG_rl_209 ;
	7'h21 :
		TR_38 = RG_rl_209 ;
	7'h22 :
		TR_38 = RG_rl_209 ;
	7'h23 :
		TR_38 = RG_rl_209 ;
	7'h24 :
		TR_38 = RG_rl_209 ;
	7'h25 :
		TR_38 = RG_rl_209 ;
	7'h26 :
		TR_38 = RG_rl_209 ;
	7'h27 :
		TR_38 = RG_rl_209 ;
	7'h28 :
		TR_38 = RG_rl_209 ;
	7'h29 :
		TR_38 = RG_rl_209 ;
	7'h2a :
		TR_38 = RG_rl_209 ;
	7'h2b :
		TR_38 = RG_rl_209 ;
	7'h2c :
		TR_38 = RG_rl_209 ;
	7'h2d :
		TR_38 = RG_rl_209 ;
	7'h2e :
		TR_38 = RG_rl_209 ;
	7'h2f :
		TR_38 = RG_rl_209 ;
	7'h30 :
		TR_38 = RG_rl_209 ;
	7'h31 :
		TR_38 = RG_rl_209 ;
	7'h32 :
		TR_38 = RG_rl_209 ;
	7'h33 :
		TR_38 = RG_rl_209 ;
	7'h34 :
		TR_38 = RG_rl_209 ;
	7'h35 :
		TR_38 = RG_rl_209 ;
	7'h36 :
		TR_38 = RG_rl_209 ;
	7'h37 :
		TR_38 = RG_rl_209 ;
	7'h38 :
		TR_38 = RG_rl_209 ;
	7'h39 :
		TR_38 = RG_rl_209 ;
	7'h3a :
		TR_38 = RG_rl_209 ;
	7'h3b :
		TR_38 = RG_rl_209 ;
	7'h3c :
		TR_38 = RG_rl_209 ;
	7'h3d :
		TR_38 = RG_rl_209 ;
	7'h3e :
		TR_38 = RG_rl_209 ;
	7'h3f :
		TR_38 = RG_rl_209 ;
	7'h40 :
		TR_38 = RG_rl_209 ;
	7'h41 :
		TR_38 = RG_rl_209 ;
	7'h42 :
		TR_38 = RG_rl_209 ;
	7'h43 :
		TR_38 = RG_rl_209 ;
	7'h44 :
		TR_38 = RG_rl_209 ;
	7'h45 :
		TR_38 = RG_rl_209 ;
	7'h46 :
		TR_38 = RG_rl_209 ;
	7'h47 :
		TR_38 = RG_rl_209 ;
	7'h48 :
		TR_38 = RG_rl_209 ;
	7'h49 :
		TR_38 = RG_rl_209 ;
	7'h4a :
		TR_38 = RG_rl_209 ;
	7'h4b :
		TR_38 = RG_rl_209 ;
	7'h4c :
		TR_38 = RG_rl_209 ;
	7'h4d :
		TR_38 = RG_rl_209 ;
	7'h4e :
		TR_38 = RG_rl_209 ;
	7'h4f :
		TR_38 = RG_rl_209 ;
	7'h50 :
		TR_38 = RG_rl_209 ;
	7'h51 :
		TR_38 = RG_rl_209 ;
	7'h52 :
		TR_38 = RG_rl_209 ;
	7'h53 :
		TR_38 = RG_rl_209 ;
	7'h54 :
		TR_38 = RG_rl_209 ;
	7'h55 :
		TR_38 = RG_rl_209 ;
	7'h56 :
		TR_38 = RG_rl_209 ;
	7'h57 :
		TR_38 = RG_rl_209 ;
	7'h58 :
		TR_38 = RG_rl_209 ;
	7'h59 :
		TR_38 = RG_rl_209 ;
	7'h5a :
		TR_38 = RG_rl_209 ;
	7'h5b :
		TR_38 = RG_rl_209 ;
	7'h5c :
		TR_38 = RG_rl_209 ;
	7'h5d :
		TR_38 = RG_rl_209 ;
	7'h5e :
		TR_38 = RG_rl_209 ;
	7'h5f :
		TR_38 = RG_rl_209 ;
	7'h60 :
		TR_38 = RG_rl_209 ;
	7'h61 :
		TR_38 = RG_rl_209 ;
	7'h62 :
		TR_38 = RG_rl_209 ;
	7'h63 :
		TR_38 = RG_rl_209 ;
	7'h64 :
		TR_38 = RG_rl_209 ;
	7'h65 :
		TR_38 = RG_rl_209 ;
	7'h66 :
		TR_38 = RG_rl_209 ;
	7'h67 :
		TR_38 = RG_rl_209 ;
	7'h68 :
		TR_38 = RG_rl_209 ;
	7'h69 :
		TR_38 = RG_rl_209 ;
	7'h6a :
		TR_38 = RG_rl_209 ;
	7'h6b :
		TR_38 = RG_rl_209 ;
	7'h6c :
		TR_38 = RG_rl_209 ;
	7'h6d :
		TR_38 = RG_rl_209 ;
	7'h6e :
		TR_38 = RG_rl_209 ;
	7'h6f :
		TR_38 = RG_rl_209 ;
	7'h70 :
		TR_38 = RG_rl_209 ;
	7'h71 :
		TR_38 = RG_rl_209 ;
	7'h72 :
		TR_38 = RG_rl_209 ;
	7'h73 :
		TR_38 = RG_rl_209 ;
	7'h74 :
		TR_38 = RG_rl_209 ;
	7'h75 :
		TR_38 = RG_rl_209 ;
	7'h76 :
		TR_38 = RG_rl_209 ;
	7'h77 :
		TR_38 = RG_rl_209 ;
	7'h78 :
		TR_38 = RG_rl_209 ;
	7'h79 :
		TR_38 = RG_rl_209 ;
	7'h7a :
		TR_38 = RG_rl_209 ;
	7'h7b :
		TR_38 = RG_rl_209 ;
	7'h7c :
		TR_38 = RG_rl_209 ;
	7'h7d :
		TR_38 = RG_rl_209 ;
	7'h7e :
		TR_38 = RG_rl_209 ;
	7'h7f :
		TR_38 = RG_rl_209 ;
	default :
		TR_38 = 9'hx ;
	endcase
always @ ( RG_rl_210 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_39 = RG_rl_210 ;
	7'h01 :
		TR_39 = RG_rl_210 ;
	7'h02 :
		TR_39 = RG_rl_210 ;
	7'h03 :
		TR_39 = RG_rl_210 ;
	7'h04 :
		TR_39 = RG_rl_210 ;
	7'h05 :
		TR_39 = RG_rl_210 ;
	7'h06 :
		TR_39 = RG_rl_210 ;
	7'h07 :
		TR_39 = RG_rl_210 ;
	7'h08 :
		TR_39 = RG_rl_210 ;
	7'h09 :
		TR_39 = RG_rl_210 ;
	7'h0a :
		TR_39 = RG_rl_210 ;
	7'h0b :
		TR_39 = RG_rl_210 ;
	7'h0c :
		TR_39 = RG_rl_210 ;
	7'h0d :
		TR_39 = RG_rl_210 ;
	7'h0e :
		TR_39 = RG_rl_210 ;
	7'h0f :
		TR_39 = RG_rl_210 ;
	7'h10 :
		TR_39 = RG_rl_210 ;
	7'h11 :
		TR_39 = RG_rl_210 ;
	7'h12 :
		TR_39 = RG_rl_210 ;
	7'h13 :
		TR_39 = RG_rl_210 ;
	7'h14 :
		TR_39 = RG_rl_210 ;
	7'h15 :
		TR_39 = RG_rl_210 ;
	7'h16 :
		TR_39 = RG_rl_210 ;
	7'h17 :
		TR_39 = RG_rl_210 ;
	7'h18 :
		TR_39 = RG_rl_210 ;
	7'h19 :
		TR_39 = RG_rl_210 ;
	7'h1a :
		TR_39 = RG_rl_210 ;
	7'h1b :
		TR_39 = 9'h000 ;	// line#=../rle.cpp:68
	7'h1c :
		TR_39 = RG_rl_210 ;
	7'h1d :
		TR_39 = RG_rl_210 ;
	7'h1e :
		TR_39 = RG_rl_210 ;
	7'h1f :
		TR_39 = RG_rl_210 ;
	7'h20 :
		TR_39 = RG_rl_210 ;
	7'h21 :
		TR_39 = RG_rl_210 ;
	7'h22 :
		TR_39 = RG_rl_210 ;
	7'h23 :
		TR_39 = RG_rl_210 ;
	7'h24 :
		TR_39 = RG_rl_210 ;
	7'h25 :
		TR_39 = RG_rl_210 ;
	7'h26 :
		TR_39 = RG_rl_210 ;
	7'h27 :
		TR_39 = RG_rl_210 ;
	7'h28 :
		TR_39 = RG_rl_210 ;
	7'h29 :
		TR_39 = RG_rl_210 ;
	7'h2a :
		TR_39 = RG_rl_210 ;
	7'h2b :
		TR_39 = RG_rl_210 ;
	7'h2c :
		TR_39 = RG_rl_210 ;
	7'h2d :
		TR_39 = RG_rl_210 ;
	7'h2e :
		TR_39 = RG_rl_210 ;
	7'h2f :
		TR_39 = RG_rl_210 ;
	7'h30 :
		TR_39 = RG_rl_210 ;
	7'h31 :
		TR_39 = RG_rl_210 ;
	7'h32 :
		TR_39 = RG_rl_210 ;
	7'h33 :
		TR_39 = RG_rl_210 ;
	7'h34 :
		TR_39 = RG_rl_210 ;
	7'h35 :
		TR_39 = RG_rl_210 ;
	7'h36 :
		TR_39 = RG_rl_210 ;
	7'h37 :
		TR_39 = RG_rl_210 ;
	7'h38 :
		TR_39 = RG_rl_210 ;
	7'h39 :
		TR_39 = RG_rl_210 ;
	7'h3a :
		TR_39 = RG_rl_210 ;
	7'h3b :
		TR_39 = RG_rl_210 ;
	7'h3c :
		TR_39 = RG_rl_210 ;
	7'h3d :
		TR_39 = RG_rl_210 ;
	7'h3e :
		TR_39 = RG_rl_210 ;
	7'h3f :
		TR_39 = RG_rl_210 ;
	7'h40 :
		TR_39 = RG_rl_210 ;
	7'h41 :
		TR_39 = RG_rl_210 ;
	7'h42 :
		TR_39 = RG_rl_210 ;
	7'h43 :
		TR_39 = RG_rl_210 ;
	7'h44 :
		TR_39 = RG_rl_210 ;
	7'h45 :
		TR_39 = RG_rl_210 ;
	7'h46 :
		TR_39 = RG_rl_210 ;
	7'h47 :
		TR_39 = RG_rl_210 ;
	7'h48 :
		TR_39 = RG_rl_210 ;
	7'h49 :
		TR_39 = RG_rl_210 ;
	7'h4a :
		TR_39 = RG_rl_210 ;
	7'h4b :
		TR_39 = RG_rl_210 ;
	7'h4c :
		TR_39 = RG_rl_210 ;
	7'h4d :
		TR_39 = RG_rl_210 ;
	7'h4e :
		TR_39 = RG_rl_210 ;
	7'h4f :
		TR_39 = RG_rl_210 ;
	7'h50 :
		TR_39 = RG_rl_210 ;
	7'h51 :
		TR_39 = RG_rl_210 ;
	7'h52 :
		TR_39 = RG_rl_210 ;
	7'h53 :
		TR_39 = RG_rl_210 ;
	7'h54 :
		TR_39 = RG_rl_210 ;
	7'h55 :
		TR_39 = RG_rl_210 ;
	7'h56 :
		TR_39 = RG_rl_210 ;
	7'h57 :
		TR_39 = RG_rl_210 ;
	7'h58 :
		TR_39 = RG_rl_210 ;
	7'h59 :
		TR_39 = RG_rl_210 ;
	7'h5a :
		TR_39 = RG_rl_210 ;
	7'h5b :
		TR_39 = RG_rl_210 ;
	7'h5c :
		TR_39 = RG_rl_210 ;
	7'h5d :
		TR_39 = RG_rl_210 ;
	7'h5e :
		TR_39 = RG_rl_210 ;
	7'h5f :
		TR_39 = RG_rl_210 ;
	7'h60 :
		TR_39 = RG_rl_210 ;
	7'h61 :
		TR_39 = RG_rl_210 ;
	7'h62 :
		TR_39 = RG_rl_210 ;
	7'h63 :
		TR_39 = RG_rl_210 ;
	7'h64 :
		TR_39 = RG_rl_210 ;
	7'h65 :
		TR_39 = RG_rl_210 ;
	7'h66 :
		TR_39 = RG_rl_210 ;
	7'h67 :
		TR_39 = RG_rl_210 ;
	7'h68 :
		TR_39 = RG_rl_210 ;
	7'h69 :
		TR_39 = RG_rl_210 ;
	7'h6a :
		TR_39 = RG_rl_210 ;
	7'h6b :
		TR_39 = RG_rl_210 ;
	7'h6c :
		TR_39 = RG_rl_210 ;
	7'h6d :
		TR_39 = RG_rl_210 ;
	7'h6e :
		TR_39 = RG_rl_210 ;
	7'h6f :
		TR_39 = RG_rl_210 ;
	7'h70 :
		TR_39 = RG_rl_210 ;
	7'h71 :
		TR_39 = RG_rl_210 ;
	7'h72 :
		TR_39 = RG_rl_210 ;
	7'h73 :
		TR_39 = RG_rl_210 ;
	7'h74 :
		TR_39 = RG_rl_210 ;
	7'h75 :
		TR_39 = RG_rl_210 ;
	7'h76 :
		TR_39 = RG_rl_210 ;
	7'h77 :
		TR_39 = RG_rl_210 ;
	7'h78 :
		TR_39 = RG_rl_210 ;
	7'h79 :
		TR_39 = RG_rl_210 ;
	7'h7a :
		TR_39 = RG_rl_210 ;
	7'h7b :
		TR_39 = RG_rl_210 ;
	7'h7c :
		TR_39 = RG_rl_210 ;
	7'h7d :
		TR_39 = RG_rl_210 ;
	7'h7e :
		TR_39 = RG_rl_210 ;
	7'h7f :
		TR_39 = RG_rl_210 ;
	default :
		TR_39 = 9'hx ;
	endcase
always @ ( RG_rl_211 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_40 = RG_rl_211 ;
	7'h01 :
		TR_40 = RG_rl_211 ;
	7'h02 :
		TR_40 = RG_rl_211 ;
	7'h03 :
		TR_40 = RG_rl_211 ;
	7'h04 :
		TR_40 = RG_rl_211 ;
	7'h05 :
		TR_40 = RG_rl_211 ;
	7'h06 :
		TR_40 = RG_rl_211 ;
	7'h07 :
		TR_40 = RG_rl_211 ;
	7'h08 :
		TR_40 = RG_rl_211 ;
	7'h09 :
		TR_40 = RG_rl_211 ;
	7'h0a :
		TR_40 = RG_rl_211 ;
	7'h0b :
		TR_40 = RG_rl_211 ;
	7'h0c :
		TR_40 = RG_rl_211 ;
	7'h0d :
		TR_40 = RG_rl_211 ;
	7'h0e :
		TR_40 = RG_rl_211 ;
	7'h0f :
		TR_40 = RG_rl_211 ;
	7'h10 :
		TR_40 = RG_rl_211 ;
	7'h11 :
		TR_40 = RG_rl_211 ;
	7'h12 :
		TR_40 = RG_rl_211 ;
	7'h13 :
		TR_40 = RG_rl_211 ;
	7'h14 :
		TR_40 = RG_rl_211 ;
	7'h15 :
		TR_40 = RG_rl_211 ;
	7'h16 :
		TR_40 = RG_rl_211 ;
	7'h17 :
		TR_40 = RG_rl_211 ;
	7'h18 :
		TR_40 = RG_rl_211 ;
	7'h19 :
		TR_40 = RG_rl_211 ;
	7'h1a :
		TR_40 = RG_rl_211 ;
	7'h1b :
		TR_40 = RG_rl_211 ;
	7'h1c :
		TR_40 = 9'h000 ;	// line#=../rle.cpp:68
	7'h1d :
		TR_40 = RG_rl_211 ;
	7'h1e :
		TR_40 = RG_rl_211 ;
	7'h1f :
		TR_40 = RG_rl_211 ;
	7'h20 :
		TR_40 = RG_rl_211 ;
	7'h21 :
		TR_40 = RG_rl_211 ;
	7'h22 :
		TR_40 = RG_rl_211 ;
	7'h23 :
		TR_40 = RG_rl_211 ;
	7'h24 :
		TR_40 = RG_rl_211 ;
	7'h25 :
		TR_40 = RG_rl_211 ;
	7'h26 :
		TR_40 = RG_rl_211 ;
	7'h27 :
		TR_40 = RG_rl_211 ;
	7'h28 :
		TR_40 = RG_rl_211 ;
	7'h29 :
		TR_40 = RG_rl_211 ;
	7'h2a :
		TR_40 = RG_rl_211 ;
	7'h2b :
		TR_40 = RG_rl_211 ;
	7'h2c :
		TR_40 = RG_rl_211 ;
	7'h2d :
		TR_40 = RG_rl_211 ;
	7'h2e :
		TR_40 = RG_rl_211 ;
	7'h2f :
		TR_40 = RG_rl_211 ;
	7'h30 :
		TR_40 = RG_rl_211 ;
	7'h31 :
		TR_40 = RG_rl_211 ;
	7'h32 :
		TR_40 = RG_rl_211 ;
	7'h33 :
		TR_40 = RG_rl_211 ;
	7'h34 :
		TR_40 = RG_rl_211 ;
	7'h35 :
		TR_40 = RG_rl_211 ;
	7'h36 :
		TR_40 = RG_rl_211 ;
	7'h37 :
		TR_40 = RG_rl_211 ;
	7'h38 :
		TR_40 = RG_rl_211 ;
	7'h39 :
		TR_40 = RG_rl_211 ;
	7'h3a :
		TR_40 = RG_rl_211 ;
	7'h3b :
		TR_40 = RG_rl_211 ;
	7'h3c :
		TR_40 = RG_rl_211 ;
	7'h3d :
		TR_40 = RG_rl_211 ;
	7'h3e :
		TR_40 = RG_rl_211 ;
	7'h3f :
		TR_40 = RG_rl_211 ;
	7'h40 :
		TR_40 = RG_rl_211 ;
	7'h41 :
		TR_40 = RG_rl_211 ;
	7'h42 :
		TR_40 = RG_rl_211 ;
	7'h43 :
		TR_40 = RG_rl_211 ;
	7'h44 :
		TR_40 = RG_rl_211 ;
	7'h45 :
		TR_40 = RG_rl_211 ;
	7'h46 :
		TR_40 = RG_rl_211 ;
	7'h47 :
		TR_40 = RG_rl_211 ;
	7'h48 :
		TR_40 = RG_rl_211 ;
	7'h49 :
		TR_40 = RG_rl_211 ;
	7'h4a :
		TR_40 = RG_rl_211 ;
	7'h4b :
		TR_40 = RG_rl_211 ;
	7'h4c :
		TR_40 = RG_rl_211 ;
	7'h4d :
		TR_40 = RG_rl_211 ;
	7'h4e :
		TR_40 = RG_rl_211 ;
	7'h4f :
		TR_40 = RG_rl_211 ;
	7'h50 :
		TR_40 = RG_rl_211 ;
	7'h51 :
		TR_40 = RG_rl_211 ;
	7'h52 :
		TR_40 = RG_rl_211 ;
	7'h53 :
		TR_40 = RG_rl_211 ;
	7'h54 :
		TR_40 = RG_rl_211 ;
	7'h55 :
		TR_40 = RG_rl_211 ;
	7'h56 :
		TR_40 = RG_rl_211 ;
	7'h57 :
		TR_40 = RG_rl_211 ;
	7'h58 :
		TR_40 = RG_rl_211 ;
	7'h59 :
		TR_40 = RG_rl_211 ;
	7'h5a :
		TR_40 = RG_rl_211 ;
	7'h5b :
		TR_40 = RG_rl_211 ;
	7'h5c :
		TR_40 = RG_rl_211 ;
	7'h5d :
		TR_40 = RG_rl_211 ;
	7'h5e :
		TR_40 = RG_rl_211 ;
	7'h5f :
		TR_40 = RG_rl_211 ;
	7'h60 :
		TR_40 = RG_rl_211 ;
	7'h61 :
		TR_40 = RG_rl_211 ;
	7'h62 :
		TR_40 = RG_rl_211 ;
	7'h63 :
		TR_40 = RG_rl_211 ;
	7'h64 :
		TR_40 = RG_rl_211 ;
	7'h65 :
		TR_40 = RG_rl_211 ;
	7'h66 :
		TR_40 = RG_rl_211 ;
	7'h67 :
		TR_40 = RG_rl_211 ;
	7'h68 :
		TR_40 = RG_rl_211 ;
	7'h69 :
		TR_40 = RG_rl_211 ;
	7'h6a :
		TR_40 = RG_rl_211 ;
	7'h6b :
		TR_40 = RG_rl_211 ;
	7'h6c :
		TR_40 = RG_rl_211 ;
	7'h6d :
		TR_40 = RG_rl_211 ;
	7'h6e :
		TR_40 = RG_rl_211 ;
	7'h6f :
		TR_40 = RG_rl_211 ;
	7'h70 :
		TR_40 = RG_rl_211 ;
	7'h71 :
		TR_40 = RG_rl_211 ;
	7'h72 :
		TR_40 = RG_rl_211 ;
	7'h73 :
		TR_40 = RG_rl_211 ;
	7'h74 :
		TR_40 = RG_rl_211 ;
	7'h75 :
		TR_40 = RG_rl_211 ;
	7'h76 :
		TR_40 = RG_rl_211 ;
	7'h77 :
		TR_40 = RG_rl_211 ;
	7'h78 :
		TR_40 = RG_rl_211 ;
	7'h79 :
		TR_40 = RG_rl_211 ;
	7'h7a :
		TR_40 = RG_rl_211 ;
	7'h7b :
		TR_40 = RG_rl_211 ;
	7'h7c :
		TR_40 = RG_rl_211 ;
	7'h7d :
		TR_40 = RG_rl_211 ;
	7'h7e :
		TR_40 = RG_rl_211 ;
	7'h7f :
		TR_40 = RG_rl_211 ;
	default :
		TR_40 = 9'hx ;
	endcase
always @ ( RG_rl_212 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_41 = RG_rl_212 ;
	7'h01 :
		TR_41 = RG_rl_212 ;
	7'h02 :
		TR_41 = RG_rl_212 ;
	7'h03 :
		TR_41 = RG_rl_212 ;
	7'h04 :
		TR_41 = RG_rl_212 ;
	7'h05 :
		TR_41 = RG_rl_212 ;
	7'h06 :
		TR_41 = RG_rl_212 ;
	7'h07 :
		TR_41 = RG_rl_212 ;
	7'h08 :
		TR_41 = RG_rl_212 ;
	7'h09 :
		TR_41 = RG_rl_212 ;
	7'h0a :
		TR_41 = RG_rl_212 ;
	7'h0b :
		TR_41 = RG_rl_212 ;
	7'h0c :
		TR_41 = RG_rl_212 ;
	7'h0d :
		TR_41 = RG_rl_212 ;
	7'h0e :
		TR_41 = RG_rl_212 ;
	7'h0f :
		TR_41 = RG_rl_212 ;
	7'h10 :
		TR_41 = RG_rl_212 ;
	7'h11 :
		TR_41 = RG_rl_212 ;
	7'h12 :
		TR_41 = RG_rl_212 ;
	7'h13 :
		TR_41 = RG_rl_212 ;
	7'h14 :
		TR_41 = RG_rl_212 ;
	7'h15 :
		TR_41 = RG_rl_212 ;
	7'h16 :
		TR_41 = RG_rl_212 ;
	7'h17 :
		TR_41 = RG_rl_212 ;
	7'h18 :
		TR_41 = RG_rl_212 ;
	7'h19 :
		TR_41 = RG_rl_212 ;
	7'h1a :
		TR_41 = RG_rl_212 ;
	7'h1b :
		TR_41 = RG_rl_212 ;
	7'h1c :
		TR_41 = RG_rl_212 ;
	7'h1d :
		TR_41 = 9'h000 ;	// line#=../rle.cpp:68
	7'h1e :
		TR_41 = RG_rl_212 ;
	7'h1f :
		TR_41 = RG_rl_212 ;
	7'h20 :
		TR_41 = RG_rl_212 ;
	7'h21 :
		TR_41 = RG_rl_212 ;
	7'h22 :
		TR_41 = RG_rl_212 ;
	7'h23 :
		TR_41 = RG_rl_212 ;
	7'h24 :
		TR_41 = RG_rl_212 ;
	7'h25 :
		TR_41 = RG_rl_212 ;
	7'h26 :
		TR_41 = RG_rl_212 ;
	7'h27 :
		TR_41 = RG_rl_212 ;
	7'h28 :
		TR_41 = RG_rl_212 ;
	7'h29 :
		TR_41 = RG_rl_212 ;
	7'h2a :
		TR_41 = RG_rl_212 ;
	7'h2b :
		TR_41 = RG_rl_212 ;
	7'h2c :
		TR_41 = RG_rl_212 ;
	7'h2d :
		TR_41 = RG_rl_212 ;
	7'h2e :
		TR_41 = RG_rl_212 ;
	7'h2f :
		TR_41 = RG_rl_212 ;
	7'h30 :
		TR_41 = RG_rl_212 ;
	7'h31 :
		TR_41 = RG_rl_212 ;
	7'h32 :
		TR_41 = RG_rl_212 ;
	7'h33 :
		TR_41 = RG_rl_212 ;
	7'h34 :
		TR_41 = RG_rl_212 ;
	7'h35 :
		TR_41 = RG_rl_212 ;
	7'h36 :
		TR_41 = RG_rl_212 ;
	7'h37 :
		TR_41 = RG_rl_212 ;
	7'h38 :
		TR_41 = RG_rl_212 ;
	7'h39 :
		TR_41 = RG_rl_212 ;
	7'h3a :
		TR_41 = RG_rl_212 ;
	7'h3b :
		TR_41 = RG_rl_212 ;
	7'h3c :
		TR_41 = RG_rl_212 ;
	7'h3d :
		TR_41 = RG_rl_212 ;
	7'h3e :
		TR_41 = RG_rl_212 ;
	7'h3f :
		TR_41 = RG_rl_212 ;
	7'h40 :
		TR_41 = RG_rl_212 ;
	7'h41 :
		TR_41 = RG_rl_212 ;
	7'h42 :
		TR_41 = RG_rl_212 ;
	7'h43 :
		TR_41 = RG_rl_212 ;
	7'h44 :
		TR_41 = RG_rl_212 ;
	7'h45 :
		TR_41 = RG_rl_212 ;
	7'h46 :
		TR_41 = RG_rl_212 ;
	7'h47 :
		TR_41 = RG_rl_212 ;
	7'h48 :
		TR_41 = RG_rl_212 ;
	7'h49 :
		TR_41 = RG_rl_212 ;
	7'h4a :
		TR_41 = RG_rl_212 ;
	7'h4b :
		TR_41 = RG_rl_212 ;
	7'h4c :
		TR_41 = RG_rl_212 ;
	7'h4d :
		TR_41 = RG_rl_212 ;
	7'h4e :
		TR_41 = RG_rl_212 ;
	7'h4f :
		TR_41 = RG_rl_212 ;
	7'h50 :
		TR_41 = RG_rl_212 ;
	7'h51 :
		TR_41 = RG_rl_212 ;
	7'h52 :
		TR_41 = RG_rl_212 ;
	7'h53 :
		TR_41 = RG_rl_212 ;
	7'h54 :
		TR_41 = RG_rl_212 ;
	7'h55 :
		TR_41 = RG_rl_212 ;
	7'h56 :
		TR_41 = RG_rl_212 ;
	7'h57 :
		TR_41 = RG_rl_212 ;
	7'h58 :
		TR_41 = RG_rl_212 ;
	7'h59 :
		TR_41 = RG_rl_212 ;
	7'h5a :
		TR_41 = RG_rl_212 ;
	7'h5b :
		TR_41 = RG_rl_212 ;
	7'h5c :
		TR_41 = RG_rl_212 ;
	7'h5d :
		TR_41 = RG_rl_212 ;
	7'h5e :
		TR_41 = RG_rl_212 ;
	7'h5f :
		TR_41 = RG_rl_212 ;
	7'h60 :
		TR_41 = RG_rl_212 ;
	7'h61 :
		TR_41 = RG_rl_212 ;
	7'h62 :
		TR_41 = RG_rl_212 ;
	7'h63 :
		TR_41 = RG_rl_212 ;
	7'h64 :
		TR_41 = RG_rl_212 ;
	7'h65 :
		TR_41 = RG_rl_212 ;
	7'h66 :
		TR_41 = RG_rl_212 ;
	7'h67 :
		TR_41 = RG_rl_212 ;
	7'h68 :
		TR_41 = RG_rl_212 ;
	7'h69 :
		TR_41 = RG_rl_212 ;
	7'h6a :
		TR_41 = RG_rl_212 ;
	7'h6b :
		TR_41 = RG_rl_212 ;
	7'h6c :
		TR_41 = RG_rl_212 ;
	7'h6d :
		TR_41 = RG_rl_212 ;
	7'h6e :
		TR_41 = RG_rl_212 ;
	7'h6f :
		TR_41 = RG_rl_212 ;
	7'h70 :
		TR_41 = RG_rl_212 ;
	7'h71 :
		TR_41 = RG_rl_212 ;
	7'h72 :
		TR_41 = RG_rl_212 ;
	7'h73 :
		TR_41 = RG_rl_212 ;
	7'h74 :
		TR_41 = RG_rl_212 ;
	7'h75 :
		TR_41 = RG_rl_212 ;
	7'h76 :
		TR_41 = RG_rl_212 ;
	7'h77 :
		TR_41 = RG_rl_212 ;
	7'h78 :
		TR_41 = RG_rl_212 ;
	7'h79 :
		TR_41 = RG_rl_212 ;
	7'h7a :
		TR_41 = RG_rl_212 ;
	7'h7b :
		TR_41 = RG_rl_212 ;
	7'h7c :
		TR_41 = RG_rl_212 ;
	7'h7d :
		TR_41 = RG_rl_212 ;
	7'h7e :
		TR_41 = RG_rl_212 ;
	7'h7f :
		TR_41 = RG_rl_212 ;
	default :
		TR_41 = 9'hx ;
	endcase
always @ ( RG_rl_213 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_42 = RG_rl_213 ;
	7'h01 :
		TR_42 = RG_rl_213 ;
	7'h02 :
		TR_42 = RG_rl_213 ;
	7'h03 :
		TR_42 = RG_rl_213 ;
	7'h04 :
		TR_42 = RG_rl_213 ;
	7'h05 :
		TR_42 = RG_rl_213 ;
	7'h06 :
		TR_42 = RG_rl_213 ;
	7'h07 :
		TR_42 = RG_rl_213 ;
	7'h08 :
		TR_42 = RG_rl_213 ;
	7'h09 :
		TR_42 = RG_rl_213 ;
	7'h0a :
		TR_42 = RG_rl_213 ;
	7'h0b :
		TR_42 = RG_rl_213 ;
	7'h0c :
		TR_42 = RG_rl_213 ;
	7'h0d :
		TR_42 = RG_rl_213 ;
	7'h0e :
		TR_42 = RG_rl_213 ;
	7'h0f :
		TR_42 = RG_rl_213 ;
	7'h10 :
		TR_42 = RG_rl_213 ;
	7'h11 :
		TR_42 = RG_rl_213 ;
	7'h12 :
		TR_42 = RG_rl_213 ;
	7'h13 :
		TR_42 = RG_rl_213 ;
	7'h14 :
		TR_42 = RG_rl_213 ;
	7'h15 :
		TR_42 = RG_rl_213 ;
	7'h16 :
		TR_42 = RG_rl_213 ;
	7'h17 :
		TR_42 = RG_rl_213 ;
	7'h18 :
		TR_42 = RG_rl_213 ;
	7'h19 :
		TR_42 = RG_rl_213 ;
	7'h1a :
		TR_42 = RG_rl_213 ;
	7'h1b :
		TR_42 = RG_rl_213 ;
	7'h1c :
		TR_42 = RG_rl_213 ;
	7'h1d :
		TR_42 = RG_rl_213 ;
	7'h1e :
		TR_42 = 9'h000 ;	// line#=../rle.cpp:68
	7'h1f :
		TR_42 = RG_rl_213 ;
	7'h20 :
		TR_42 = RG_rl_213 ;
	7'h21 :
		TR_42 = RG_rl_213 ;
	7'h22 :
		TR_42 = RG_rl_213 ;
	7'h23 :
		TR_42 = RG_rl_213 ;
	7'h24 :
		TR_42 = RG_rl_213 ;
	7'h25 :
		TR_42 = RG_rl_213 ;
	7'h26 :
		TR_42 = RG_rl_213 ;
	7'h27 :
		TR_42 = RG_rl_213 ;
	7'h28 :
		TR_42 = RG_rl_213 ;
	7'h29 :
		TR_42 = RG_rl_213 ;
	7'h2a :
		TR_42 = RG_rl_213 ;
	7'h2b :
		TR_42 = RG_rl_213 ;
	7'h2c :
		TR_42 = RG_rl_213 ;
	7'h2d :
		TR_42 = RG_rl_213 ;
	7'h2e :
		TR_42 = RG_rl_213 ;
	7'h2f :
		TR_42 = RG_rl_213 ;
	7'h30 :
		TR_42 = RG_rl_213 ;
	7'h31 :
		TR_42 = RG_rl_213 ;
	7'h32 :
		TR_42 = RG_rl_213 ;
	7'h33 :
		TR_42 = RG_rl_213 ;
	7'h34 :
		TR_42 = RG_rl_213 ;
	7'h35 :
		TR_42 = RG_rl_213 ;
	7'h36 :
		TR_42 = RG_rl_213 ;
	7'h37 :
		TR_42 = RG_rl_213 ;
	7'h38 :
		TR_42 = RG_rl_213 ;
	7'h39 :
		TR_42 = RG_rl_213 ;
	7'h3a :
		TR_42 = RG_rl_213 ;
	7'h3b :
		TR_42 = RG_rl_213 ;
	7'h3c :
		TR_42 = RG_rl_213 ;
	7'h3d :
		TR_42 = RG_rl_213 ;
	7'h3e :
		TR_42 = RG_rl_213 ;
	7'h3f :
		TR_42 = RG_rl_213 ;
	7'h40 :
		TR_42 = RG_rl_213 ;
	7'h41 :
		TR_42 = RG_rl_213 ;
	7'h42 :
		TR_42 = RG_rl_213 ;
	7'h43 :
		TR_42 = RG_rl_213 ;
	7'h44 :
		TR_42 = RG_rl_213 ;
	7'h45 :
		TR_42 = RG_rl_213 ;
	7'h46 :
		TR_42 = RG_rl_213 ;
	7'h47 :
		TR_42 = RG_rl_213 ;
	7'h48 :
		TR_42 = RG_rl_213 ;
	7'h49 :
		TR_42 = RG_rl_213 ;
	7'h4a :
		TR_42 = RG_rl_213 ;
	7'h4b :
		TR_42 = RG_rl_213 ;
	7'h4c :
		TR_42 = RG_rl_213 ;
	7'h4d :
		TR_42 = RG_rl_213 ;
	7'h4e :
		TR_42 = RG_rl_213 ;
	7'h4f :
		TR_42 = RG_rl_213 ;
	7'h50 :
		TR_42 = RG_rl_213 ;
	7'h51 :
		TR_42 = RG_rl_213 ;
	7'h52 :
		TR_42 = RG_rl_213 ;
	7'h53 :
		TR_42 = RG_rl_213 ;
	7'h54 :
		TR_42 = RG_rl_213 ;
	7'h55 :
		TR_42 = RG_rl_213 ;
	7'h56 :
		TR_42 = RG_rl_213 ;
	7'h57 :
		TR_42 = RG_rl_213 ;
	7'h58 :
		TR_42 = RG_rl_213 ;
	7'h59 :
		TR_42 = RG_rl_213 ;
	7'h5a :
		TR_42 = RG_rl_213 ;
	7'h5b :
		TR_42 = RG_rl_213 ;
	7'h5c :
		TR_42 = RG_rl_213 ;
	7'h5d :
		TR_42 = RG_rl_213 ;
	7'h5e :
		TR_42 = RG_rl_213 ;
	7'h5f :
		TR_42 = RG_rl_213 ;
	7'h60 :
		TR_42 = RG_rl_213 ;
	7'h61 :
		TR_42 = RG_rl_213 ;
	7'h62 :
		TR_42 = RG_rl_213 ;
	7'h63 :
		TR_42 = RG_rl_213 ;
	7'h64 :
		TR_42 = RG_rl_213 ;
	7'h65 :
		TR_42 = RG_rl_213 ;
	7'h66 :
		TR_42 = RG_rl_213 ;
	7'h67 :
		TR_42 = RG_rl_213 ;
	7'h68 :
		TR_42 = RG_rl_213 ;
	7'h69 :
		TR_42 = RG_rl_213 ;
	7'h6a :
		TR_42 = RG_rl_213 ;
	7'h6b :
		TR_42 = RG_rl_213 ;
	7'h6c :
		TR_42 = RG_rl_213 ;
	7'h6d :
		TR_42 = RG_rl_213 ;
	7'h6e :
		TR_42 = RG_rl_213 ;
	7'h6f :
		TR_42 = RG_rl_213 ;
	7'h70 :
		TR_42 = RG_rl_213 ;
	7'h71 :
		TR_42 = RG_rl_213 ;
	7'h72 :
		TR_42 = RG_rl_213 ;
	7'h73 :
		TR_42 = RG_rl_213 ;
	7'h74 :
		TR_42 = RG_rl_213 ;
	7'h75 :
		TR_42 = RG_rl_213 ;
	7'h76 :
		TR_42 = RG_rl_213 ;
	7'h77 :
		TR_42 = RG_rl_213 ;
	7'h78 :
		TR_42 = RG_rl_213 ;
	7'h79 :
		TR_42 = RG_rl_213 ;
	7'h7a :
		TR_42 = RG_rl_213 ;
	7'h7b :
		TR_42 = RG_rl_213 ;
	7'h7c :
		TR_42 = RG_rl_213 ;
	7'h7d :
		TR_42 = RG_rl_213 ;
	7'h7e :
		TR_42 = RG_rl_213 ;
	7'h7f :
		TR_42 = RG_rl_213 ;
	default :
		TR_42 = 9'hx ;
	endcase
always @ ( RG_rl_214 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_43 = RG_rl_214 ;
	7'h01 :
		TR_43 = RG_rl_214 ;
	7'h02 :
		TR_43 = RG_rl_214 ;
	7'h03 :
		TR_43 = RG_rl_214 ;
	7'h04 :
		TR_43 = RG_rl_214 ;
	7'h05 :
		TR_43 = RG_rl_214 ;
	7'h06 :
		TR_43 = RG_rl_214 ;
	7'h07 :
		TR_43 = RG_rl_214 ;
	7'h08 :
		TR_43 = RG_rl_214 ;
	7'h09 :
		TR_43 = RG_rl_214 ;
	7'h0a :
		TR_43 = RG_rl_214 ;
	7'h0b :
		TR_43 = RG_rl_214 ;
	7'h0c :
		TR_43 = RG_rl_214 ;
	7'h0d :
		TR_43 = RG_rl_214 ;
	7'h0e :
		TR_43 = RG_rl_214 ;
	7'h0f :
		TR_43 = RG_rl_214 ;
	7'h10 :
		TR_43 = RG_rl_214 ;
	7'h11 :
		TR_43 = RG_rl_214 ;
	7'h12 :
		TR_43 = RG_rl_214 ;
	7'h13 :
		TR_43 = RG_rl_214 ;
	7'h14 :
		TR_43 = RG_rl_214 ;
	7'h15 :
		TR_43 = RG_rl_214 ;
	7'h16 :
		TR_43 = RG_rl_214 ;
	7'h17 :
		TR_43 = RG_rl_214 ;
	7'h18 :
		TR_43 = RG_rl_214 ;
	7'h19 :
		TR_43 = RG_rl_214 ;
	7'h1a :
		TR_43 = RG_rl_214 ;
	7'h1b :
		TR_43 = RG_rl_214 ;
	7'h1c :
		TR_43 = RG_rl_214 ;
	7'h1d :
		TR_43 = RG_rl_214 ;
	7'h1e :
		TR_43 = RG_rl_214 ;
	7'h1f :
		TR_43 = 9'h000 ;	// line#=../rle.cpp:68
	7'h20 :
		TR_43 = RG_rl_214 ;
	7'h21 :
		TR_43 = RG_rl_214 ;
	7'h22 :
		TR_43 = RG_rl_214 ;
	7'h23 :
		TR_43 = RG_rl_214 ;
	7'h24 :
		TR_43 = RG_rl_214 ;
	7'h25 :
		TR_43 = RG_rl_214 ;
	7'h26 :
		TR_43 = RG_rl_214 ;
	7'h27 :
		TR_43 = RG_rl_214 ;
	7'h28 :
		TR_43 = RG_rl_214 ;
	7'h29 :
		TR_43 = RG_rl_214 ;
	7'h2a :
		TR_43 = RG_rl_214 ;
	7'h2b :
		TR_43 = RG_rl_214 ;
	7'h2c :
		TR_43 = RG_rl_214 ;
	7'h2d :
		TR_43 = RG_rl_214 ;
	7'h2e :
		TR_43 = RG_rl_214 ;
	7'h2f :
		TR_43 = RG_rl_214 ;
	7'h30 :
		TR_43 = RG_rl_214 ;
	7'h31 :
		TR_43 = RG_rl_214 ;
	7'h32 :
		TR_43 = RG_rl_214 ;
	7'h33 :
		TR_43 = RG_rl_214 ;
	7'h34 :
		TR_43 = RG_rl_214 ;
	7'h35 :
		TR_43 = RG_rl_214 ;
	7'h36 :
		TR_43 = RG_rl_214 ;
	7'h37 :
		TR_43 = RG_rl_214 ;
	7'h38 :
		TR_43 = RG_rl_214 ;
	7'h39 :
		TR_43 = RG_rl_214 ;
	7'h3a :
		TR_43 = RG_rl_214 ;
	7'h3b :
		TR_43 = RG_rl_214 ;
	7'h3c :
		TR_43 = RG_rl_214 ;
	7'h3d :
		TR_43 = RG_rl_214 ;
	7'h3e :
		TR_43 = RG_rl_214 ;
	7'h3f :
		TR_43 = RG_rl_214 ;
	7'h40 :
		TR_43 = RG_rl_214 ;
	7'h41 :
		TR_43 = RG_rl_214 ;
	7'h42 :
		TR_43 = RG_rl_214 ;
	7'h43 :
		TR_43 = RG_rl_214 ;
	7'h44 :
		TR_43 = RG_rl_214 ;
	7'h45 :
		TR_43 = RG_rl_214 ;
	7'h46 :
		TR_43 = RG_rl_214 ;
	7'h47 :
		TR_43 = RG_rl_214 ;
	7'h48 :
		TR_43 = RG_rl_214 ;
	7'h49 :
		TR_43 = RG_rl_214 ;
	7'h4a :
		TR_43 = RG_rl_214 ;
	7'h4b :
		TR_43 = RG_rl_214 ;
	7'h4c :
		TR_43 = RG_rl_214 ;
	7'h4d :
		TR_43 = RG_rl_214 ;
	7'h4e :
		TR_43 = RG_rl_214 ;
	7'h4f :
		TR_43 = RG_rl_214 ;
	7'h50 :
		TR_43 = RG_rl_214 ;
	7'h51 :
		TR_43 = RG_rl_214 ;
	7'h52 :
		TR_43 = RG_rl_214 ;
	7'h53 :
		TR_43 = RG_rl_214 ;
	7'h54 :
		TR_43 = RG_rl_214 ;
	7'h55 :
		TR_43 = RG_rl_214 ;
	7'h56 :
		TR_43 = RG_rl_214 ;
	7'h57 :
		TR_43 = RG_rl_214 ;
	7'h58 :
		TR_43 = RG_rl_214 ;
	7'h59 :
		TR_43 = RG_rl_214 ;
	7'h5a :
		TR_43 = RG_rl_214 ;
	7'h5b :
		TR_43 = RG_rl_214 ;
	7'h5c :
		TR_43 = RG_rl_214 ;
	7'h5d :
		TR_43 = RG_rl_214 ;
	7'h5e :
		TR_43 = RG_rl_214 ;
	7'h5f :
		TR_43 = RG_rl_214 ;
	7'h60 :
		TR_43 = RG_rl_214 ;
	7'h61 :
		TR_43 = RG_rl_214 ;
	7'h62 :
		TR_43 = RG_rl_214 ;
	7'h63 :
		TR_43 = RG_rl_214 ;
	7'h64 :
		TR_43 = RG_rl_214 ;
	7'h65 :
		TR_43 = RG_rl_214 ;
	7'h66 :
		TR_43 = RG_rl_214 ;
	7'h67 :
		TR_43 = RG_rl_214 ;
	7'h68 :
		TR_43 = RG_rl_214 ;
	7'h69 :
		TR_43 = RG_rl_214 ;
	7'h6a :
		TR_43 = RG_rl_214 ;
	7'h6b :
		TR_43 = RG_rl_214 ;
	7'h6c :
		TR_43 = RG_rl_214 ;
	7'h6d :
		TR_43 = RG_rl_214 ;
	7'h6e :
		TR_43 = RG_rl_214 ;
	7'h6f :
		TR_43 = RG_rl_214 ;
	7'h70 :
		TR_43 = RG_rl_214 ;
	7'h71 :
		TR_43 = RG_rl_214 ;
	7'h72 :
		TR_43 = RG_rl_214 ;
	7'h73 :
		TR_43 = RG_rl_214 ;
	7'h74 :
		TR_43 = RG_rl_214 ;
	7'h75 :
		TR_43 = RG_rl_214 ;
	7'h76 :
		TR_43 = RG_rl_214 ;
	7'h77 :
		TR_43 = RG_rl_214 ;
	7'h78 :
		TR_43 = RG_rl_214 ;
	7'h79 :
		TR_43 = RG_rl_214 ;
	7'h7a :
		TR_43 = RG_rl_214 ;
	7'h7b :
		TR_43 = RG_rl_214 ;
	7'h7c :
		TR_43 = RG_rl_214 ;
	7'h7d :
		TR_43 = RG_rl_214 ;
	7'h7e :
		TR_43 = RG_rl_214 ;
	7'h7f :
		TR_43 = RG_rl_214 ;
	default :
		TR_43 = 9'hx ;
	endcase
always @ ( RG_rl_215 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_44 = RG_rl_215 ;
	7'h01 :
		TR_44 = RG_rl_215 ;
	7'h02 :
		TR_44 = RG_rl_215 ;
	7'h03 :
		TR_44 = RG_rl_215 ;
	7'h04 :
		TR_44 = RG_rl_215 ;
	7'h05 :
		TR_44 = RG_rl_215 ;
	7'h06 :
		TR_44 = RG_rl_215 ;
	7'h07 :
		TR_44 = RG_rl_215 ;
	7'h08 :
		TR_44 = RG_rl_215 ;
	7'h09 :
		TR_44 = RG_rl_215 ;
	7'h0a :
		TR_44 = RG_rl_215 ;
	7'h0b :
		TR_44 = RG_rl_215 ;
	7'h0c :
		TR_44 = RG_rl_215 ;
	7'h0d :
		TR_44 = RG_rl_215 ;
	7'h0e :
		TR_44 = RG_rl_215 ;
	7'h0f :
		TR_44 = RG_rl_215 ;
	7'h10 :
		TR_44 = RG_rl_215 ;
	7'h11 :
		TR_44 = RG_rl_215 ;
	7'h12 :
		TR_44 = RG_rl_215 ;
	7'h13 :
		TR_44 = RG_rl_215 ;
	7'h14 :
		TR_44 = RG_rl_215 ;
	7'h15 :
		TR_44 = RG_rl_215 ;
	7'h16 :
		TR_44 = RG_rl_215 ;
	7'h17 :
		TR_44 = RG_rl_215 ;
	7'h18 :
		TR_44 = RG_rl_215 ;
	7'h19 :
		TR_44 = RG_rl_215 ;
	7'h1a :
		TR_44 = RG_rl_215 ;
	7'h1b :
		TR_44 = RG_rl_215 ;
	7'h1c :
		TR_44 = RG_rl_215 ;
	7'h1d :
		TR_44 = RG_rl_215 ;
	7'h1e :
		TR_44 = RG_rl_215 ;
	7'h1f :
		TR_44 = RG_rl_215 ;
	7'h20 :
		TR_44 = 9'h000 ;	// line#=../rle.cpp:68
	7'h21 :
		TR_44 = RG_rl_215 ;
	7'h22 :
		TR_44 = RG_rl_215 ;
	7'h23 :
		TR_44 = RG_rl_215 ;
	7'h24 :
		TR_44 = RG_rl_215 ;
	7'h25 :
		TR_44 = RG_rl_215 ;
	7'h26 :
		TR_44 = RG_rl_215 ;
	7'h27 :
		TR_44 = RG_rl_215 ;
	7'h28 :
		TR_44 = RG_rl_215 ;
	7'h29 :
		TR_44 = RG_rl_215 ;
	7'h2a :
		TR_44 = RG_rl_215 ;
	7'h2b :
		TR_44 = RG_rl_215 ;
	7'h2c :
		TR_44 = RG_rl_215 ;
	7'h2d :
		TR_44 = RG_rl_215 ;
	7'h2e :
		TR_44 = RG_rl_215 ;
	7'h2f :
		TR_44 = RG_rl_215 ;
	7'h30 :
		TR_44 = RG_rl_215 ;
	7'h31 :
		TR_44 = RG_rl_215 ;
	7'h32 :
		TR_44 = RG_rl_215 ;
	7'h33 :
		TR_44 = RG_rl_215 ;
	7'h34 :
		TR_44 = RG_rl_215 ;
	7'h35 :
		TR_44 = RG_rl_215 ;
	7'h36 :
		TR_44 = RG_rl_215 ;
	7'h37 :
		TR_44 = RG_rl_215 ;
	7'h38 :
		TR_44 = RG_rl_215 ;
	7'h39 :
		TR_44 = RG_rl_215 ;
	7'h3a :
		TR_44 = RG_rl_215 ;
	7'h3b :
		TR_44 = RG_rl_215 ;
	7'h3c :
		TR_44 = RG_rl_215 ;
	7'h3d :
		TR_44 = RG_rl_215 ;
	7'h3e :
		TR_44 = RG_rl_215 ;
	7'h3f :
		TR_44 = RG_rl_215 ;
	7'h40 :
		TR_44 = RG_rl_215 ;
	7'h41 :
		TR_44 = RG_rl_215 ;
	7'h42 :
		TR_44 = RG_rl_215 ;
	7'h43 :
		TR_44 = RG_rl_215 ;
	7'h44 :
		TR_44 = RG_rl_215 ;
	7'h45 :
		TR_44 = RG_rl_215 ;
	7'h46 :
		TR_44 = RG_rl_215 ;
	7'h47 :
		TR_44 = RG_rl_215 ;
	7'h48 :
		TR_44 = RG_rl_215 ;
	7'h49 :
		TR_44 = RG_rl_215 ;
	7'h4a :
		TR_44 = RG_rl_215 ;
	7'h4b :
		TR_44 = RG_rl_215 ;
	7'h4c :
		TR_44 = RG_rl_215 ;
	7'h4d :
		TR_44 = RG_rl_215 ;
	7'h4e :
		TR_44 = RG_rl_215 ;
	7'h4f :
		TR_44 = RG_rl_215 ;
	7'h50 :
		TR_44 = RG_rl_215 ;
	7'h51 :
		TR_44 = RG_rl_215 ;
	7'h52 :
		TR_44 = RG_rl_215 ;
	7'h53 :
		TR_44 = RG_rl_215 ;
	7'h54 :
		TR_44 = RG_rl_215 ;
	7'h55 :
		TR_44 = RG_rl_215 ;
	7'h56 :
		TR_44 = RG_rl_215 ;
	7'h57 :
		TR_44 = RG_rl_215 ;
	7'h58 :
		TR_44 = RG_rl_215 ;
	7'h59 :
		TR_44 = RG_rl_215 ;
	7'h5a :
		TR_44 = RG_rl_215 ;
	7'h5b :
		TR_44 = RG_rl_215 ;
	7'h5c :
		TR_44 = RG_rl_215 ;
	7'h5d :
		TR_44 = RG_rl_215 ;
	7'h5e :
		TR_44 = RG_rl_215 ;
	7'h5f :
		TR_44 = RG_rl_215 ;
	7'h60 :
		TR_44 = RG_rl_215 ;
	7'h61 :
		TR_44 = RG_rl_215 ;
	7'h62 :
		TR_44 = RG_rl_215 ;
	7'h63 :
		TR_44 = RG_rl_215 ;
	7'h64 :
		TR_44 = RG_rl_215 ;
	7'h65 :
		TR_44 = RG_rl_215 ;
	7'h66 :
		TR_44 = RG_rl_215 ;
	7'h67 :
		TR_44 = RG_rl_215 ;
	7'h68 :
		TR_44 = RG_rl_215 ;
	7'h69 :
		TR_44 = RG_rl_215 ;
	7'h6a :
		TR_44 = RG_rl_215 ;
	7'h6b :
		TR_44 = RG_rl_215 ;
	7'h6c :
		TR_44 = RG_rl_215 ;
	7'h6d :
		TR_44 = RG_rl_215 ;
	7'h6e :
		TR_44 = RG_rl_215 ;
	7'h6f :
		TR_44 = RG_rl_215 ;
	7'h70 :
		TR_44 = RG_rl_215 ;
	7'h71 :
		TR_44 = RG_rl_215 ;
	7'h72 :
		TR_44 = RG_rl_215 ;
	7'h73 :
		TR_44 = RG_rl_215 ;
	7'h74 :
		TR_44 = RG_rl_215 ;
	7'h75 :
		TR_44 = RG_rl_215 ;
	7'h76 :
		TR_44 = RG_rl_215 ;
	7'h77 :
		TR_44 = RG_rl_215 ;
	7'h78 :
		TR_44 = RG_rl_215 ;
	7'h79 :
		TR_44 = RG_rl_215 ;
	7'h7a :
		TR_44 = RG_rl_215 ;
	7'h7b :
		TR_44 = RG_rl_215 ;
	7'h7c :
		TR_44 = RG_rl_215 ;
	7'h7d :
		TR_44 = RG_rl_215 ;
	7'h7e :
		TR_44 = RG_rl_215 ;
	7'h7f :
		TR_44 = RG_rl_215 ;
	default :
		TR_44 = 9'hx ;
	endcase
always @ ( RG_rl_216 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_45 = RG_rl_216 ;
	7'h01 :
		TR_45 = RG_rl_216 ;
	7'h02 :
		TR_45 = RG_rl_216 ;
	7'h03 :
		TR_45 = RG_rl_216 ;
	7'h04 :
		TR_45 = RG_rl_216 ;
	7'h05 :
		TR_45 = RG_rl_216 ;
	7'h06 :
		TR_45 = RG_rl_216 ;
	7'h07 :
		TR_45 = RG_rl_216 ;
	7'h08 :
		TR_45 = RG_rl_216 ;
	7'h09 :
		TR_45 = RG_rl_216 ;
	7'h0a :
		TR_45 = RG_rl_216 ;
	7'h0b :
		TR_45 = RG_rl_216 ;
	7'h0c :
		TR_45 = RG_rl_216 ;
	7'h0d :
		TR_45 = RG_rl_216 ;
	7'h0e :
		TR_45 = RG_rl_216 ;
	7'h0f :
		TR_45 = RG_rl_216 ;
	7'h10 :
		TR_45 = RG_rl_216 ;
	7'h11 :
		TR_45 = RG_rl_216 ;
	7'h12 :
		TR_45 = RG_rl_216 ;
	7'h13 :
		TR_45 = RG_rl_216 ;
	7'h14 :
		TR_45 = RG_rl_216 ;
	7'h15 :
		TR_45 = RG_rl_216 ;
	7'h16 :
		TR_45 = RG_rl_216 ;
	7'h17 :
		TR_45 = RG_rl_216 ;
	7'h18 :
		TR_45 = RG_rl_216 ;
	7'h19 :
		TR_45 = RG_rl_216 ;
	7'h1a :
		TR_45 = RG_rl_216 ;
	7'h1b :
		TR_45 = RG_rl_216 ;
	7'h1c :
		TR_45 = RG_rl_216 ;
	7'h1d :
		TR_45 = RG_rl_216 ;
	7'h1e :
		TR_45 = RG_rl_216 ;
	7'h1f :
		TR_45 = RG_rl_216 ;
	7'h20 :
		TR_45 = RG_rl_216 ;
	7'h21 :
		TR_45 = 9'h000 ;	// line#=../rle.cpp:68
	7'h22 :
		TR_45 = RG_rl_216 ;
	7'h23 :
		TR_45 = RG_rl_216 ;
	7'h24 :
		TR_45 = RG_rl_216 ;
	7'h25 :
		TR_45 = RG_rl_216 ;
	7'h26 :
		TR_45 = RG_rl_216 ;
	7'h27 :
		TR_45 = RG_rl_216 ;
	7'h28 :
		TR_45 = RG_rl_216 ;
	7'h29 :
		TR_45 = RG_rl_216 ;
	7'h2a :
		TR_45 = RG_rl_216 ;
	7'h2b :
		TR_45 = RG_rl_216 ;
	7'h2c :
		TR_45 = RG_rl_216 ;
	7'h2d :
		TR_45 = RG_rl_216 ;
	7'h2e :
		TR_45 = RG_rl_216 ;
	7'h2f :
		TR_45 = RG_rl_216 ;
	7'h30 :
		TR_45 = RG_rl_216 ;
	7'h31 :
		TR_45 = RG_rl_216 ;
	7'h32 :
		TR_45 = RG_rl_216 ;
	7'h33 :
		TR_45 = RG_rl_216 ;
	7'h34 :
		TR_45 = RG_rl_216 ;
	7'h35 :
		TR_45 = RG_rl_216 ;
	7'h36 :
		TR_45 = RG_rl_216 ;
	7'h37 :
		TR_45 = RG_rl_216 ;
	7'h38 :
		TR_45 = RG_rl_216 ;
	7'h39 :
		TR_45 = RG_rl_216 ;
	7'h3a :
		TR_45 = RG_rl_216 ;
	7'h3b :
		TR_45 = RG_rl_216 ;
	7'h3c :
		TR_45 = RG_rl_216 ;
	7'h3d :
		TR_45 = RG_rl_216 ;
	7'h3e :
		TR_45 = RG_rl_216 ;
	7'h3f :
		TR_45 = RG_rl_216 ;
	7'h40 :
		TR_45 = RG_rl_216 ;
	7'h41 :
		TR_45 = RG_rl_216 ;
	7'h42 :
		TR_45 = RG_rl_216 ;
	7'h43 :
		TR_45 = RG_rl_216 ;
	7'h44 :
		TR_45 = RG_rl_216 ;
	7'h45 :
		TR_45 = RG_rl_216 ;
	7'h46 :
		TR_45 = RG_rl_216 ;
	7'h47 :
		TR_45 = RG_rl_216 ;
	7'h48 :
		TR_45 = RG_rl_216 ;
	7'h49 :
		TR_45 = RG_rl_216 ;
	7'h4a :
		TR_45 = RG_rl_216 ;
	7'h4b :
		TR_45 = RG_rl_216 ;
	7'h4c :
		TR_45 = RG_rl_216 ;
	7'h4d :
		TR_45 = RG_rl_216 ;
	7'h4e :
		TR_45 = RG_rl_216 ;
	7'h4f :
		TR_45 = RG_rl_216 ;
	7'h50 :
		TR_45 = RG_rl_216 ;
	7'h51 :
		TR_45 = RG_rl_216 ;
	7'h52 :
		TR_45 = RG_rl_216 ;
	7'h53 :
		TR_45 = RG_rl_216 ;
	7'h54 :
		TR_45 = RG_rl_216 ;
	7'h55 :
		TR_45 = RG_rl_216 ;
	7'h56 :
		TR_45 = RG_rl_216 ;
	7'h57 :
		TR_45 = RG_rl_216 ;
	7'h58 :
		TR_45 = RG_rl_216 ;
	7'h59 :
		TR_45 = RG_rl_216 ;
	7'h5a :
		TR_45 = RG_rl_216 ;
	7'h5b :
		TR_45 = RG_rl_216 ;
	7'h5c :
		TR_45 = RG_rl_216 ;
	7'h5d :
		TR_45 = RG_rl_216 ;
	7'h5e :
		TR_45 = RG_rl_216 ;
	7'h5f :
		TR_45 = RG_rl_216 ;
	7'h60 :
		TR_45 = RG_rl_216 ;
	7'h61 :
		TR_45 = RG_rl_216 ;
	7'h62 :
		TR_45 = RG_rl_216 ;
	7'h63 :
		TR_45 = RG_rl_216 ;
	7'h64 :
		TR_45 = RG_rl_216 ;
	7'h65 :
		TR_45 = RG_rl_216 ;
	7'h66 :
		TR_45 = RG_rl_216 ;
	7'h67 :
		TR_45 = RG_rl_216 ;
	7'h68 :
		TR_45 = RG_rl_216 ;
	7'h69 :
		TR_45 = RG_rl_216 ;
	7'h6a :
		TR_45 = RG_rl_216 ;
	7'h6b :
		TR_45 = RG_rl_216 ;
	7'h6c :
		TR_45 = RG_rl_216 ;
	7'h6d :
		TR_45 = RG_rl_216 ;
	7'h6e :
		TR_45 = RG_rl_216 ;
	7'h6f :
		TR_45 = RG_rl_216 ;
	7'h70 :
		TR_45 = RG_rl_216 ;
	7'h71 :
		TR_45 = RG_rl_216 ;
	7'h72 :
		TR_45 = RG_rl_216 ;
	7'h73 :
		TR_45 = RG_rl_216 ;
	7'h74 :
		TR_45 = RG_rl_216 ;
	7'h75 :
		TR_45 = RG_rl_216 ;
	7'h76 :
		TR_45 = RG_rl_216 ;
	7'h77 :
		TR_45 = RG_rl_216 ;
	7'h78 :
		TR_45 = RG_rl_216 ;
	7'h79 :
		TR_45 = RG_rl_216 ;
	7'h7a :
		TR_45 = RG_rl_216 ;
	7'h7b :
		TR_45 = RG_rl_216 ;
	7'h7c :
		TR_45 = RG_rl_216 ;
	7'h7d :
		TR_45 = RG_rl_216 ;
	7'h7e :
		TR_45 = RG_rl_216 ;
	7'h7f :
		TR_45 = RG_rl_216 ;
	default :
		TR_45 = 9'hx ;
	endcase
always @ ( RG_rl_217 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_46 = RG_rl_217 ;
	7'h01 :
		TR_46 = RG_rl_217 ;
	7'h02 :
		TR_46 = RG_rl_217 ;
	7'h03 :
		TR_46 = RG_rl_217 ;
	7'h04 :
		TR_46 = RG_rl_217 ;
	7'h05 :
		TR_46 = RG_rl_217 ;
	7'h06 :
		TR_46 = RG_rl_217 ;
	7'h07 :
		TR_46 = RG_rl_217 ;
	7'h08 :
		TR_46 = RG_rl_217 ;
	7'h09 :
		TR_46 = RG_rl_217 ;
	7'h0a :
		TR_46 = RG_rl_217 ;
	7'h0b :
		TR_46 = RG_rl_217 ;
	7'h0c :
		TR_46 = RG_rl_217 ;
	7'h0d :
		TR_46 = RG_rl_217 ;
	7'h0e :
		TR_46 = RG_rl_217 ;
	7'h0f :
		TR_46 = RG_rl_217 ;
	7'h10 :
		TR_46 = RG_rl_217 ;
	7'h11 :
		TR_46 = RG_rl_217 ;
	7'h12 :
		TR_46 = RG_rl_217 ;
	7'h13 :
		TR_46 = RG_rl_217 ;
	7'h14 :
		TR_46 = RG_rl_217 ;
	7'h15 :
		TR_46 = RG_rl_217 ;
	7'h16 :
		TR_46 = RG_rl_217 ;
	7'h17 :
		TR_46 = RG_rl_217 ;
	7'h18 :
		TR_46 = RG_rl_217 ;
	7'h19 :
		TR_46 = RG_rl_217 ;
	7'h1a :
		TR_46 = RG_rl_217 ;
	7'h1b :
		TR_46 = RG_rl_217 ;
	7'h1c :
		TR_46 = RG_rl_217 ;
	7'h1d :
		TR_46 = RG_rl_217 ;
	7'h1e :
		TR_46 = RG_rl_217 ;
	7'h1f :
		TR_46 = RG_rl_217 ;
	7'h20 :
		TR_46 = RG_rl_217 ;
	7'h21 :
		TR_46 = RG_rl_217 ;
	7'h22 :
		TR_46 = 9'h000 ;	// line#=../rle.cpp:68
	7'h23 :
		TR_46 = RG_rl_217 ;
	7'h24 :
		TR_46 = RG_rl_217 ;
	7'h25 :
		TR_46 = RG_rl_217 ;
	7'h26 :
		TR_46 = RG_rl_217 ;
	7'h27 :
		TR_46 = RG_rl_217 ;
	7'h28 :
		TR_46 = RG_rl_217 ;
	7'h29 :
		TR_46 = RG_rl_217 ;
	7'h2a :
		TR_46 = RG_rl_217 ;
	7'h2b :
		TR_46 = RG_rl_217 ;
	7'h2c :
		TR_46 = RG_rl_217 ;
	7'h2d :
		TR_46 = RG_rl_217 ;
	7'h2e :
		TR_46 = RG_rl_217 ;
	7'h2f :
		TR_46 = RG_rl_217 ;
	7'h30 :
		TR_46 = RG_rl_217 ;
	7'h31 :
		TR_46 = RG_rl_217 ;
	7'h32 :
		TR_46 = RG_rl_217 ;
	7'h33 :
		TR_46 = RG_rl_217 ;
	7'h34 :
		TR_46 = RG_rl_217 ;
	7'h35 :
		TR_46 = RG_rl_217 ;
	7'h36 :
		TR_46 = RG_rl_217 ;
	7'h37 :
		TR_46 = RG_rl_217 ;
	7'h38 :
		TR_46 = RG_rl_217 ;
	7'h39 :
		TR_46 = RG_rl_217 ;
	7'h3a :
		TR_46 = RG_rl_217 ;
	7'h3b :
		TR_46 = RG_rl_217 ;
	7'h3c :
		TR_46 = RG_rl_217 ;
	7'h3d :
		TR_46 = RG_rl_217 ;
	7'h3e :
		TR_46 = RG_rl_217 ;
	7'h3f :
		TR_46 = RG_rl_217 ;
	7'h40 :
		TR_46 = RG_rl_217 ;
	7'h41 :
		TR_46 = RG_rl_217 ;
	7'h42 :
		TR_46 = RG_rl_217 ;
	7'h43 :
		TR_46 = RG_rl_217 ;
	7'h44 :
		TR_46 = RG_rl_217 ;
	7'h45 :
		TR_46 = RG_rl_217 ;
	7'h46 :
		TR_46 = RG_rl_217 ;
	7'h47 :
		TR_46 = RG_rl_217 ;
	7'h48 :
		TR_46 = RG_rl_217 ;
	7'h49 :
		TR_46 = RG_rl_217 ;
	7'h4a :
		TR_46 = RG_rl_217 ;
	7'h4b :
		TR_46 = RG_rl_217 ;
	7'h4c :
		TR_46 = RG_rl_217 ;
	7'h4d :
		TR_46 = RG_rl_217 ;
	7'h4e :
		TR_46 = RG_rl_217 ;
	7'h4f :
		TR_46 = RG_rl_217 ;
	7'h50 :
		TR_46 = RG_rl_217 ;
	7'h51 :
		TR_46 = RG_rl_217 ;
	7'h52 :
		TR_46 = RG_rl_217 ;
	7'h53 :
		TR_46 = RG_rl_217 ;
	7'h54 :
		TR_46 = RG_rl_217 ;
	7'h55 :
		TR_46 = RG_rl_217 ;
	7'h56 :
		TR_46 = RG_rl_217 ;
	7'h57 :
		TR_46 = RG_rl_217 ;
	7'h58 :
		TR_46 = RG_rl_217 ;
	7'h59 :
		TR_46 = RG_rl_217 ;
	7'h5a :
		TR_46 = RG_rl_217 ;
	7'h5b :
		TR_46 = RG_rl_217 ;
	7'h5c :
		TR_46 = RG_rl_217 ;
	7'h5d :
		TR_46 = RG_rl_217 ;
	7'h5e :
		TR_46 = RG_rl_217 ;
	7'h5f :
		TR_46 = RG_rl_217 ;
	7'h60 :
		TR_46 = RG_rl_217 ;
	7'h61 :
		TR_46 = RG_rl_217 ;
	7'h62 :
		TR_46 = RG_rl_217 ;
	7'h63 :
		TR_46 = RG_rl_217 ;
	7'h64 :
		TR_46 = RG_rl_217 ;
	7'h65 :
		TR_46 = RG_rl_217 ;
	7'h66 :
		TR_46 = RG_rl_217 ;
	7'h67 :
		TR_46 = RG_rl_217 ;
	7'h68 :
		TR_46 = RG_rl_217 ;
	7'h69 :
		TR_46 = RG_rl_217 ;
	7'h6a :
		TR_46 = RG_rl_217 ;
	7'h6b :
		TR_46 = RG_rl_217 ;
	7'h6c :
		TR_46 = RG_rl_217 ;
	7'h6d :
		TR_46 = RG_rl_217 ;
	7'h6e :
		TR_46 = RG_rl_217 ;
	7'h6f :
		TR_46 = RG_rl_217 ;
	7'h70 :
		TR_46 = RG_rl_217 ;
	7'h71 :
		TR_46 = RG_rl_217 ;
	7'h72 :
		TR_46 = RG_rl_217 ;
	7'h73 :
		TR_46 = RG_rl_217 ;
	7'h74 :
		TR_46 = RG_rl_217 ;
	7'h75 :
		TR_46 = RG_rl_217 ;
	7'h76 :
		TR_46 = RG_rl_217 ;
	7'h77 :
		TR_46 = RG_rl_217 ;
	7'h78 :
		TR_46 = RG_rl_217 ;
	7'h79 :
		TR_46 = RG_rl_217 ;
	7'h7a :
		TR_46 = RG_rl_217 ;
	7'h7b :
		TR_46 = RG_rl_217 ;
	7'h7c :
		TR_46 = RG_rl_217 ;
	7'h7d :
		TR_46 = RG_rl_217 ;
	7'h7e :
		TR_46 = RG_rl_217 ;
	7'h7f :
		TR_46 = RG_rl_217 ;
	default :
		TR_46 = 9'hx ;
	endcase
always @ ( RG_rl_218 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_47 = RG_rl_218 ;
	7'h01 :
		TR_47 = RG_rl_218 ;
	7'h02 :
		TR_47 = RG_rl_218 ;
	7'h03 :
		TR_47 = RG_rl_218 ;
	7'h04 :
		TR_47 = RG_rl_218 ;
	7'h05 :
		TR_47 = RG_rl_218 ;
	7'h06 :
		TR_47 = RG_rl_218 ;
	7'h07 :
		TR_47 = RG_rl_218 ;
	7'h08 :
		TR_47 = RG_rl_218 ;
	7'h09 :
		TR_47 = RG_rl_218 ;
	7'h0a :
		TR_47 = RG_rl_218 ;
	7'h0b :
		TR_47 = RG_rl_218 ;
	7'h0c :
		TR_47 = RG_rl_218 ;
	7'h0d :
		TR_47 = RG_rl_218 ;
	7'h0e :
		TR_47 = RG_rl_218 ;
	7'h0f :
		TR_47 = RG_rl_218 ;
	7'h10 :
		TR_47 = RG_rl_218 ;
	7'h11 :
		TR_47 = RG_rl_218 ;
	7'h12 :
		TR_47 = RG_rl_218 ;
	7'h13 :
		TR_47 = RG_rl_218 ;
	7'h14 :
		TR_47 = RG_rl_218 ;
	7'h15 :
		TR_47 = RG_rl_218 ;
	7'h16 :
		TR_47 = RG_rl_218 ;
	7'h17 :
		TR_47 = RG_rl_218 ;
	7'h18 :
		TR_47 = RG_rl_218 ;
	7'h19 :
		TR_47 = RG_rl_218 ;
	7'h1a :
		TR_47 = RG_rl_218 ;
	7'h1b :
		TR_47 = RG_rl_218 ;
	7'h1c :
		TR_47 = RG_rl_218 ;
	7'h1d :
		TR_47 = RG_rl_218 ;
	7'h1e :
		TR_47 = RG_rl_218 ;
	7'h1f :
		TR_47 = RG_rl_218 ;
	7'h20 :
		TR_47 = RG_rl_218 ;
	7'h21 :
		TR_47 = RG_rl_218 ;
	7'h22 :
		TR_47 = RG_rl_218 ;
	7'h23 :
		TR_47 = 9'h000 ;	// line#=../rle.cpp:68
	7'h24 :
		TR_47 = RG_rl_218 ;
	7'h25 :
		TR_47 = RG_rl_218 ;
	7'h26 :
		TR_47 = RG_rl_218 ;
	7'h27 :
		TR_47 = RG_rl_218 ;
	7'h28 :
		TR_47 = RG_rl_218 ;
	7'h29 :
		TR_47 = RG_rl_218 ;
	7'h2a :
		TR_47 = RG_rl_218 ;
	7'h2b :
		TR_47 = RG_rl_218 ;
	7'h2c :
		TR_47 = RG_rl_218 ;
	7'h2d :
		TR_47 = RG_rl_218 ;
	7'h2e :
		TR_47 = RG_rl_218 ;
	7'h2f :
		TR_47 = RG_rl_218 ;
	7'h30 :
		TR_47 = RG_rl_218 ;
	7'h31 :
		TR_47 = RG_rl_218 ;
	7'h32 :
		TR_47 = RG_rl_218 ;
	7'h33 :
		TR_47 = RG_rl_218 ;
	7'h34 :
		TR_47 = RG_rl_218 ;
	7'h35 :
		TR_47 = RG_rl_218 ;
	7'h36 :
		TR_47 = RG_rl_218 ;
	7'h37 :
		TR_47 = RG_rl_218 ;
	7'h38 :
		TR_47 = RG_rl_218 ;
	7'h39 :
		TR_47 = RG_rl_218 ;
	7'h3a :
		TR_47 = RG_rl_218 ;
	7'h3b :
		TR_47 = RG_rl_218 ;
	7'h3c :
		TR_47 = RG_rl_218 ;
	7'h3d :
		TR_47 = RG_rl_218 ;
	7'h3e :
		TR_47 = RG_rl_218 ;
	7'h3f :
		TR_47 = RG_rl_218 ;
	7'h40 :
		TR_47 = RG_rl_218 ;
	7'h41 :
		TR_47 = RG_rl_218 ;
	7'h42 :
		TR_47 = RG_rl_218 ;
	7'h43 :
		TR_47 = RG_rl_218 ;
	7'h44 :
		TR_47 = RG_rl_218 ;
	7'h45 :
		TR_47 = RG_rl_218 ;
	7'h46 :
		TR_47 = RG_rl_218 ;
	7'h47 :
		TR_47 = RG_rl_218 ;
	7'h48 :
		TR_47 = RG_rl_218 ;
	7'h49 :
		TR_47 = RG_rl_218 ;
	7'h4a :
		TR_47 = RG_rl_218 ;
	7'h4b :
		TR_47 = RG_rl_218 ;
	7'h4c :
		TR_47 = RG_rl_218 ;
	7'h4d :
		TR_47 = RG_rl_218 ;
	7'h4e :
		TR_47 = RG_rl_218 ;
	7'h4f :
		TR_47 = RG_rl_218 ;
	7'h50 :
		TR_47 = RG_rl_218 ;
	7'h51 :
		TR_47 = RG_rl_218 ;
	7'h52 :
		TR_47 = RG_rl_218 ;
	7'h53 :
		TR_47 = RG_rl_218 ;
	7'h54 :
		TR_47 = RG_rl_218 ;
	7'h55 :
		TR_47 = RG_rl_218 ;
	7'h56 :
		TR_47 = RG_rl_218 ;
	7'h57 :
		TR_47 = RG_rl_218 ;
	7'h58 :
		TR_47 = RG_rl_218 ;
	7'h59 :
		TR_47 = RG_rl_218 ;
	7'h5a :
		TR_47 = RG_rl_218 ;
	7'h5b :
		TR_47 = RG_rl_218 ;
	7'h5c :
		TR_47 = RG_rl_218 ;
	7'h5d :
		TR_47 = RG_rl_218 ;
	7'h5e :
		TR_47 = RG_rl_218 ;
	7'h5f :
		TR_47 = RG_rl_218 ;
	7'h60 :
		TR_47 = RG_rl_218 ;
	7'h61 :
		TR_47 = RG_rl_218 ;
	7'h62 :
		TR_47 = RG_rl_218 ;
	7'h63 :
		TR_47 = RG_rl_218 ;
	7'h64 :
		TR_47 = RG_rl_218 ;
	7'h65 :
		TR_47 = RG_rl_218 ;
	7'h66 :
		TR_47 = RG_rl_218 ;
	7'h67 :
		TR_47 = RG_rl_218 ;
	7'h68 :
		TR_47 = RG_rl_218 ;
	7'h69 :
		TR_47 = RG_rl_218 ;
	7'h6a :
		TR_47 = RG_rl_218 ;
	7'h6b :
		TR_47 = RG_rl_218 ;
	7'h6c :
		TR_47 = RG_rl_218 ;
	7'h6d :
		TR_47 = RG_rl_218 ;
	7'h6e :
		TR_47 = RG_rl_218 ;
	7'h6f :
		TR_47 = RG_rl_218 ;
	7'h70 :
		TR_47 = RG_rl_218 ;
	7'h71 :
		TR_47 = RG_rl_218 ;
	7'h72 :
		TR_47 = RG_rl_218 ;
	7'h73 :
		TR_47 = RG_rl_218 ;
	7'h74 :
		TR_47 = RG_rl_218 ;
	7'h75 :
		TR_47 = RG_rl_218 ;
	7'h76 :
		TR_47 = RG_rl_218 ;
	7'h77 :
		TR_47 = RG_rl_218 ;
	7'h78 :
		TR_47 = RG_rl_218 ;
	7'h79 :
		TR_47 = RG_rl_218 ;
	7'h7a :
		TR_47 = RG_rl_218 ;
	7'h7b :
		TR_47 = RG_rl_218 ;
	7'h7c :
		TR_47 = RG_rl_218 ;
	7'h7d :
		TR_47 = RG_rl_218 ;
	7'h7e :
		TR_47 = RG_rl_218 ;
	7'h7f :
		TR_47 = RG_rl_218 ;
	default :
		TR_47 = 9'hx ;
	endcase
always @ ( RG_rl_219 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_48 = RG_rl_219 ;
	7'h01 :
		TR_48 = RG_rl_219 ;
	7'h02 :
		TR_48 = RG_rl_219 ;
	7'h03 :
		TR_48 = RG_rl_219 ;
	7'h04 :
		TR_48 = RG_rl_219 ;
	7'h05 :
		TR_48 = RG_rl_219 ;
	7'h06 :
		TR_48 = RG_rl_219 ;
	7'h07 :
		TR_48 = RG_rl_219 ;
	7'h08 :
		TR_48 = RG_rl_219 ;
	7'h09 :
		TR_48 = RG_rl_219 ;
	7'h0a :
		TR_48 = RG_rl_219 ;
	7'h0b :
		TR_48 = RG_rl_219 ;
	7'h0c :
		TR_48 = RG_rl_219 ;
	7'h0d :
		TR_48 = RG_rl_219 ;
	7'h0e :
		TR_48 = RG_rl_219 ;
	7'h0f :
		TR_48 = RG_rl_219 ;
	7'h10 :
		TR_48 = RG_rl_219 ;
	7'h11 :
		TR_48 = RG_rl_219 ;
	7'h12 :
		TR_48 = RG_rl_219 ;
	7'h13 :
		TR_48 = RG_rl_219 ;
	7'h14 :
		TR_48 = RG_rl_219 ;
	7'h15 :
		TR_48 = RG_rl_219 ;
	7'h16 :
		TR_48 = RG_rl_219 ;
	7'h17 :
		TR_48 = RG_rl_219 ;
	7'h18 :
		TR_48 = RG_rl_219 ;
	7'h19 :
		TR_48 = RG_rl_219 ;
	7'h1a :
		TR_48 = RG_rl_219 ;
	7'h1b :
		TR_48 = RG_rl_219 ;
	7'h1c :
		TR_48 = RG_rl_219 ;
	7'h1d :
		TR_48 = RG_rl_219 ;
	7'h1e :
		TR_48 = RG_rl_219 ;
	7'h1f :
		TR_48 = RG_rl_219 ;
	7'h20 :
		TR_48 = RG_rl_219 ;
	7'h21 :
		TR_48 = RG_rl_219 ;
	7'h22 :
		TR_48 = RG_rl_219 ;
	7'h23 :
		TR_48 = RG_rl_219 ;
	7'h24 :
		TR_48 = 9'h000 ;	// line#=../rle.cpp:68
	7'h25 :
		TR_48 = RG_rl_219 ;
	7'h26 :
		TR_48 = RG_rl_219 ;
	7'h27 :
		TR_48 = RG_rl_219 ;
	7'h28 :
		TR_48 = RG_rl_219 ;
	7'h29 :
		TR_48 = RG_rl_219 ;
	7'h2a :
		TR_48 = RG_rl_219 ;
	7'h2b :
		TR_48 = RG_rl_219 ;
	7'h2c :
		TR_48 = RG_rl_219 ;
	7'h2d :
		TR_48 = RG_rl_219 ;
	7'h2e :
		TR_48 = RG_rl_219 ;
	7'h2f :
		TR_48 = RG_rl_219 ;
	7'h30 :
		TR_48 = RG_rl_219 ;
	7'h31 :
		TR_48 = RG_rl_219 ;
	7'h32 :
		TR_48 = RG_rl_219 ;
	7'h33 :
		TR_48 = RG_rl_219 ;
	7'h34 :
		TR_48 = RG_rl_219 ;
	7'h35 :
		TR_48 = RG_rl_219 ;
	7'h36 :
		TR_48 = RG_rl_219 ;
	7'h37 :
		TR_48 = RG_rl_219 ;
	7'h38 :
		TR_48 = RG_rl_219 ;
	7'h39 :
		TR_48 = RG_rl_219 ;
	7'h3a :
		TR_48 = RG_rl_219 ;
	7'h3b :
		TR_48 = RG_rl_219 ;
	7'h3c :
		TR_48 = RG_rl_219 ;
	7'h3d :
		TR_48 = RG_rl_219 ;
	7'h3e :
		TR_48 = RG_rl_219 ;
	7'h3f :
		TR_48 = RG_rl_219 ;
	7'h40 :
		TR_48 = RG_rl_219 ;
	7'h41 :
		TR_48 = RG_rl_219 ;
	7'h42 :
		TR_48 = RG_rl_219 ;
	7'h43 :
		TR_48 = RG_rl_219 ;
	7'h44 :
		TR_48 = RG_rl_219 ;
	7'h45 :
		TR_48 = RG_rl_219 ;
	7'h46 :
		TR_48 = RG_rl_219 ;
	7'h47 :
		TR_48 = RG_rl_219 ;
	7'h48 :
		TR_48 = RG_rl_219 ;
	7'h49 :
		TR_48 = RG_rl_219 ;
	7'h4a :
		TR_48 = RG_rl_219 ;
	7'h4b :
		TR_48 = RG_rl_219 ;
	7'h4c :
		TR_48 = RG_rl_219 ;
	7'h4d :
		TR_48 = RG_rl_219 ;
	7'h4e :
		TR_48 = RG_rl_219 ;
	7'h4f :
		TR_48 = RG_rl_219 ;
	7'h50 :
		TR_48 = RG_rl_219 ;
	7'h51 :
		TR_48 = RG_rl_219 ;
	7'h52 :
		TR_48 = RG_rl_219 ;
	7'h53 :
		TR_48 = RG_rl_219 ;
	7'h54 :
		TR_48 = RG_rl_219 ;
	7'h55 :
		TR_48 = RG_rl_219 ;
	7'h56 :
		TR_48 = RG_rl_219 ;
	7'h57 :
		TR_48 = RG_rl_219 ;
	7'h58 :
		TR_48 = RG_rl_219 ;
	7'h59 :
		TR_48 = RG_rl_219 ;
	7'h5a :
		TR_48 = RG_rl_219 ;
	7'h5b :
		TR_48 = RG_rl_219 ;
	7'h5c :
		TR_48 = RG_rl_219 ;
	7'h5d :
		TR_48 = RG_rl_219 ;
	7'h5e :
		TR_48 = RG_rl_219 ;
	7'h5f :
		TR_48 = RG_rl_219 ;
	7'h60 :
		TR_48 = RG_rl_219 ;
	7'h61 :
		TR_48 = RG_rl_219 ;
	7'h62 :
		TR_48 = RG_rl_219 ;
	7'h63 :
		TR_48 = RG_rl_219 ;
	7'h64 :
		TR_48 = RG_rl_219 ;
	7'h65 :
		TR_48 = RG_rl_219 ;
	7'h66 :
		TR_48 = RG_rl_219 ;
	7'h67 :
		TR_48 = RG_rl_219 ;
	7'h68 :
		TR_48 = RG_rl_219 ;
	7'h69 :
		TR_48 = RG_rl_219 ;
	7'h6a :
		TR_48 = RG_rl_219 ;
	7'h6b :
		TR_48 = RG_rl_219 ;
	7'h6c :
		TR_48 = RG_rl_219 ;
	7'h6d :
		TR_48 = RG_rl_219 ;
	7'h6e :
		TR_48 = RG_rl_219 ;
	7'h6f :
		TR_48 = RG_rl_219 ;
	7'h70 :
		TR_48 = RG_rl_219 ;
	7'h71 :
		TR_48 = RG_rl_219 ;
	7'h72 :
		TR_48 = RG_rl_219 ;
	7'h73 :
		TR_48 = RG_rl_219 ;
	7'h74 :
		TR_48 = RG_rl_219 ;
	7'h75 :
		TR_48 = RG_rl_219 ;
	7'h76 :
		TR_48 = RG_rl_219 ;
	7'h77 :
		TR_48 = RG_rl_219 ;
	7'h78 :
		TR_48 = RG_rl_219 ;
	7'h79 :
		TR_48 = RG_rl_219 ;
	7'h7a :
		TR_48 = RG_rl_219 ;
	7'h7b :
		TR_48 = RG_rl_219 ;
	7'h7c :
		TR_48 = RG_rl_219 ;
	7'h7d :
		TR_48 = RG_rl_219 ;
	7'h7e :
		TR_48 = RG_rl_219 ;
	7'h7f :
		TR_48 = RG_rl_219 ;
	default :
		TR_48 = 9'hx ;
	endcase
always @ ( RG_rl_220 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_49 = RG_rl_220 ;
	7'h01 :
		TR_49 = RG_rl_220 ;
	7'h02 :
		TR_49 = RG_rl_220 ;
	7'h03 :
		TR_49 = RG_rl_220 ;
	7'h04 :
		TR_49 = RG_rl_220 ;
	7'h05 :
		TR_49 = RG_rl_220 ;
	7'h06 :
		TR_49 = RG_rl_220 ;
	7'h07 :
		TR_49 = RG_rl_220 ;
	7'h08 :
		TR_49 = RG_rl_220 ;
	7'h09 :
		TR_49 = RG_rl_220 ;
	7'h0a :
		TR_49 = RG_rl_220 ;
	7'h0b :
		TR_49 = RG_rl_220 ;
	7'h0c :
		TR_49 = RG_rl_220 ;
	7'h0d :
		TR_49 = RG_rl_220 ;
	7'h0e :
		TR_49 = RG_rl_220 ;
	7'h0f :
		TR_49 = RG_rl_220 ;
	7'h10 :
		TR_49 = RG_rl_220 ;
	7'h11 :
		TR_49 = RG_rl_220 ;
	7'h12 :
		TR_49 = RG_rl_220 ;
	7'h13 :
		TR_49 = RG_rl_220 ;
	7'h14 :
		TR_49 = RG_rl_220 ;
	7'h15 :
		TR_49 = RG_rl_220 ;
	7'h16 :
		TR_49 = RG_rl_220 ;
	7'h17 :
		TR_49 = RG_rl_220 ;
	7'h18 :
		TR_49 = RG_rl_220 ;
	7'h19 :
		TR_49 = RG_rl_220 ;
	7'h1a :
		TR_49 = RG_rl_220 ;
	7'h1b :
		TR_49 = RG_rl_220 ;
	7'h1c :
		TR_49 = RG_rl_220 ;
	7'h1d :
		TR_49 = RG_rl_220 ;
	7'h1e :
		TR_49 = RG_rl_220 ;
	7'h1f :
		TR_49 = RG_rl_220 ;
	7'h20 :
		TR_49 = RG_rl_220 ;
	7'h21 :
		TR_49 = RG_rl_220 ;
	7'h22 :
		TR_49 = RG_rl_220 ;
	7'h23 :
		TR_49 = RG_rl_220 ;
	7'h24 :
		TR_49 = RG_rl_220 ;
	7'h25 :
		TR_49 = 9'h000 ;	// line#=../rle.cpp:68
	7'h26 :
		TR_49 = RG_rl_220 ;
	7'h27 :
		TR_49 = RG_rl_220 ;
	7'h28 :
		TR_49 = RG_rl_220 ;
	7'h29 :
		TR_49 = RG_rl_220 ;
	7'h2a :
		TR_49 = RG_rl_220 ;
	7'h2b :
		TR_49 = RG_rl_220 ;
	7'h2c :
		TR_49 = RG_rl_220 ;
	7'h2d :
		TR_49 = RG_rl_220 ;
	7'h2e :
		TR_49 = RG_rl_220 ;
	7'h2f :
		TR_49 = RG_rl_220 ;
	7'h30 :
		TR_49 = RG_rl_220 ;
	7'h31 :
		TR_49 = RG_rl_220 ;
	7'h32 :
		TR_49 = RG_rl_220 ;
	7'h33 :
		TR_49 = RG_rl_220 ;
	7'h34 :
		TR_49 = RG_rl_220 ;
	7'h35 :
		TR_49 = RG_rl_220 ;
	7'h36 :
		TR_49 = RG_rl_220 ;
	7'h37 :
		TR_49 = RG_rl_220 ;
	7'h38 :
		TR_49 = RG_rl_220 ;
	7'h39 :
		TR_49 = RG_rl_220 ;
	7'h3a :
		TR_49 = RG_rl_220 ;
	7'h3b :
		TR_49 = RG_rl_220 ;
	7'h3c :
		TR_49 = RG_rl_220 ;
	7'h3d :
		TR_49 = RG_rl_220 ;
	7'h3e :
		TR_49 = RG_rl_220 ;
	7'h3f :
		TR_49 = RG_rl_220 ;
	7'h40 :
		TR_49 = RG_rl_220 ;
	7'h41 :
		TR_49 = RG_rl_220 ;
	7'h42 :
		TR_49 = RG_rl_220 ;
	7'h43 :
		TR_49 = RG_rl_220 ;
	7'h44 :
		TR_49 = RG_rl_220 ;
	7'h45 :
		TR_49 = RG_rl_220 ;
	7'h46 :
		TR_49 = RG_rl_220 ;
	7'h47 :
		TR_49 = RG_rl_220 ;
	7'h48 :
		TR_49 = RG_rl_220 ;
	7'h49 :
		TR_49 = RG_rl_220 ;
	7'h4a :
		TR_49 = RG_rl_220 ;
	7'h4b :
		TR_49 = RG_rl_220 ;
	7'h4c :
		TR_49 = RG_rl_220 ;
	7'h4d :
		TR_49 = RG_rl_220 ;
	7'h4e :
		TR_49 = RG_rl_220 ;
	7'h4f :
		TR_49 = RG_rl_220 ;
	7'h50 :
		TR_49 = RG_rl_220 ;
	7'h51 :
		TR_49 = RG_rl_220 ;
	7'h52 :
		TR_49 = RG_rl_220 ;
	7'h53 :
		TR_49 = RG_rl_220 ;
	7'h54 :
		TR_49 = RG_rl_220 ;
	7'h55 :
		TR_49 = RG_rl_220 ;
	7'h56 :
		TR_49 = RG_rl_220 ;
	7'h57 :
		TR_49 = RG_rl_220 ;
	7'h58 :
		TR_49 = RG_rl_220 ;
	7'h59 :
		TR_49 = RG_rl_220 ;
	7'h5a :
		TR_49 = RG_rl_220 ;
	7'h5b :
		TR_49 = RG_rl_220 ;
	7'h5c :
		TR_49 = RG_rl_220 ;
	7'h5d :
		TR_49 = RG_rl_220 ;
	7'h5e :
		TR_49 = RG_rl_220 ;
	7'h5f :
		TR_49 = RG_rl_220 ;
	7'h60 :
		TR_49 = RG_rl_220 ;
	7'h61 :
		TR_49 = RG_rl_220 ;
	7'h62 :
		TR_49 = RG_rl_220 ;
	7'h63 :
		TR_49 = RG_rl_220 ;
	7'h64 :
		TR_49 = RG_rl_220 ;
	7'h65 :
		TR_49 = RG_rl_220 ;
	7'h66 :
		TR_49 = RG_rl_220 ;
	7'h67 :
		TR_49 = RG_rl_220 ;
	7'h68 :
		TR_49 = RG_rl_220 ;
	7'h69 :
		TR_49 = RG_rl_220 ;
	7'h6a :
		TR_49 = RG_rl_220 ;
	7'h6b :
		TR_49 = RG_rl_220 ;
	7'h6c :
		TR_49 = RG_rl_220 ;
	7'h6d :
		TR_49 = RG_rl_220 ;
	7'h6e :
		TR_49 = RG_rl_220 ;
	7'h6f :
		TR_49 = RG_rl_220 ;
	7'h70 :
		TR_49 = RG_rl_220 ;
	7'h71 :
		TR_49 = RG_rl_220 ;
	7'h72 :
		TR_49 = RG_rl_220 ;
	7'h73 :
		TR_49 = RG_rl_220 ;
	7'h74 :
		TR_49 = RG_rl_220 ;
	7'h75 :
		TR_49 = RG_rl_220 ;
	7'h76 :
		TR_49 = RG_rl_220 ;
	7'h77 :
		TR_49 = RG_rl_220 ;
	7'h78 :
		TR_49 = RG_rl_220 ;
	7'h79 :
		TR_49 = RG_rl_220 ;
	7'h7a :
		TR_49 = RG_rl_220 ;
	7'h7b :
		TR_49 = RG_rl_220 ;
	7'h7c :
		TR_49 = RG_rl_220 ;
	7'h7d :
		TR_49 = RG_rl_220 ;
	7'h7e :
		TR_49 = RG_rl_220 ;
	7'h7f :
		TR_49 = RG_rl_220 ;
	default :
		TR_49 = 9'hx ;
	endcase
always @ ( RG_rl_221 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_50 = RG_rl_221 ;
	7'h01 :
		TR_50 = RG_rl_221 ;
	7'h02 :
		TR_50 = RG_rl_221 ;
	7'h03 :
		TR_50 = RG_rl_221 ;
	7'h04 :
		TR_50 = RG_rl_221 ;
	7'h05 :
		TR_50 = RG_rl_221 ;
	7'h06 :
		TR_50 = RG_rl_221 ;
	7'h07 :
		TR_50 = RG_rl_221 ;
	7'h08 :
		TR_50 = RG_rl_221 ;
	7'h09 :
		TR_50 = RG_rl_221 ;
	7'h0a :
		TR_50 = RG_rl_221 ;
	7'h0b :
		TR_50 = RG_rl_221 ;
	7'h0c :
		TR_50 = RG_rl_221 ;
	7'h0d :
		TR_50 = RG_rl_221 ;
	7'h0e :
		TR_50 = RG_rl_221 ;
	7'h0f :
		TR_50 = RG_rl_221 ;
	7'h10 :
		TR_50 = RG_rl_221 ;
	7'h11 :
		TR_50 = RG_rl_221 ;
	7'h12 :
		TR_50 = RG_rl_221 ;
	7'h13 :
		TR_50 = RG_rl_221 ;
	7'h14 :
		TR_50 = RG_rl_221 ;
	7'h15 :
		TR_50 = RG_rl_221 ;
	7'h16 :
		TR_50 = RG_rl_221 ;
	7'h17 :
		TR_50 = RG_rl_221 ;
	7'h18 :
		TR_50 = RG_rl_221 ;
	7'h19 :
		TR_50 = RG_rl_221 ;
	7'h1a :
		TR_50 = RG_rl_221 ;
	7'h1b :
		TR_50 = RG_rl_221 ;
	7'h1c :
		TR_50 = RG_rl_221 ;
	7'h1d :
		TR_50 = RG_rl_221 ;
	7'h1e :
		TR_50 = RG_rl_221 ;
	7'h1f :
		TR_50 = RG_rl_221 ;
	7'h20 :
		TR_50 = RG_rl_221 ;
	7'h21 :
		TR_50 = RG_rl_221 ;
	7'h22 :
		TR_50 = RG_rl_221 ;
	7'h23 :
		TR_50 = RG_rl_221 ;
	7'h24 :
		TR_50 = RG_rl_221 ;
	7'h25 :
		TR_50 = RG_rl_221 ;
	7'h26 :
		TR_50 = 9'h000 ;	// line#=../rle.cpp:68
	7'h27 :
		TR_50 = RG_rl_221 ;
	7'h28 :
		TR_50 = RG_rl_221 ;
	7'h29 :
		TR_50 = RG_rl_221 ;
	7'h2a :
		TR_50 = RG_rl_221 ;
	7'h2b :
		TR_50 = RG_rl_221 ;
	7'h2c :
		TR_50 = RG_rl_221 ;
	7'h2d :
		TR_50 = RG_rl_221 ;
	7'h2e :
		TR_50 = RG_rl_221 ;
	7'h2f :
		TR_50 = RG_rl_221 ;
	7'h30 :
		TR_50 = RG_rl_221 ;
	7'h31 :
		TR_50 = RG_rl_221 ;
	7'h32 :
		TR_50 = RG_rl_221 ;
	7'h33 :
		TR_50 = RG_rl_221 ;
	7'h34 :
		TR_50 = RG_rl_221 ;
	7'h35 :
		TR_50 = RG_rl_221 ;
	7'h36 :
		TR_50 = RG_rl_221 ;
	7'h37 :
		TR_50 = RG_rl_221 ;
	7'h38 :
		TR_50 = RG_rl_221 ;
	7'h39 :
		TR_50 = RG_rl_221 ;
	7'h3a :
		TR_50 = RG_rl_221 ;
	7'h3b :
		TR_50 = RG_rl_221 ;
	7'h3c :
		TR_50 = RG_rl_221 ;
	7'h3d :
		TR_50 = RG_rl_221 ;
	7'h3e :
		TR_50 = RG_rl_221 ;
	7'h3f :
		TR_50 = RG_rl_221 ;
	7'h40 :
		TR_50 = RG_rl_221 ;
	7'h41 :
		TR_50 = RG_rl_221 ;
	7'h42 :
		TR_50 = RG_rl_221 ;
	7'h43 :
		TR_50 = RG_rl_221 ;
	7'h44 :
		TR_50 = RG_rl_221 ;
	7'h45 :
		TR_50 = RG_rl_221 ;
	7'h46 :
		TR_50 = RG_rl_221 ;
	7'h47 :
		TR_50 = RG_rl_221 ;
	7'h48 :
		TR_50 = RG_rl_221 ;
	7'h49 :
		TR_50 = RG_rl_221 ;
	7'h4a :
		TR_50 = RG_rl_221 ;
	7'h4b :
		TR_50 = RG_rl_221 ;
	7'h4c :
		TR_50 = RG_rl_221 ;
	7'h4d :
		TR_50 = RG_rl_221 ;
	7'h4e :
		TR_50 = RG_rl_221 ;
	7'h4f :
		TR_50 = RG_rl_221 ;
	7'h50 :
		TR_50 = RG_rl_221 ;
	7'h51 :
		TR_50 = RG_rl_221 ;
	7'h52 :
		TR_50 = RG_rl_221 ;
	7'h53 :
		TR_50 = RG_rl_221 ;
	7'h54 :
		TR_50 = RG_rl_221 ;
	7'h55 :
		TR_50 = RG_rl_221 ;
	7'h56 :
		TR_50 = RG_rl_221 ;
	7'h57 :
		TR_50 = RG_rl_221 ;
	7'h58 :
		TR_50 = RG_rl_221 ;
	7'h59 :
		TR_50 = RG_rl_221 ;
	7'h5a :
		TR_50 = RG_rl_221 ;
	7'h5b :
		TR_50 = RG_rl_221 ;
	7'h5c :
		TR_50 = RG_rl_221 ;
	7'h5d :
		TR_50 = RG_rl_221 ;
	7'h5e :
		TR_50 = RG_rl_221 ;
	7'h5f :
		TR_50 = RG_rl_221 ;
	7'h60 :
		TR_50 = RG_rl_221 ;
	7'h61 :
		TR_50 = RG_rl_221 ;
	7'h62 :
		TR_50 = RG_rl_221 ;
	7'h63 :
		TR_50 = RG_rl_221 ;
	7'h64 :
		TR_50 = RG_rl_221 ;
	7'h65 :
		TR_50 = RG_rl_221 ;
	7'h66 :
		TR_50 = RG_rl_221 ;
	7'h67 :
		TR_50 = RG_rl_221 ;
	7'h68 :
		TR_50 = RG_rl_221 ;
	7'h69 :
		TR_50 = RG_rl_221 ;
	7'h6a :
		TR_50 = RG_rl_221 ;
	7'h6b :
		TR_50 = RG_rl_221 ;
	7'h6c :
		TR_50 = RG_rl_221 ;
	7'h6d :
		TR_50 = RG_rl_221 ;
	7'h6e :
		TR_50 = RG_rl_221 ;
	7'h6f :
		TR_50 = RG_rl_221 ;
	7'h70 :
		TR_50 = RG_rl_221 ;
	7'h71 :
		TR_50 = RG_rl_221 ;
	7'h72 :
		TR_50 = RG_rl_221 ;
	7'h73 :
		TR_50 = RG_rl_221 ;
	7'h74 :
		TR_50 = RG_rl_221 ;
	7'h75 :
		TR_50 = RG_rl_221 ;
	7'h76 :
		TR_50 = RG_rl_221 ;
	7'h77 :
		TR_50 = RG_rl_221 ;
	7'h78 :
		TR_50 = RG_rl_221 ;
	7'h79 :
		TR_50 = RG_rl_221 ;
	7'h7a :
		TR_50 = RG_rl_221 ;
	7'h7b :
		TR_50 = RG_rl_221 ;
	7'h7c :
		TR_50 = RG_rl_221 ;
	7'h7d :
		TR_50 = RG_rl_221 ;
	7'h7e :
		TR_50 = RG_rl_221 ;
	7'h7f :
		TR_50 = RG_rl_221 ;
	default :
		TR_50 = 9'hx ;
	endcase
always @ ( RG_rl_222 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_51 = RG_rl_222 ;
	7'h01 :
		TR_51 = RG_rl_222 ;
	7'h02 :
		TR_51 = RG_rl_222 ;
	7'h03 :
		TR_51 = RG_rl_222 ;
	7'h04 :
		TR_51 = RG_rl_222 ;
	7'h05 :
		TR_51 = RG_rl_222 ;
	7'h06 :
		TR_51 = RG_rl_222 ;
	7'h07 :
		TR_51 = RG_rl_222 ;
	7'h08 :
		TR_51 = RG_rl_222 ;
	7'h09 :
		TR_51 = RG_rl_222 ;
	7'h0a :
		TR_51 = RG_rl_222 ;
	7'h0b :
		TR_51 = RG_rl_222 ;
	7'h0c :
		TR_51 = RG_rl_222 ;
	7'h0d :
		TR_51 = RG_rl_222 ;
	7'h0e :
		TR_51 = RG_rl_222 ;
	7'h0f :
		TR_51 = RG_rl_222 ;
	7'h10 :
		TR_51 = RG_rl_222 ;
	7'h11 :
		TR_51 = RG_rl_222 ;
	7'h12 :
		TR_51 = RG_rl_222 ;
	7'h13 :
		TR_51 = RG_rl_222 ;
	7'h14 :
		TR_51 = RG_rl_222 ;
	7'h15 :
		TR_51 = RG_rl_222 ;
	7'h16 :
		TR_51 = RG_rl_222 ;
	7'h17 :
		TR_51 = RG_rl_222 ;
	7'h18 :
		TR_51 = RG_rl_222 ;
	7'h19 :
		TR_51 = RG_rl_222 ;
	7'h1a :
		TR_51 = RG_rl_222 ;
	7'h1b :
		TR_51 = RG_rl_222 ;
	7'h1c :
		TR_51 = RG_rl_222 ;
	7'h1d :
		TR_51 = RG_rl_222 ;
	7'h1e :
		TR_51 = RG_rl_222 ;
	7'h1f :
		TR_51 = RG_rl_222 ;
	7'h20 :
		TR_51 = RG_rl_222 ;
	7'h21 :
		TR_51 = RG_rl_222 ;
	7'h22 :
		TR_51 = RG_rl_222 ;
	7'h23 :
		TR_51 = RG_rl_222 ;
	7'h24 :
		TR_51 = RG_rl_222 ;
	7'h25 :
		TR_51 = RG_rl_222 ;
	7'h26 :
		TR_51 = RG_rl_222 ;
	7'h27 :
		TR_51 = 9'h000 ;	// line#=../rle.cpp:68
	7'h28 :
		TR_51 = RG_rl_222 ;
	7'h29 :
		TR_51 = RG_rl_222 ;
	7'h2a :
		TR_51 = RG_rl_222 ;
	7'h2b :
		TR_51 = RG_rl_222 ;
	7'h2c :
		TR_51 = RG_rl_222 ;
	7'h2d :
		TR_51 = RG_rl_222 ;
	7'h2e :
		TR_51 = RG_rl_222 ;
	7'h2f :
		TR_51 = RG_rl_222 ;
	7'h30 :
		TR_51 = RG_rl_222 ;
	7'h31 :
		TR_51 = RG_rl_222 ;
	7'h32 :
		TR_51 = RG_rl_222 ;
	7'h33 :
		TR_51 = RG_rl_222 ;
	7'h34 :
		TR_51 = RG_rl_222 ;
	7'h35 :
		TR_51 = RG_rl_222 ;
	7'h36 :
		TR_51 = RG_rl_222 ;
	7'h37 :
		TR_51 = RG_rl_222 ;
	7'h38 :
		TR_51 = RG_rl_222 ;
	7'h39 :
		TR_51 = RG_rl_222 ;
	7'h3a :
		TR_51 = RG_rl_222 ;
	7'h3b :
		TR_51 = RG_rl_222 ;
	7'h3c :
		TR_51 = RG_rl_222 ;
	7'h3d :
		TR_51 = RG_rl_222 ;
	7'h3e :
		TR_51 = RG_rl_222 ;
	7'h3f :
		TR_51 = RG_rl_222 ;
	7'h40 :
		TR_51 = RG_rl_222 ;
	7'h41 :
		TR_51 = RG_rl_222 ;
	7'h42 :
		TR_51 = RG_rl_222 ;
	7'h43 :
		TR_51 = RG_rl_222 ;
	7'h44 :
		TR_51 = RG_rl_222 ;
	7'h45 :
		TR_51 = RG_rl_222 ;
	7'h46 :
		TR_51 = RG_rl_222 ;
	7'h47 :
		TR_51 = RG_rl_222 ;
	7'h48 :
		TR_51 = RG_rl_222 ;
	7'h49 :
		TR_51 = RG_rl_222 ;
	7'h4a :
		TR_51 = RG_rl_222 ;
	7'h4b :
		TR_51 = RG_rl_222 ;
	7'h4c :
		TR_51 = RG_rl_222 ;
	7'h4d :
		TR_51 = RG_rl_222 ;
	7'h4e :
		TR_51 = RG_rl_222 ;
	7'h4f :
		TR_51 = RG_rl_222 ;
	7'h50 :
		TR_51 = RG_rl_222 ;
	7'h51 :
		TR_51 = RG_rl_222 ;
	7'h52 :
		TR_51 = RG_rl_222 ;
	7'h53 :
		TR_51 = RG_rl_222 ;
	7'h54 :
		TR_51 = RG_rl_222 ;
	7'h55 :
		TR_51 = RG_rl_222 ;
	7'h56 :
		TR_51 = RG_rl_222 ;
	7'h57 :
		TR_51 = RG_rl_222 ;
	7'h58 :
		TR_51 = RG_rl_222 ;
	7'h59 :
		TR_51 = RG_rl_222 ;
	7'h5a :
		TR_51 = RG_rl_222 ;
	7'h5b :
		TR_51 = RG_rl_222 ;
	7'h5c :
		TR_51 = RG_rl_222 ;
	7'h5d :
		TR_51 = RG_rl_222 ;
	7'h5e :
		TR_51 = RG_rl_222 ;
	7'h5f :
		TR_51 = RG_rl_222 ;
	7'h60 :
		TR_51 = RG_rl_222 ;
	7'h61 :
		TR_51 = RG_rl_222 ;
	7'h62 :
		TR_51 = RG_rl_222 ;
	7'h63 :
		TR_51 = RG_rl_222 ;
	7'h64 :
		TR_51 = RG_rl_222 ;
	7'h65 :
		TR_51 = RG_rl_222 ;
	7'h66 :
		TR_51 = RG_rl_222 ;
	7'h67 :
		TR_51 = RG_rl_222 ;
	7'h68 :
		TR_51 = RG_rl_222 ;
	7'h69 :
		TR_51 = RG_rl_222 ;
	7'h6a :
		TR_51 = RG_rl_222 ;
	7'h6b :
		TR_51 = RG_rl_222 ;
	7'h6c :
		TR_51 = RG_rl_222 ;
	7'h6d :
		TR_51 = RG_rl_222 ;
	7'h6e :
		TR_51 = RG_rl_222 ;
	7'h6f :
		TR_51 = RG_rl_222 ;
	7'h70 :
		TR_51 = RG_rl_222 ;
	7'h71 :
		TR_51 = RG_rl_222 ;
	7'h72 :
		TR_51 = RG_rl_222 ;
	7'h73 :
		TR_51 = RG_rl_222 ;
	7'h74 :
		TR_51 = RG_rl_222 ;
	7'h75 :
		TR_51 = RG_rl_222 ;
	7'h76 :
		TR_51 = RG_rl_222 ;
	7'h77 :
		TR_51 = RG_rl_222 ;
	7'h78 :
		TR_51 = RG_rl_222 ;
	7'h79 :
		TR_51 = RG_rl_222 ;
	7'h7a :
		TR_51 = RG_rl_222 ;
	7'h7b :
		TR_51 = RG_rl_222 ;
	7'h7c :
		TR_51 = RG_rl_222 ;
	7'h7d :
		TR_51 = RG_rl_222 ;
	7'h7e :
		TR_51 = RG_rl_222 ;
	7'h7f :
		TR_51 = RG_rl_222 ;
	default :
		TR_51 = 9'hx ;
	endcase
always @ ( RG_rl_223 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_52 = RG_rl_223 ;
	7'h01 :
		TR_52 = RG_rl_223 ;
	7'h02 :
		TR_52 = RG_rl_223 ;
	7'h03 :
		TR_52 = RG_rl_223 ;
	7'h04 :
		TR_52 = RG_rl_223 ;
	7'h05 :
		TR_52 = RG_rl_223 ;
	7'h06 :
		TR_52 = RG_rl_223 ;
	7'h07 :
		TR_52 = RG_rl_223 ;
	7'h08 :
		TR_52 = RG_rl_223 ;
	7'h09 :
		TR_52 = RG_rl_223 ;
	7'h0a :
		TR_52 = RG_rl_223 ;
	7'h0b :
		TR_52 = RG_rl_223 ;
	7'h0c :
		TR_52 = RG_rl_223 ;
	7'h0d :
		TR_52 = RG_rl_223 ;
	7'h0e :
		TR_52 = RG_rl_223 ;
	7'h0f :
		TR_52 = RG_rl_223 ;
	7'h10 :
		TR_52 = RG_rl_223 ;
	7'h11 :
		TR_52 = RG_rl_223 ;
	7'h12 :
		TR_52 = RG_rl_223 ;
	7'h13 :
		TR_52 = RG_rl_223 ;
	7'h14 :
		TR_52 = RG_rl_223 ;
	7'h15 :
		TR_52 = RG_rl_223 ;
	7'h16 :
		TR_52 = RG_rl_223 ;
	7'h17 :
		TR_52 = RG_rl_223 ;
	7'h18 :
		TR_52 = RG_rl_223 ;
	7'h19 :
		TR_52 = RG_rl_223 ;
	7'h1a :
		TR_52 = RG_rl_223 ;
	7'h1b :
		TR_52 = RG_rl_223 ;
	7'h1c :
		TR_52 = RG_rl_223 ;
	7'h1d :
		TR_52 = RG_rl_223 ;
	7'h1e :
		TR_52 = RG_rl_223 ;
	7'h1f :
		TR_52 = RG_rl_223 ;
	7'h20 :
		TR_52 = RG_rl_223 ;
	7'h21 :
		TR_52 = RG_rl_223 ;
	7'h22 :
		TR_52 = RG_rl_223 ;
	7'h23 :
		TR_52 = RG_rl_223 ;
	7'h24 :
		TR_52 = RG_rl_223 ;
	7'h25 :
		TR_52 = RG_rl_223 ;
	7'h26 :
		TR_52 = RG_rl_223 ;
	7'h27 :
		TR_52 = RG_rl_223 ;
	7'h28 :
		TR_52 = 9'h000 ;	// line#=../rle.cpp:68
	7'h29 :
		TR_52 = RG_rl_223 ;
	7'h2a :
		TR_52 = RG_rl_223 ;
	7'h2b :
		TR_52 = RG_rl_223 ;
	7'h2c :
		TR_52 = RG_rl_223 ;
	7'h2d :
		TR_52 = RG_rl_223 ;
	7'h2e :
		TR_52 = RG_rl_223 ;
	7'h2f :
		TR_52 = RG_rl_223 ;
	7'h30 :
		TR_52 = RG_rl_223 ;
	7'h31 :
		TR_52 = RG_rl_223 ;
	7'h32 :
		TR_52 = RG_rl_223 ;
	7'h33 :
		TR_52 = RG_rl_223 ;
	7'h34 :
		TR_52 = RG_rl_223 ;
	7'h35 :
		TR_52 = RG_rl_223 ;
	7'h36 :
		TR_52 = RG_rl_223 ;
	7'h37 :
		TR_52 = RG_rl_223 ;
	7'h38 :
		TR_52 = RG_rl_223 ;
	7'h39 :
		TR_52 = RG_rl_223 ;
	7'h3a :
		TR_52 = RG_rl_223 ;
	7'h3b :
		TR_52 = RG_rl_223 ;
	7'h3c :
		TR_52 = RG_rl_223 ;
	7'h3d :
		TR_52 = RG_rl_223 ;
	7'h3e :
		TR_52 = RG_rl_223 ;
	7'h3f :
		TR_52 = RG_rl_223 ;
	7'h40 :
		TR_52 = RG_rl_223 ;
	7'h41 :
		TR_52 = RG_rl_223 ;
	7'h42 :
		TR_52 = RG_rl_223 ;
	7'h43 :
		TR_52 = RG_rl_223 ;
	7'h44 :
		TR_52 = RG_rl_223 ;
	7'h45 :
		TR_52 = RG_rl_223 ;
	7'h46 :
		TR_52 = RG_rl_223 ;
	7'h47 :
		TR_52 = RG_rl_223 ;
	7'h48 :
		TR_52 = RG_rl_223 ;
	7'h49 :
		TR_52 = RG_rl_223 ;
	7'h4a :
		TR_52 = RG_rl_223 ;
	7'h4b :
		TR_52 = RG_rl_223 ;
	7'h4c :
		TR_52 = RG_rl_223 ;
	7'h4d :
		TR_52 = RG_rl_223 ;
	7'h4e :
		TR_52 = RG_rl_223 ;
	7'h4f :
		TR_52 = RG_rl_223 ;
	7'h50 :
		TR_52 = RG_rl_223 ;
	7'h51 :
		TR_52 = RG_rl_223 ;
	7'h52 :
		TR_52 = RG_rl_223 ;
	7'h53 :
		TR_52 = RG_rl_223 ;
	7'h54 :
		TR_52 = RG_rl_223 ;
	7'h55 :
		TR_52 = RG_rl_223 ;
	7'h56 :
		TR_52 = RG_rl_223 ;
	7'h57 :
		TR_52 = RG_rl_223 ;
	7'h58 :
		TR_52 = RG_rl_223 ;
	7'h59 :
		TR_52 = RG_rl_223 ;
	7'h5a :
		TR_52 = RG_rl_223 ;
	7'h5b :
		TR_52 = RG_rl_223 ;
	7'h5c :
		TR_52 = RG_rl_223 ;
	7'h5d :
		TR_52 = RG_rl_223 ;
	7'h5e :
		TR_52 = RG_rl_223 ;
	7'h5f :
		TR_52 = RG_rl_223 ;
	7'h60 :
		TR_52 = RG_rl_223 ;
	7'h61 :
		TR_52 = RG_rl_223 ;
	7'h62 :
		TR_52 = RG_rl_223 ;
	7'h63 :
		TR_52 = RG_rl_223 ;
	7'h64 :
		TR_52 = RG_rl_223 ;
	7'h65 :
		TR_52 = RG_rl_223 ;
	7'h66 :
		TR_52 = RG_rl_223 ;
	7'h67 :
		TR_52 = RG_rl_223 ;
	7'h68 :
		TR_52 = RG_rl_223 ;
	7'h69 :
		TR_52 = RG_rl_223 ;
	7'h6a :
		TR_52 = RG_rl_223 ;
	7'h6b :
		TR_52 = RG_rl_223 ;
	7'h6c :
		TR_52 = RG_rl_223 ;
	7'h6d :
		TR_52 = RG_rl_223 ;
	7'h6e :
		TR_52 = RG_rl_223 ;
	7'h6f :
		TR_52 = RG_rl_223 ;
	7'h70 :
		TR_52 = RG_rl_223 ;
	7'h71 :
		TR_52 = RG_rl_223 ;
	7'h72 :
		TR_52 = RG_rl_223 ;
	7'h73 :
		TR_52 = RG_rl_223 ;
	7'h74 :
		TR_52 = RG_rl_223 ;
	7'h75 :
		TR_52 = RG_rl_223 ;
	7'h76 :
		TR_52 = RG_rl_223 ;
	7'h77 :
		TR_52 = RG_rl_223 ;
	7'h78 :
		TR_52 = RG_rl_223 ;
	7'h79 :
		TR_52 = RG_rl_223 ;
	7'h7a :
		TR_52 = RG_rl_223 ;
	7'h7b :
		TR_52 = RG_rl_223 ;
	7'h7c :
		TR_52 = RG_rl_223 ;
	7'h7d :
		TR_52 = RG_rl_223 ;
	7'h7e :
		TR_52 = RG_rl_223 ;
	7'h7f :
		TR_52 = RG_rl_223 ;
	default :
		TR_52 = 9'hx ;
	endcase
always @ ( RG_rl_224 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_53 = RG_rl_224 ;
	7'h01 :
		TR_53 = RG_rl_224 ;
	7'h02 :
		TR_53 = RG_rl_224 ;
	7'h03 :
		TR_53 = RG_rl_224 ;
	7'h04 :
		TR_53 = RG_rl_224 ;
	7'h05 :
		TR_53 = RG_rl_224 ;
	7'h06 :
		TR_53 = RG_rl_224 ;
	7'h07 :
		TR_53 = RG_rl_224 ;
	7'h08 :
		TR_53 = RG_rl_224 ;
	7'h09 :
		TR_53 = RG_rl_224 ;
	7'h0a :
		TR_53 = RG_rl_224 ;
	7'h0b :
		TR_53 = RG_rl_224 ;
	7'h0c :
		TR_53 = RG_rl_224 ;
	7'h0d :
		TR_53 = RG_rl_224 ;
	7'h0e :
		TR_53 = RG_rl_224 ;
	7'h0f :
		TR_53 = RG_rl_224 ;
	7'h10 :
		TR_53 = RG_rl_224 ;
	7'h11 :
		TR_53 = RG_rl_224 ;
	7'h12 :
		TR_53 = RG_rl_224 ;
	7'h13 :
		TR_53 = RG_rl_224 ;
	7'h14 :
		TR_53 = RG_rl_224 ;
	7'h15 :
		TR_53 = RG_rl_224 ;
	7'h16 :
		TR_53 = RG_rl_224 ;
	7'h17 :
		TR_53 = RG_rl_224 ;
	7'h18 :
		TR_53 = RG_rl_224 ;
	7'h19 :
		TR_53 = RG_rl_224 ;
	7'h1a :
		TR_53 = RG_rl_224 ;
	7'h1b :
		TR_53 = RG_rl_224 ;
	7'h1c :
		TR_53 = RG_rl_224 ;
	7'h1d :
		TR_53 = RG_rl_224 ;
	7'h1e :
		TR_53 = RG_rl_224 ;
	7'h1f :
		TR_53 = RG_rl_224 ;
	7'h20 :
		TR_53 = RG_rl_224 ;
	7'h21 :
		TR_53 = RG_rl_224 ;
	7'h22 :
		TR_53 = RG_rl_224 ;
	7'h23 :
		TR_53 = RG_rl_224 ;
	7'h24 :
		TR_53 = RG_rl_224 ;
	7'h25 :
		TR_53 = RG_rl_224 ;
	7'h26 :
		TR_53 = RG_rl_224 ;
	7'h27 :
		TR_53 = RG_rl_224 ;
	7'h28 :
		TR_53 = RG_rl_224 ;
	7'h29 :
		TR_53 = 9'h000 ;	// line#=../rle.cpp:68
	7'h2a :
		TR_53 = RG_rl_224 ;
	7'h2b :
		TR_53 = RG_rl_224 ;
	7'h2c :
		TR_53 = RG_rl_224 ;
	7'h2d :
		TR_53 = RG_rl_224 ;
	7'h2e :
		TR_53 = RG_rl_224 ;
	7'h2f :
		TR_53 = RG_rl_224 ;
	7'h30 :
		TR_53 = RG_rl_224 ;
	7'h31 :
		TR_53 = RG_rl_224 ;
	7'h32 :
		TR_53 = RG_rl_224 ;
	7'h33 :
		TR_53 = RG_rl_224 ;
	7'h34 :
		TR_53 = RG_rl_224 ;
	7'h35 :
		TR_53 = RG_rl_224 ;
	7'h36 :
		TR_53 = RG_rl_224 ;
	7'h37 :
		TR_53 = RG_rl_224 ;
	7'h38 :
		TR_53 = RG_rl_224 ;
	7'h39 :
		TR_53 = RG_rl_224 ;
	7'h3a :
		TR_53 = RG_rl_224 ;
	7'h3b :
		TR_53 = RG_rl_224 ;
	7'h3c :
		TR_53 = RG_rl_224 ;
	7'h3d :
		TR_53 = RG_rl_224 ;
	7'h3e :
		TR_53 = RG_rl_224 ;
	7'h3f :
		TR_53 = RG_rl_224 ;
	7'h40 :
		TR_53 = RG_rl_224 ;
	7'h41 :
		TR_53 = RG_rl_224 ;
	7'h42 :
		TR_53 = RG_rl_224 ;
	7'h43 :
		TR_53 = RG_rl_224 ;
	7'h44 :
		TR_53 = RG_rl_224 ;
	7'h45 :
		TR_53 = RG_rl_224 ;
	7'h46 :
		TR_53 = RG_rl_224 ;
	7'h47 :
		TR_53 = RG_rl_224 ;
	7'h48 :
		TR_53 = RG_rl_224 ;
	7'h49 :
		TR_53 = RG_rl_224 ;
	7'h4a :
		TR_53 = RG_rl_224 ;
	7'h4b :
		TR_53 = RG_rl_224 ;
	7'h4c :
		TR_53 = RG_rl_224 ;
	7'h4d :
		TR_53 = RG_rl_224 ;
	7'h4e :
		TR_53 = RG_rl_224 ;
	7'h4f :
		TR_53 = RG_rl_224 ;
	7'h50 :
		TR_53 = RG_rl_224 ;
	7'h51 :
		TR_53 = RG_rl_224 ;
	7'h52 :
		TR_53 = RG_rl_224 ;
	7'h53 :
		TR_53 = RG_rl_224 ;
	7'h54 :
		TR_53 = RG_rl_224 ;
	7'h55 :
		TR_53 = RG_rl_224 ;
	7'h56 :
		TR_53 = RG_rl_224 ;
	7'h57 :
		TR_53 = RG_rl_224 ;
	7'h58 :
		TR_53 = RG_rl_224 ;
	7'h59 :
		TR_53 = RG_rl_224 ;
	7'h5a :
		TR_53 = RG_rl_224 ;
	7'h5b :
		TR_53 = RG_rl_224 ;
	7'h5c :
		TR_53 = RG_rl_224 ;
	7'h5d :
		TR_53 = RG_rl_224 ;
	7'h5e :
		TR_53 = RG_rl_224 ;
	7'h5f :
		TR_53 = RG_rl_224 ;
	7'h60 :
		TR_53 = RG_rl_224 ;
	7'h61 :
		TR_53 = RG_rl_224 ;
	7'h62 :
		TR_53 = RG_rl_224 ;
	7'h63 :
		TR_53 = RG_rl_224 ;
	7'h64 :
		TR_53 = RG_rl_224 ;
	7'h65 :
		TR_53 = RG_rl_224 ;
	7'h66 :
		TR_53 = RG_rl_224 ;
	7'h67 :
		TR_53 = RG_rl_224 ;
	7'h68 :
		TR_53 = RG_rl_224 ;
	7'h69 :
		TR_53 = RG_rl_224 ;
	7'h6a :
		TR_53 = RG_rl_224 ;
	7'h6b :
		TR_53 = RG_rl_224 ;
	7'h6c :
		TR_53 = RG_rl_224 ;
	7'h6d :
		TR_53 = RG_rl_224 ;
	7'h6e :
		TR_53 = RG_rl_224 ;
	7'h6f :
		TR_53 = RG_rl_224 ;
	7'h70 :
		TR_53 = RG_rl_224 ;
	7'h71 :
		TR_53 = RG_rl_224 ;
	7'h72 :
		TR_53 = RG_rl_224 ;
	7'h73 :
		TR_53 = RG_rl_224 ;
	7'h74 :
		TR_53 = RG_rl_224 ;
	7'h75 :
		TR_53 = RG_rl_224 ;
	7'h76 :
		TR_53 = RG_rl_224 ;
	7'h77 :
		TR_53 = RG_rl_224 ;
	7'h78 :
		TR_53 = RG_rl_224 ;
	7'h79 :
		TR_53 = RG_rl_224 ;
	7'h7a :
		TR_53 = RG_rl_224 ;
	7'h7b :
		TR_53 = RG_rl_224 ;
	7'h7c :
		TR_53 = RG_rl_224 ;
	7'h7d :
		TR_53 = RG_rl_224 ;
	7'h7e :
		TR_53 = RG_rl_224 ;
	7'h7f :
		TR_53 = RG_rl_224 ;
	default :
		TR_53 = 9'hx ;
	endcase
always @ ( RG_rl_225 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_54 = RG_rl_225 ;
	7'h01 :
		TR_54 = RG_rl_225 ;
	7'h02 :
		TR_54 = RG_rl_225 ;
	7'h03 :
		TR_54 = RG_rl_225 ;
	7'h04 :
		TR_54 = RG_rl_225 ;
	7'h05 :
		TR_54 = RG_rl_225 ;
	7'h06 :
		TR_54 = RG_rl_225 ;
	7'h07 :
		TR_54 = RG_rl_225 ;
	7'h08 :
		TR_54 = RG_rl_225 ;
	7'h09 :
		TR_54 = RG_rl_225 ;
	7'h0a :
		TR_54 = RG_rl_225 ;
	7'h0b :
		TR_54 = RG_rl_225 ;
	7'h0c :
		TR_54 = RG_rl_225 ;
	7'h0d :
		TR_54 = RG_rl_225 ;
	7'h0e :
		TR_54 = RG_rl_225 ;
	7'h0f :
		TR_54 = RG_rl_225 ;
	7'h10 :
		TR_54 = RG_rl_225 ;
	7'h11 :
		TR_54 = RG_rl_225 ;
	7'h12 :
		TR_54 = RG_rl_225 ;
	7'h13 :
		TR_54 = RG_rl_225 ;
	7'h14 :
		TR_54 = RG_rl_225 ;
	7'h15 :
		TR_54 = RG_rl_225 ;
	7'h16 :
		TR_54 = RG_rl_225 ;
	7'h17 :
		TR_54 = RG_rl_225 ;
	7'h18 :
		TR_54 = RG_rl_225 ;
	7'h19 :
		TR_54 = RG_rl_225 ;
	7'h1a :
		TR_54 = RG_rl_225 ;
	7'h1b :
		TR_54 = RG_rl_225 ;
	7'h1c :
		TR_54 = RG_rl_225 ;
	7'h1d :
		TR_54 = RG_rl_225 ;
	7'h1e :
		TR_54 = RG_rl_225 ;
	7'h1f :
		TR_54 = RG_rl_225 ;
	7'h20 :
		TR_54 = RG_rl_225 ;
	7'h21 :
		TR_54 = RG_rl_225 ;
	7'h22 :
		TR_54 = RG_rl_225 ;
	7'h23 :
		TR_54 = RG_rl_225 ;
	7'h24 :
		TR_54 = RG_rl_225 ;
	7'h25 :
		TR_54 = RG_rl_225 ;
	7'h26 :
		TR_54 = RG_rl_225 ;
	7'h27 :
		TR_54 = RG_rl_225 ;
	7'h28 :
		TR_54 = RG_rl_225 ;
	7'h29 :
		TR_54 = RG_rl_225 ;
	7'h2a :
		TR_54 = 9'h000 ;	// line#=../rle.cpp:68
	7'h2b :
		TR_54 = RG_rl_225 ;
	7'h2c :
		TR_54 = RG_rl_225 ;
	7'h2d :
		TR_54 = RG_rl_225 ;
	7'h2e :
		TR_54 = RG_rl_225 ;
	7'h2f :
		TR_54 = RG_rl_225 ;
	7'h30 :
		TR_54 = RG_rl_225 ;
	7'h31 :
		TR_54 = RG_rl_225 ;
	7'h32 :
		TR_54 = RG_rl_225 ;
	7'h33 :
		TR_54 = RG_rl_225 ;
	7'h34 :
		TR_54 = RG_rl_225 ;
	7'h35 :
		TR_54 = RG_rl_225 ;
	7'h36 :
		TR_54 = RG_rl_225 ;
	7'h37 :
		TR_54 = RG_rl_225 ;
	7'h38 :
		TR_54 = RG_rl_225 ;
	7'h39 :
		TR_54 = RG_rl_225 ;
	7'h3a :
		TR_54 = RG_rl_225 ;
	7'h3b :
		TR_54 = RG_rl_225 ;
	7'h3c :
		TR_54 = RG_rl_225 ;
	7'h3d :
		TR_54 = RG_rl_225 ;
	7'h3e :
		TR_54 = RG_rl_225 ;
	7'h3f :
		TR_54 = RG_rl_225 ;
	7'h40 :
		TR_54 = RG_rl_225 ;
	7'h41 :
		TR_54 = RG_rl_225 ;
	7'h42 :
		TR_54 = RG_rl_225 ;
	7'h43 :
		TR_54 = RG_rl_225 ;
	7'h44 :
		TR_54 = RG_rl_225 ;
	7'h45 :
		TR_54 = RG_rl_225 ;
	7'h46 :
		TR_54 = RG_rl_225 ;
	7'h47 :
		TR_54 = RG_rl_225 ;
	7'h48 :
		TR_54 = RG_rl_225 ;
	7'h49 :
		TR_54 = RG_rl_225 ;
	7'h4a :
		TR_54 = RG_rl_225 ;
	7'h4b :
		TR_54 = RG_rl_225 ;
	7'h4c :
		TR_54 = RG_rl_225 ;
	7'h4d :
		TR_54 = RG_rl_225 ;
	7'h4e :
		TR_54 = RG_rl_225 ;
	7'h4f :
		TR_54 = RG_rl_225 ;
	7'h50 :
		TR_54 = RG_rl_225 ;
	7'h51 :
		TR_54 = RG_rl_225 ;
	7'h52 :
		TR_54 = RG_rl_225 ;
	7'h53 :
		TR_54 = RG_rl_225 ;
	7'h54 :
		TR_54 = RG_rl_225 ;
	7'h55 :
		TR_54 = RG_rl_225 ;
	7'h56 :
		TR_54 = RG_rl_225 ;
	7'h57 :
		TR_54 = RG_rl_225 ;
	7'h58 :
		TR_54 = RG_rl_225 ;
	7'h59 :
		TR_54 = RG_rl_225 ;
	7'h5a :
		TR_54 = RG_rl_225 ;
	7'h5b :
		TR_54 = RG_rl_225 ;
	7'h5c :
		TR_54 = RG_rl_225 ;
	7'h5d :
		TR_54 = RG_rl_225 ;
	7'h5e :
		TR_54 = RG_rl_225 ;
	7'h5f :
		TR_54 = RG_rl_225 ;
	7'h60 :
		TR_54 = RG_rl_225 ;
	7'h61 :
		TR_54 = RG_rl_225 ;
	7'h62 :
		TR_54 = RG_rl_225 ;
	7'h63 :
		TR_54 = RG_rl_225 ;
	7'h64 :
		TR_54 = RG_rl_225 ;
	7'h65 :
		TR_54 = RG_rl_225 ;
	7'h66 :
		TR_54 = RG_rl_225 ;
	7'h67 :
		TR_54 = RG_rl_225 ;
	7'h68 :
		TR_54 = RG_rl_225 ;
	7'h69 :
		TR_54 = RG_rl_225 ;
	7'h6a :
		TR_54 = RG_rl_225 ;
	7'h6b :
		TR_54 = RG_rl_225 ;
	7'h6c :
		TR_54 = RG_rl_225 ;
	7'h6d :
		TR_54 = RG_rl_225 ;
	7'h6e :
		TR_54 = RG_rl_225 ;
	7'h6f :
		TR_54 = RG_rl_225 ;
	7'h70 :
		TR_54 = RG_rl_225 ;
	7'h71 :
		TR_54 = RG_rl_225 ;
	7'h72 :
		TR_54 = RG_rl_225 ;
	7'h73 :
		TR_54 = RG_rl_225 ;
	7'h74 :
		TR_54 = RG_rl_225 ;
	7'h75 :
		TR_54 = RG_rl_225 ;
	7'h76 :
		TR_54 = RG_rl_225 ;
	7'h77 :
		TR_54 = RG_rl_225 ;
	7'h78 :
		TR_54 = RG_rl_225 ;
	7'h79 :
		TR_54 = RG_rl_225 ;
	7'h7a :
		TR_54 = RG_rl_225 ;
	7'h7b :
		TR_54 = RG_rl_225 ;
	7'h7c :
		TR_54 = RG_rl_225 ;
	7'h7d :
		TR_54 = RG_rl_225 ;
	7'h7e :
		TR_54 = RG_rl_225 ;
	7'h7f :
		TR_54 = RG_rl_225 ;
	default :
		TR_54 = 9'hx ;
	endcase
always @ ( RG_rl_226 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_55 = RG_rl_226 ;
	7'h01 :
		TR_55 = RG_rl_226 ;
	7'h02 :
		TR_55 = RG_rl_226 ;
	7'h03 :
		TR_55 = RG_rl_226 ;
	7'h04 :
		TR_55 = RG_rl_226 ;
	7'h05 :
		TR_55 = RG_rl_226 ;
	7'h06 :
		TR_55 = RG_rl_226 ;
	7'h07 :
		TR_55 = RG_rl_226 ;
	7'h08 :
		TR_55 = RG_rl_226 ;
	7'h09 :
		TR_55 = RG_rl_226 ;
	7'h0a :
		TR_55 = RG_rl_226 ;
	7'h0b :
		TR_55 = RG_rl_226 ;
	7'h0c :
		TR_55 = RG_rl_226 ;
	7'h0d :
		TR_55 = RG_rl_226 ;
	7'h0e :
		TR_55 = RG_rl_226 ;
	7'h0f :
		TR_55 = RG_rl_226 ;
	7'h10 :
		TR_55 = RG_rl_226 ;
	7'h11 :
		TR_55 = RG_rl_226 ;
	7'h12 :
		TR_55 = RG_rl_226 ;
	7'h13 :
		TR_55 = RG_rl_226 ;
	7'h14 :
		TR_55 = RG_rl_226 ;
	7'h15 :
		TR_55 = RG_rl_226 ;
	7'h16 :
		TR_55 = RG_rl_226 ;
	7'h17 :
		TR_55 = RG_rl_226 ;
	7'h18 :
		TR_55 = RG_rl_226 ;
	7'h19 :
		TR_55 = RG_rl_226 ;
	7'h1a :
		TR_55 = RG_rl_226 ;
	7'h1b :
		TR_55 = RG_rl_226 ;
	7'h1c :
		TR_55 = RG_rl_226 ;
	7'h1d :
		TR_55 = RG_rl_226 ;
	7'h1e :
		TR_55 = RG_rl_226 ;
	7'h1f :
		TR_55 = RG_rl_226 ;
	7'h20 :
		TR_55 = RG_rl_226 ;
	7'h21 :
		TR_55 = RG_rl_226 ;
	7'h22 :
		TR_55 = RG_rl_226 ;
	7'h23 :
		TR_55 = RG_rl_226 ;
	7'h24 :
		TR_55 = RG_rl_226 ;
	7'h25 :
		TR_55 = RG_rl_226 ;
	7'h26 :
		TR_55 = RG_rl_226 ;
	7'h27 :
		TR_55 = RG_rl_226 ;
	7'h28 :
		TR_55 = RG_rl_226 ;
	7'h29 :
		TR_55 = RG_rl_226 ;
	7'h2a :
		TR_55 = RG_rl_226 ;
	7'h2b :
		TR_55 = 9'h000 ;	// line#=../rle.cpp:68
	7'h2c :
		TR_55 = RG_rl_226 ;
	7'h2d :
		TR_55 = RG_rl_226 ;
	7'h2e :
		TR_55 = RG_rl_226 ;
	7'h2f :
		TR_55 = RG_rl_226 ;
	7'h30 :
		TR_55 = RG_rl_226 ;
	7'h31 :
		TR_55 = RG_rl_226 ;
	7'h32 :
		TR_55 = RG_rl_226 ;
	7'h33 :
		TR_55 = RG_rl_226 ;
	7'h34 :
		TR_55 = RG_rl_226 ;
	7'h35 :
		TR_55 = RG_rl_226 ;
	7'h36 :
		TR_55 = RG_rl_226 ;
	7'h37 :
		TR_55 = RG_rl_226 ;
	7'h38 :
		TR_55 = RG_rl_226 ;
	7'h39 :
		TR_55 = RG_rl_226 ;
	7'h3a :
		TR_55 = RG_rl_226 ;
	7'h3b :
		TR_55 = RG_rl_226 ;
	7'h3c :
		TR_55 = RG_rl_226 ;
	7'h3d :
		TR_55 = RG_rl_226 ;
	7'h3e :
		TR_55 = RG_rl_226 ;
	7'h3f :
		TR_55 = RG_rl_226 ;
	7'h40 :
		TR_55 = RG_rl_226 ;
	7'h41 :
		TR_55 = RG_rl_226 ;
	7'h42 :
		TR_55 = RG_rl_226 ;
	7'h43 :
		TR_55 = RG_rl_226 ;
	7'h44 :
		TR_55 = RG_rl_226 ;
	7'h45 :
		TR_55 = RG_rl_226 ;
	7'h46 :
		TR_55 = RG_rl_226 ;
	7'h47 :
		TR_55 = RG_rl_226 ;
	7'h48 :
		TR_55 = RG_rl_226 ;
	7'h49 :
		TR_55 = RG_rl_226 ;
	7'h4a :
		TR_55 = RG_rl_226 ;
	7'h4b :
		TR_55 = RG_rl_226 ;
	7'h4c :
		TR_55 = RG_rl_226 ;
	7'h4d :
		TR_55 = RG_rl_226 ;
	7'h4e :
		TR_55 = RG_rl_226 ;
	7'h4f :
		TR_55 = RG_rl_226 ;
	7'h50 :
		TR_55 = RG_rl_226 ;
	7'h51 :
		TR_55 = RG_rl_226 ;
	7'h52 :
		TR_55 = RG_rl_226 ;
	7'h53 :
		TR_55 = RG_rl_226 ;
	7'h54 :
		TR_55 = RG_rl_226 ;
	7'h55 :
		TR_55 = RG_rl_226 ;
	7'h56 :
		TR_55 = RG_rl_226 ;
	7'h57 :
		TR_55 = RG_rl_226 ;
	7'h58 :
		TR_55 = RG_rl_226 ;
	7'h59 :
		TR_55 = RG_rl_226 ;
	7'h5a :
		TR_55 = RG_rl_226 ;
	7'h5b :
		TR_55 = RG_rl_226 ;
	7'h5c :
		TR_55 = RG_rl_226 ;
	7'h5d :
		TR_55 = RG_rl_226 ;
	7'h5e :
		TR_55 = RG_rl_226 ;
	7'h5f :
		TR_55 = RG_rl_226 ;
	7'h60 :
		TR_55 = RG_rl_226 ;
	7'h61 :
		TR_55 = RG_rl_226 ;
	7'h62 :
		TR_55 = RG_rl_226 ;
	7'h63 :
		TR_55 = RG_rl_226 ;
	7'h64 :
		TR_55 = RG_rl_226 ;
	7'h65 :
		TR_55 = RG_rl_226 ;
	7'h66 :
		TR_55 = RG_rl_226 ;
	7'h67 :
		TR_55 = RG_rl_226 ;
	7'h68 :
		TR_55 = RG_rl_226 ;
	7'h69 :
		TR_55 = RG_rl_226 ;
	7'h6a :
		TR_55 = RG_rl_226 ;
	7'h6b :
		TR_55 = RG_rl_226 ;
	7'h6c :
		TR_55 = RG_rl_226 ;
	7'h6d :
		TR_55 = RG_rl_226 ;
	7'h6e :
		TR_55 = RG_rl_226 ;
	7'h6f :
		TR_55 = RG_rl_226 ;
	7'h70 :
		TR_55 = RG_rl_226 ;
	7'h71 :
		TR_55 = RG_rl_226 ;
	7'h72 :
		TR_55 = RG_rl_226 ;
	7'h73 :
		TR_55 = RG_rl_226 ;
	7'h74 :
		TR_55 = RG_rl_226 ;
	7'h75 :
		TR_55 = RG_rl_226 ;
	7'h76 :
		TR_55 = RG_rl_226 ;
	7'h77 :
		TR_55 = RG_rl_226 ;
	7'h78 :
		TR_55 = RG_rl_226 ;
	7'h79 :
		TR_55 = RG_rl_226 ;
	7'h7a :
		TR_55 = RG_rl_226 ;
	7'h7b :
		TR_55 = RG_rl_226 ;
	7'h7c :
		TR_55 = RG_rl_226 ;
	7'h7d :
		TR_55 = RG_rl_226 ;
	7'h7e :
		TR_55 = RG_rl_226 ;
	7'h7f :
		TR_55 = RG_rl_226 ;
	default :
		TR_55 = 9'hx ;
	endcase
always @ ( RG_rl_227 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_56 = RG_rl_227 ;
	7'h01 :
		TR_56 = RG_rl_227 ;
	7'h02 :
		TR_56 = RG_rl_227 ;
	7'h03 :
		TR_56 = RG_rl_227 ;
	7'h04 :
		TR_56 = RG_rl_227 ;
	7'h05 :
		TR_56 = RG_rl_227 ;
	7'h06 :
		TR_56 = RG_rl_227 ;
	7'h07 :
		TR_56 = RG_rl_227 ;
	7'h08 :
		TR_56 = RG_rl_227 ;
	7'h09 :
		TR_56 = RG_rl_227 ;
	7'h0a :
		TR_56 = RG_rl_227 ;
	7'h0b :
		TR_56 = RG_rl_227 ;
	7'h0c :
		TR_56 = RG_rl_227 ;
	7'h0d :
		TR_56 = RG_rl_227 ;
	7'h0e :
		TR_56 = RG_rl_227 ;
	7'h0f :
		TR_56 = RG_rl_227 ;
	7'h10 :
		TR_56 = RG_rl_227 ;
	7'h11 :
		TR_56 = RG_rl_227 ;
	7'h12 :
		TR_56 = RG_rl_227 ;
	7'h13 :
		TR_56 = RG_rl_227 ;
	7'h14 :
		TR_56 = RG_rl_227 ;
	7'h15 :
		TR_56 = RG_rl_227 ;
	7'h16 :
		TR_56 = RG_rl_227 ;
	7'h17 :
		TR_56 = RG_rl_227 ;
	7'h18 :
		TR_56 = RG_rl_227 ;
	7'h19 :
		TR_56 = RG_rl_227 ;
	7'h1a :
		TR_56 = RG_rl_227 ;
	7'h1b :
		TR_56 = RG_rl_227 ;
	7'h1c :
		TR_56 = RG_rl_227 ;
	7'h1d :
		TR_56 = RG_rl_227 ;
	7'h1e :
		TR_56 = RG_rl_227 ;
	7'h1f :
		TR_56 = RG_rl_227 ;
	7'h20 :
		TR_56 = RG_rl_227 ;
	7'h21 :
		TR_56 = RG_rl_227 ;
	7'h22 :
		TR_56 = RG_rl_227 ;
	7'h23 :
		TR_56 = RG_rl_227 ;
	7'h24 :
		TR_56 = RG_rl_227 ;
	7'h25 :
		TR_56 = RG_rl_227 ;
	7'h26 :
		TR_56 = RG_rl_227 ;
	7'h27 :
		TR_56 = RG_rl_227 ;
	7'h28 :
		TR_56 = RG_rl_227 ;
	7'h29 :
		TR_56 = RG_rl_227 ;
	7'h2a :
		TR_56 = RG_rl_227 ;
	7'h2b :
		TR_56 = RG_rl_227 ;
	7'h2c :
		TR_56 = 9'h000 ;	// line#=../rle.cpp:68
	7'h2d :
		TR_56 = RG_rl_227 ;
	7'h2e :
		TR_56 = RG_rl_227 ;
	7'h2f :
		TR_56 = RG_rl_227 ;
	7'h30 :
		TR_56 = RG_rl_227 ;
	7'h31 :
		TR_56 = RG_rl_227 ;
	7'h32 :
		TR_56 = RG_rl_227 ;
	7'h33 :
		TR_56 = RG_rl_227 ;
	7'h34 :
		TR_56 = RG_rl_227 ;
	7'h35 :
		TR_56 = RG_rl_227 ;
	7'h36 :
		TR_56 = RG_rl_227 ;
	7'h37 :
		TR_56 = RG_rl_227 ;
	7'h38 :
		TR_56 = RG_rl_227 ;
	7'h39 :
		TR_56 = RG_rl_227 ;
	7'h3a :
		TR_56 = RG_rl_227 ;
	7'h3b :
		TR_56 = RG_rl_227 ;
	7'h3c :
		TR_56 = RG_rl_227 ;
	7'h3d :
		TR_56 = RG_rl_227 ;
	7'h3e :
		TR_56 = RG_rl_227 ;
	7'h3f :
		TR_56 = RG_rl_227 ;
	7'h40 :
		TR_56 = RG_rl_227 ;
	7'h41 :
		TR_56 = RG_rl_227 ;
	7'h42 :
		TR_56 = RG_rl_227 ;
	7'h43 :
		TR_56 = RG_rl_227 ;
	7'h44 :
		TR_56 = RG_rl_227 ;
	7'h45 :
		TR_56 = RG_rl_227 ;
	7'h46 :
		TR_56 = RG_rl_227 ;
	7'h47 :
		TR_56 = RG_rl_227 ;
	7'h48 :
		TR_56 = RG_rl_227 ;
	7'h49 :
		TR_56 = RG_rl_227 ;
	7'h4a :
		TR_56 = RG_rl_227 ;
	7'h4b :
		TR_56 = RG_rl_227 ;
	7'h4c :
		TR_56 = RG_rl_227 ;
	7'h4d :
		TR_56 = RG_rl_227 ;
	7'h4e :
		TR_56 = RG_rl_227 ;
	7'h4f :
		TR_56 = RG_rl_227 ;
	7'h50 :
		TR_56 = RG_rl_227 ;
	7'h51 :
		TR_56 = RG_rl_227 ;
	7'h52 :
		TR_56 = RG_rl_227 ;
	7'h53 :
		TR_56 = RG_rl_227 ;
	7'h54 :
		TR_56 = RG_rl_227 ;
	7'h55 :
		TR_56 = RG_rl_227 ;
	7'h56 :
		TR_56 = RG_rl_227 ;
	7'h57 :
		TR_56 = RG_rl_227 ;
	7'h58 :
		TR_56 = RG_rl_227 ;
	7'h59 :
		TR_56 = RG_rl_227 ;
	7'h5a :
		TR_56 = RG_rl_227 ;
	7'h5b :
		TR_56 = RG_rl_227 ;
	7'h5c :
		TR_56 = RG_rl_227 ;
	7'h5d :
		TR_56 = RG_rl_227 ;
	7'h5e :
		TR_56 = RG_rl_227 ;
	7'h5f :
		TR_56 = RG_rl_227 ;
	7'h60 :
		TR_56 = RG_rl_227 ;
	7'h61 :
		TR_56 = RG_rl_227 ;
	7'h62 :
		TR_56 = RG_rl_227 ;
	7'h63 :
		TR_56 = RG_rl_227 ;
	7'h64 :
		TR_56 = RG_rl_227 ;
	7'h65 :
		TR_56 = RG_rl_227 ;
	7'h66 :
		TR_56 = RG_rl_227 ;
	7'h67 :
		TR_56 = RG_rl_227 ;
	7'h68 :
		TR_56 = RG_rl_227 ;
	7'h69 :
		TR_56 = RG_rl_227 ;
	7'h6a :
		TR_56 = RG_rl_227 ;
	7'h6b :
		TR_56 = RG_rl_227 ;
	7'h6c :
		TR_56 = RG_rl_227 ;
	7'h6d :
		TR_56 = RG_rl_227 ;
	7'h6e :
		TR_56 = RG_rl_227 ;
	7'h6f :
		TR_56 = RG_rl_227 ;
	7'h70 :
		TR_56 = RG_rl_227 ;
	7'h71 :
		TR_56 = RG_rl_227 ;
	7'h72 :
		TR_56 = RG_rl_227 ;
	7'h73 :
		TR_56 = RG_rl_227 ;
	7'h74 :
		TR_56 = RG_rl_227 ;
	7'h75 :
		TR_56 = RG_rl_227 ;
	7'h76 :
		TR_56 = RG_rl_227 ;
	7'h77 :
		TR_56 = RG_rl_227 ;
	7'h78 :
		TR_56 = RG_rl_227 ;
	7'h79 :
		TR_56 = RG_rl_227 ;
	7'h7a :
		TR_56 = RG_rl_227 ;
	7'h7b :
		TR_56 = RG_rl_227 ;
	7'h7c :
		TR_56 = RG_rl_227 ;
	7'h7d :
		TR_56 = RG_rl_227 ;
	7'h7e :
		TR_56 = RG_rl_227 ;
	7'h7f :
		TR_56 = RG_rl_227 ;
	default :
		TR_56 = 9'hx ;
	endcase
always @ ( RG_rl_228 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_57 = RG_rl_228 ;
	7'h01 :
		TR_57 = RG_rl_228 ;
	7'h02 :
		TR_57 = RG_rl_228 ;
	7'h03 :
		TR_57 = RG_rl_228 ;
	7'h04 :
		TR_57 = RG_rl_228 ;
	7'h05 :
		TR_57 = RG_rl_228 ;
	7'h06 :
		TR_57 = RG_rl_228 ;
	7'h07 :
		TR_57 = RG_rl_228 ;
	7'h08 :
		TR_57 = RG_rl_228 ;
	7'h09 :
		TR_57 = RG_rl_228 ;
	7'h0a :
		TR_57 = RG_rl_228 ;
	7'h0b :
		TR_57 = RG_rl_228 ;
	7'h0c :
		TR_57 = RG_rl_228 ;
	7'h0d :
		TR_57 = RG_rl_228 ;
	7'h0e :
		TR_57 = RG_rl_228 ;
	7'h0f :
		TR_57 = RG_rl_228 ;
	7'h10 :
		TR_57 = RG_rl_228 ;
	7'h11 :
		TR_57 = RG_rl_228 ;
	7'h12 :
		TR_57 = RG_rl_228 ;
	7'h13 :
		TR_57 = RG_rl_228 ;
	7'h14 :
		TR_57 = RG_rl_228 ;
	7'h15 :
		TR_57 = RG_rl_228 ;
	7'h16 :
		TR_57 = RG_rl_228 ;
	7'h17 :
		TR_57 = RG_rl_228 ;
	7'h18 :
		TR_57 = RG_rl_228 ;
	7'h19 :
		TR_57 = RG_rl_228 ;
	7'h1a :
		TR_57 = RG_rl_228 ;
	7'h1b :
		TR_57 = RG_rl_228 ;
	7'h1c :
		TR_57 = RG_rl_228 ;
	7'h1d :
		TR_57 = RG_rl_228 ;
	7'h1e :
		TR_57 = RG_rl_228 ;
	7'h1f :
		TR_57 = RG_rl_228 ;
	7'h20 :
		TR_57 = RG_rl_228 ;
	7'h21 :
		TR_57 = RG_rl_228 ;
	7'h22 :
		TR_57 = RG_rl_228 ;
	7'h23 :
		TR_57 = RG_rl_228 ;
	7'h24 :
		TR_57 = RG_rl_228 ;
	7'h25 :
		TR_57 = RG_rl_228 ;
	7'h26 :
		TR_57 = RG_rl_228 ;
	7'h27 :
		TR_57 = RG_rl_228 ;
	7'h28 :
		TR_57 = RG_rl_228 ;
	7'h29 :
		TR_57 = RG_rl_228 ;
	7'h2a :
		TR_57 = RG_rl_228 ;
	7'h2b :
		TR_57 = RG_rl_228 ;
	7'h2c :
		TR_57 = RG_rl_228 ;
	7'h2d :
		TR_57 = 9'h000 ;	// line#=../rle.cpp:68
	7'h2e :
		TR_57 = RG_rl_228 ;
	7'h2f :
		TR_57 = RG_rl_228 ;
	7'h30 :
		TR_57 = RG_rl_228 ;
	7'h31 :
		TR_57 = RG_rl_228 ;
	7'h32 :
		TR_57 = RG_rl_228 ;
	7'h33 :
		TR_57 = RG_rl_228 ;
	7'h34 :
		TR_57 = RG_rl_228 ;
	7'h35 :
		TR_57 = RG_rl_228 ;
	7'h36 :
		TR_57 = RG_rl_228 ;
	7'h37 :
		TR_57 = RG_rl_228 ;
	7'h38 :
		TR_57 = RG_rl_228 ;
	7'h39 :
		TR_57 = RG_rl_228 ;
	7'h3a :
		TR_57 = RG_rl_228 ;
	7'h3b :
		TR_57 = RG_rl_228 ;
	7'h3c :
		TR_57 = RG_rl_228 ;
	7'h3d :
		TR_57 = RG_rl_228 ;
	7'h3e :
		TR_57 = RG_rl_228 ;
	7'h3f :
		TR_57 = RG_rl_228 ;
	7'h40 :
		TR_57 = RG_rl_228 ;
	7'h41 :
		TR_57 = RG_rl_228 ;
	7'h42 :
		TR_57 = RG_rl_228 ;
	7'h43 :
		TR_57 = RG_rl_228 ;
	7'h44 :
		TR_57 = RG_rl_228 ;
	7'h45 :
		TR_57 = RG_rl_228 ;
	7'h46 :
		TR_57 = RG_rl_228 ;
	7'h47 :
		TR_57 = RG_rl_228 ;
	7'h48 :
		TR_57 = RG_rl_228 ;
	7'h49 :
		TR_57 = RG_rl_228 ;
	7'h4a :
		TR_57 = RG_rl_228 ;
	7'h4b :
		TR_57 = RG_rl_228 ;
	7'h4c :
		TR_57 = RG_rl_228 ;
	7'h4d :
		TR_57 = RG_rl_228 ;
	7'h4e :
		TR_57 = RG_rl_228 ;
	7'h4f :
		TR_57 = RG_rl_228 ;
	7'h50 :
		TR_57 = RG_rl_228 ;
	7'h51 :
		TR_57 = RG_rl_228 ;
	7'h52 :
		TR_57 = RG_rl_228 ;
	7'h53 :
		TR_57 = RG_rl_228 ;
	7'h54 :
		TR_57 = RG_rl_228 ;
	7'h55 :
		TR_57 = RG_rl_228 ;
	7'h56 :
		TR_57 = RG_rl_228 ;
	7'h57 :
		TR_57 = RG_rl_228 ;
	7'h58 :
		TR_57 = RG_rl_228 ;
	7'h59 :
		TR_57 = RG_rl_228 ;
	7'h5a :
		TR_57 = RG_rl_228 ;
	7'h5b :
		TR_57 = RG_rl_228 ;
	7'h5c :
		TR_57 = RG_rl_228 ;
	7'h5d :
		TR_57 = RG_rl_228 ;
	7'h5e :
		TR_57 = RG_rl_228 ;
	7'h5f :
		TR_57 = RG_rl_228 ;
	7'h60 :
		TR_57 = RG_rl_228 ;
	7'h61 :
		TR_57 = RG_rl_228 ;
	7'h62 :
		TR_57 = RG_rl_228 ;
	7'h63 :
		TR_57 = RG_rl_228 ;
	7'h64 :
		TR_57 = RG_rl_228 ;
	7'h65 :
		TR_57 = RG_rl_228 ;
	7'h66 :
		TR_57 = RG_rl_228 ;
	7'h67 :
		TR_57 = RG_rl_228 ;
	7'h68 :
		TR_57 = RG_rl_228 ;
	7'h69 :
		TR_57 = RG_rl_228 ;
	7'h6a :
		TR_57 = RG_rl_228 ;
	7'h6b :
		TR_57 = RG_rl_228 ;
	7'h6c :
		TR_57 = RG_rl_228 ;
	7'h6d :
		TR_57 = RG_rl_228 ;
	7'h6e :
		TR_57 = RG_rl_228 ;
	7'h6f :
		TR_57 = RG_rl_228 ;
	7'h70 :
		TR_57 = RG_rl_228 ;
	7'h71 :
		TR_57 = RG_rl_228 ;
	7'h72 :
		TR_57 = RG_rl_228 ;
	7'h73 :
		TR_57 = RG_rl_228 ;
	7'h74 :
		TR_57 = RG_rl_228 ;
	7'h75 :
		TR_57 = RG_rl_228 ;
	7'h76 :
		TR_57 = RG_rl_228 ;
	7'h77 :
		TR_57 = RG_rl_228 ;
	7'h78 :
		TR_57 = RG_rl_228 ;
	7'h79 :
		TR_57 = RG_rl_228 ;
	7'h7a :
		TR_57 = RG_rl_228 ;
	7'h7b :
		TR_57 = RG_rl_228 ;
	7'h7c :
		TR_57 = RG_rl_228 ;
	7'h7d :
		TR_57 = RG_rl_228 ;
	7'h7e :
		TR_57 = RG_rl_228 ;
	7'h7f :
		TR_57 = RG_rl_228 ;
	default :
		TR_57 = 9'hx ;
	endcase
always @ ( RG_rl_229 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_58 = RG_rl_229 ;
	7'h01 :
		TR_58 = RG_rl_229 ;
	7'h02 :
		TR_58 = RG_rl_229 ;
	7'h03 :
		TR_58 = RG_rl_229 ;
	7'h04 :
		TR_58 = RG_rl_229 ;
	7'h05 :
		TR_58 = RG_rl_229 ;
	7'h06 :
		TR_58 = RG_rl_229 ;
	7'h07 :
		TR_58 = RG_rl_229 ;
	7'h08 :
		TR_58 = RG_rl_229 ;
	7'h09 :
		TR_58 = RG_rl_229 ;
	7'h0a :
		TR_58 = RG_rl_229 ;
	7'h0b :
		TR_58 = RG_rl_229 ;
	7'h0c :
		TR_58 = RG_rl_229 ;
	7'h0d :
		TR_58 = RG_rl_229 ;
	7'h0e :
		TR_58 = RG_rl_229 ;
	7'h0f :
		TR_58 = RG_rl_229 ;
	7'h10 :
		TR_58 = RG_rl_229 ;
	7'h11 :
		TR_58 = RG_rl_229 ;
	7'h12 :
		TR_58 = RG_rl_229 ;
	7'h13 :
		TR_58 = RG_rl_229 ;
	7'h14 :
		TR_58 = RG_rl_229 ;
	7'h15 :
		TR_58 = RG_rl_229 ;
	7'h16 :
		TR_58 = RG_rl_229 ;
	7'h17 :
		TR_58 = RG_rl_229 ;
	7'h18 :
		TR_58 = RG_rl_229 ;
	7'h19 :
		TR_58 = RG_rl_229 ;
	7'h1a :
		TR_58 = RG_rl_229 ;
	7'h1b :
		TR_58 = RG_rl_229 ;
	7'h1c :
		TR_58 = RG_rl_229 ;
	7'h1d :
		TR_58 = RG_rl_229 ;
	7'h1e :
		TR_58 = RG_rl_229 ;
	7'h1f :
		TR_58 = RG_rl_229 ;
	7'h20 :
		TR_58 = RG_rl_229 ;
	7'h21 :
		TR_58 = RG_rl_229 ;
	7'h22 :
		TR_58 = RG_rl_229 ;
	7'h23 :
		TR_58 = RG_rl_229 ;
	7'h24 :
		TR_58 = RG_rl_229 ;
	7'h25 :
		TR_58 = RG_rl_229 ;
	7'h26 :
		TR_58 = RG_rl_229 ;
	7'h27 :
		TR_58 = RG_rl_229 ;
	7'h28 :
		TR_58 = RG_rl_229 ;
	7'h29 :
		TR_58 = RG_rl_229 ;
	7'h2a :
		TR_58 = RG_rl_229 ;
	7'h2b :
		TR_58 = RG_rl_229 ;
	7'h2c :
		TR_58 = RG_rl_229 ;
	7'h2d :
		TR_58 = RG_rl_229 ;
	7'h2e :
		TR_58 = 9'h000 ;	// line#=../rle.cpp:68
	7'h2f :
		TR_58 = RG_rl_229 ;
	7'h30 :
		TR_58 = RG_rl_229 ;
	7'h31 :
		TR_58 = RG_rl_229 ;
	7'h32 :
		TR_58 = RG_rl_229 ;
	7'h33 :
		TR_58 = RG_rl_229 ;
	7'h34 :
		TR_58 = RG_rl_229 ;
	7'h35 :
		TR_58 = RG_rl_229 ;
	7'h36 :
		TR_58 = RG_rl_229 ;
	7'h37 :
		TR_58 = RG_rl_229 ;
	7'h38 :
		TR_58 = RG_rl_229 ;
	7'h39 :
		TR_58 = RG_rl_229 ;
	7'h3a :
		TR_58 = RG_rl_229 ;
	7'h3b :
		TR_58 = RG_rl_229 ;
	7'h3c :
		TR_58 = RG_rl_229 ;
	7'h3d :
		TR_58 = RG_rl_229 ;
	7'h3e :
		TR_58 = RG_rl_229 ;
	7'h3f :
		TR_58 = RG_rl_229 ;
	7'h40 :
		TR_58 = RG_rl_229 ;
	7'h41 :
		TR_58 = RG_rl_229 ;
	7'h42 :
		TR_58 = RG_rl_229 ;
	7'h43 :
		TR_58 = RG_rl_229 ;
	7'h44 :
		TR_58 = RG_rl_229 ;
	7'h45 :
		TR_58 = RG_rl_229 ;
	7'h46 :
		TR_58 = RG_rl_229 ;
	7'h47 :
		TR_58 = RG_rl_229 ;
	7'h48 :
		TR_58 = RG_rl_229 ;
	7'h49 :
		TR_58 = RG_rl_229 ;
	7'h4a :
		TR_58 = RG_rl_229 ;
	7'h4b :
		TR_58 = RG_rl_229 ;
	7'h4c :
		TR_58 = RG_rl_229 ;
	7'h4d :
		TR_58 = RG_rl_229 ;
	7'h4e :
		TR_58 = RG_rl_229 ;
	7'h4f :
		TR_58 = RG_rl_229 ;
	7'h50 :
		TR_58 = RG_rl_229 ;
	7'h51 :
		TR_58 = RG_rl_229 ;
	7'h52 :
		TR_58 = RG_rl_229 ;
	7'h53 :
		TR_58 = RG_rl_229 ;
	7'h54 :
		TR_58 = RG_rl_229 ;
	7'h55 :
		TR_58 = RG_rl_229 ;
	7'h56 :
		TR_58 = RG_rl_229 ;
	7'h57 :
		TR_58 = RG_rl_229 ;
	7'h58 :
		TR_58 = RG_rl_229 ;
	7'h59 :
		TR_58 = RG_rl_229 ;
	7'h5a :
		TR_58 = RG_rl_229 ;
	7'h5b :
		TR_58 = RG_rl_229 ;
	7'h5c :
		TR_58 = RG_rl_229 ;
	7'h5d :
		TR_58 = RG_rl_229 ;
	7'h5e :
		TR_58 = RG_rl_229 ;
	7'h5f :
		TR_58 = RG_rl_229 ;
	7'h60 :
		TR_58 = RG_rl_229 ;
	7'h61 :
		TR_58 = RG_rl_229 ;
	7'h62 :
		TR_58 = RG_rl_229 ;
	7'h63 :
		TR_58 = RG_rl_229 ;
	7'h64 :
		TR_58 = RG_rl_229 ;
	7'h65 :
		TR_58 = RG_rl_229 ;
	7'h66 :
		TR_58 = RG_rl_229 ;
	7'h67 :
		TR_58 = RG_rl_229 ;
	7'h68 :
		TR_58 = RG_rl_229 ;
	7'h69 :
		TR_58 = RG_rl_229 ;
	7'h6a :
		TR_58 = RG_rl_229 ;
	7'h6b :
		TR_58 = RG_rl_229 ;
	7'h6c :
		TR_58 = RG_rl_229 ;
	7'h6d :
		TR_58 = RG_rl_229 ;
	7'h6e :
		TR_58 = RG_rl_229 ;
	7'h6f :
		TR_58 = RG_rl_229 ;
	7'h70 :
		TR_58 = RG_rl_229 ;
	7'h71 :
		TR_58 = RG_rl_229 ;
	7'h72 :
		TR_58 = RG_rl_229 ;
	7'h73 :
		TR_58 = RG_rl_229 ;
	7'h74 :
		TR_58 = RG_rl_229 ;
	7'h75 :
		TR_58 = RG_rl_229 ;
	7'h76 :
		TR_58 = RG_rl_229 ;
	7'h77 :
		TR_58 = RG_rl_229 ;
	7'h78 :
		TR_58 = RG_rl_229 ;
	7'h79 :
		TR_58 = RG_rl_229 ;
	7'h7a :
		TR_58 = RG_rl_229 ;
	7'h7b :
		TR_58 = RG_rl_229 ;
	7'h7c :
		TR_58 = RG_rl_229 ;
	7'h7d :
		TR_58 = RG_rl_229 ;
	7'h7e :
		TR_58 = RG_rl_229 ;
	7'h7f :
		TR_58 = RG_rl_229 ;
	default :
		TR_58 = 9'hx ;
	endcase
always @ ( RG_rl_230 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_59 = RG_rl_230 ;
	7'h01 :
		TR_59 = RG_rl_230 ;
	7'h02 :
		TR_59 = RG_rl_230 ;
	7'h03 :
		TR_59 = RG_rl_230 ;
	7'h04 :
		TR_59 = RG_rl_230 ;
	7'h05 :
		TR_59 = RG_rl_230 ;
	7'h06 :
		TR_59 = RG_rl_230 ;
	7'h07 :
		TR_59 = RG_rl_230 ;
	7'h08 :
		TR_59 = RG_rl_230 ;
	7'h09 :
		TR_59 = RG_rl_230 ;
	7'h0a :
		TR_59 = RG_rl_230 ;
	7'h0b :
		TR_59 = RG_rl_230 ;
	7'h0c :
		TR_59 = RG_rl_230 ;
	7'h0d :
		TR_59 = RG_rl_230 ;
	7'h0e :
		TR_59 = RG_rl_230 ;
	7'h0f :
		TR_59 = RG_rl_230 ;
	7'h10 :
		TR_59 = RG_rl_230 ;
	7'h11 :
		TR_59 = RG_rl_230 ;
	7'h12 :
		TR_59 = RG_rl_230 ;
	7'h13 :
		TR_59 = RG_rl_230 ;
	7'h14 :
		TR_59 = RG_rl_230 ;
	7'h15 :
		TR_59 = RG_rl_230 ;
	7'h16 :
		TR_59 = RG_rl_230 ;
	7'h17 :
		TR_59 = RG_rl_230 ;
	7'h18 :
		TR_59 = RG_rl_230 ;
	7'h19 :
		TR_59 = RG_rl_230 ;
	7'h1a :
		TR_59 = RG_rl_230 ;
	7'h1b :
		TR_59 = RG_rl_230 ;
	7'h1c :
		TR_59 = RG_rl_230 ;
	7'h1d :
		TR_59 = RG_rl_230 ;
	7'h1e :
		TR_59 = RG_rl_230 ;
	7'h1f :
		TR_59 = RG_rl_230 ;
	7'h20 :
		TR_59 = RG_rl_230 ;
	7'h21 :
		TR_59 = RG_rl_230 ;
	7'h22 :
		TR_59 = RG_rl_230 ;
	7'h23 :
		TR_59 = RG_rl_230 ;
	7'h24 :
		TR_59 = RG_rl_230 ;
	7'h25 :
		TR_59 = RG_rl_230 ;
	7'h26 :
		TR_59 = RG_rl_230 ;
	7'h27 :
		TR_59 = RG_rl_230 ;
	7'h28 :
		TR_59 = RG_rl_230 ;
	7'h29 :
		TR_59 = RG_rl_230 ;
	7'h2a :
		TR_59 = RG_rl_230 ;
	7'h2b :
		TR_59 = RG_rl_230 ;
	7'h2c :
		TR_59 = RG_rl_230 ;
	7'h2d :
		TR_59 = RG_rl_230 ;
	7'h2e :
		TR_59 = RG_rl_230 ;
	7'h2f :
		TR_59 = 9'h000 ;	// line#=../rle.cpp:68
	7'h30 :
		TR_59 = RG_rl_230 ;
	7'h31 :
		TR_59 = RG_rl_230 ;
	7'h32 :
		TR_59 = RG_rl_230 ;
	7'h33 :
		TR_59 = RG_rl_230 ;
	7'h34 :
		TR_59 = RG_rl_230 ;
	7'h35 :
		TR_59 = RG_rl_230 ;
	7'h36 :
		TR_59 = RG_rl_230 ;
	7'h37 :
		TR_59 = RG_rl_230 ;
	7'h38 :
		TR_59 = RG_rl_230 ;
	7'h39 :
		TR_59 = RG_rl_230 ;
	7'h3a :
		TR_59 = RG_rl_230 ;
	7'h3b :
		TR_59 = RG_rl_230 ;
	7'h3c :
		TR_59 = RG_rl_230 ;
	7'h3d :
		TR_59 = RG_rl_230 ;
	7'h3e :
		TR_59 = RG_rl_230 ;
	7'h3f :
		TR_59 = RG_rl_230 ;
	7'h40 :
		TR_59 = RG_rl_230 ;
	7'h41 :
		TR_59 = RG_rl_230 ;
	7'h42 :
		TR_59 = RG_rl_230 ;
	7'h43 :
		TR_59 = RG_rl_230 ;
	7'h44 :
		TR_59 = RG_rl_230 ;
	7'h45 :
		TR_59 = RG_rl_230 ;
	7'h46 :
		TR_59 = RG_rl_230 ;
	7'h47 :
		TR_59 = RG_rl_230 ;
	7'h48 :
		TR_59 = RG_rl_230 ;
	7'h49 :
		TR_59 = RG_rl_230 ;
	7'h4a :
		TR_59 = RG_rl_230 ;
	7'h4b :
		TR_59 = RG_rl_230 ;
	7'h4c :
		TR_59 = RG_rl_230 ;
	7'h4d :
		TR_59 = RG_rl_230 ;
	7'h4e :
		TR_59 = RG_rl_230 ;
	7'h4f :
		TR_59 = RG_rl_230 ;
	7'h50 :
		TR_59 = RG_rl_230 ;
	7'h51 :
		TR_59 = RG_rl_230 ;
	7'h52 :
		TR_59 = RG_rl_230 ;
	7'h53 :
		TR_59 = RG_rl_230 ;
	7'h54 :
		TR_59 = RG_rl_230 ;
	7'h55 :
		TR_59 = RG_rl_230 ;
	7'h56 :
		TR_59 = RG_rl_230 ;
	7'h57 :
		TR_59 = RG_rl_230 ;
	7'h58 :
		TR_59 = RG_rl_230 ;
	7'h59 :
		TR_59 = RG_rl_230 ;
	7'h5a :
		TR_59 = RG_rl_230 ;
	7'h5b :
		TR_59 = RG_rl_230 ;
	7'h5c :
		TR_59 = RG_rl_230 ;
	7'h5d :
		TR_59 = RG_rl_230 ;
	7'h5e :
		TR_59 = RG_rl_230 ;
	7'h5f :
		TR_59 = RG_rl_230 ;
	7'h60 :
		TR_59 = RG_rl_230 ;
	7'h61 :
		TR_59 = RG_rl_230 ;
	7'h62 :
		TR_59 = RG_rl_230 ;
	7'h63 :
		TR_59 = RG_rl_230 ;
	7'h64 :
		TR_59 = RG_rl_230 ;
	7'h65 :
		TR_59 = RG_rl_230 ;
	7'h66 :
		TR_59 = RG_rl_230 ;
	7'h67 :
		TR_59 = RG_rl_230 ;
	7'h68 :
		TR_59 = RG_rl_230 ;
	7'h69 :
		TR_59 = RG_rl_230 ;
	7'h6a :
		TR_59 = RG_rl_230 ;
	7'h6b :
		TR_59 = RG_rl_230 ;
	7'h6c :
		TR_59 = RG_rl_230 ;
	7'h6d :
		TR_59 = RG_rl_230 ;
	7'h6e :
		TR_59 = RG_rl_230 ;
	7'h6f :
		TR_59 = RG_rl_230 ;
	7'h70 :
		TR_59 = RG_rl_230 ;
	7'h71 :
		TR_59 = RG_rl_230 ;
	7'h72 :
		TR_59 = RG_rl_230 ;
	7'h73 :
		TR_59 = RG_rl_230 ;
	7'h74 :
		TR_59 = RG_rl_230 ;
	7'h75 :
		TR_59 = RG_rl_230 ;
	7'h76 :
		TR_59 = RG_rl_230 ;
	7'h77 :
		TR_59 = RG_rl_230 ;
	7'h78 :
		TR_59 = RG_rl_230 ;
	7'h79 :
		TR_59 = RG_rl_230 ;
	7'h7a :
		TR_59 = RG_rl_230 ;
	7'h7b :
		TR_59 = RG_rl_230 ;
	7'h7c :
		TR_59 = RG_rl_230 ;
	7'h7d :
		TR_59 = RG_rl_230 ;
	7'h7e :
		TR_59 = RG_rl_230 ;
	7'h7f :
		TR_59 = RG_rl_230 ;
	default :
		TR_59 = 9'hx ;
	endcase
always @ ( RG_rl_231 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_60 = RG_rl_231 ;
	7'h01 :
		TR_60 = RG_rl_231 ;
	7'h02 :
		TR_60 = RG_rl_231 ;
	7'h03 :
		TR_60 = RG_rl_231 ;
	7'h04 :
		TR_60 = RG_rl_231 ;
	7'h05 :
		TR_60 = RG_rl_231 ;
	7'h06 :
		TR_60 = RG_rl_231 ;
	7'h07 :
		TR_60 = RG_rl_231 ;
	7'h08 :
		TR_60 = RG_rl_231 ;
	7'h09 :
		TR_60 = RG_rl_231 ;
	7'h0a :
		TR_60 = RG_rl_231 ;
	7'h0b :
		TR_60 = RG_rl_231 ;
	7'h0c :
		TR_60 = RG_rl_231 ;
	7'h0d :
		TR_60 = RG_rl_231 ;
	7'h0e :
		TR_60 = RG_rl_231 ;
	7'h0f :
		TR_60 = RG_rl_231 ;
	7'h10 :
		TR_60 = RG_rl_231 ;
	7'h11 :
		TR_60 = RG_rl_231 ;
	7'h12 :
		TR_60 = RG_rl_231 ;
	7'h13 :
		TR_60 = RG_rl_231 ;
	7'h14 :
		TR_60 = RG_rl_231 ;
	7'h15 :
		TR_60 = RG_rl_231 ;
	7'h16 :
		TR_60 = RG_rl_231 ;
	7'h17 :
		TR_60 = RG_rl_231 ;
	7'h18 :
		TR_60 = RG_rl_231 ;
	7'h19 :
		TR_60 = RG_rl_231 ;
	7'h1a :
		TR_60 = RG_rl_231 ;
	7'h1b :
		TR_60 = RG_rl_231 ;
	7'h1c :
		TR_60 = RG_rl_231 ;
	7'h1d :
		TR_60 = RG_rl_231 ;
	7'h1e :
		TR_60 = RG_rl_231 ;
	7'h1f :
		TR_60 = RG_rl_231 ;
	7'h20 :
		TR_60 = RG_rl_231 ;
	7'h21 :
		TR_60 = RG_rl_231 ;
	7'h22 :
		TR_60 = RG_rl_231 ;
	7'h23 :
		TR_60 = RG_rl_231 ;
	7'h24 :
		TR_60 = RG_rl_231 ;
	7'h25 :
		TR_60 = RG_rl_231 ;
	7'h26 :
		TR_60 = RG_rl_231 ;
	7'h27 :
		TR_60 = RG_rl_231 ;
	7'h28 :
		TR_60 = RG_rl_231 ;
	7'h29 :
		TR_60 = RG_rl_231 ;
	7'h2a :
		TR_60 = RG_rl_231 ;
	7'h2b :
		TR_60 = RG_rl_231 ;
	7'h2c :
		TR_60 = RG_rl_231 ;
	7'h2d :
		TR_60 = RG_rl_231 ;
	7'h2e :
		TR_60 = RG_rl_231 ;
	7'h2f :
		TR_60 = RG_rl_231 ;
	7'h30 :
		TR_60 = 9'h000 ;	// line#=../rle.cpp:68
	7'h31 :
		TR_60 = RG_rl_231 ;
	7'h32 :
		TR_60 = RG_rl_231 ;
	7'h33 :
		TR_60 = RG_rl_231 ;
	7'h34 :
		TR_60 = RG_rl_231 ;
	7'h35 :
		TR_60 = RG_rl_231 ;
	7'h36 :
		TR_60 = RG_rl_231 ;
	7'h37 :
		TR_60 = RG_rl_231 ;
	7'h38 :
		TR_60 = RG_rl_231 ;
	7'h39 :
		TR_60 = RG_rl_231 ;
	7'h3a :
		TR_60 = RG_rl_231 ;
	7'h3b :
		TR_60 = RG_rl_231 ;
	7'h3c :
		TR_60 = RG_rl_231 ;
	7'h3d :
		TR_60 = RG_rl_231 ;
	7'h3e :
		TR_60 = RG_rl_231 ;
	7'h3f :
		TR_60 = RG_rl_231 ;
	7'h40 :
		TR_60 = RG_rl_231 ;
	7'h41 :
		TR_60 = RG_rl_231 ;
	7'h42 :
		TR_60 = RG_rl_231 ;
	7'h43 :
		TR_60 = RG_rl_231 ;
	7'h44 :
		TR_60 = RG_rl_231 ;
	7'h45 :
		TR_60 = RG_rl_231 ;
	7'h46 :
		TR_60 = RG_rl_231 ;
	7'h47 :
		TR_60 = RG_rl_231 ;
	7'h48 :
		TR_60 = RG_rl_231 ;
	7'h49 :
		TR_60 = RG_rl_231 ;
	7'h4a :
		TR_60 = RG_rl_231 ;
	7'h4b :
		TR_60 = RG_rl_231 ;
	7'h4c :
		TR_60 = RG_rl_231 ;
	7'h4d :
		TR_60 = RG_rl_231 ;
	7'h4e :
		TR_60 = RG_rl_231 ;
	7'h4f :
		TR_60 = RG_rl_231 ;
	7'h50 :
		TR_60 = RG_rl_231 ;
	7'h51 :
		TR_60 = RG_rl_231 ;
	7'h52 :
		TR_60 = RG_rl_231 ;
	7'h53 :
		TR_60 = RG_rl_231 ;
	7'h54 :
		TR_60 = RG_rl_231 ;
	7'h55 :
		TR_60 = RG_rl_231 ;
	7'h56 :
		TR_60 = RG_rl_231 ;
	7'h57 :
		TR_60 = RG_rl_231 ;
	7'h58 :
		TR_60 = RG_rl_231 ;
	7'h59 :
		TR_60 = RG_rl_231 ;
	7'h5a :
		TR_60 = RG_rl_231 ;
	7'h5b :
		TR_60 = RG_rl_231 ;
	7'h5c :
		TR_60 = RG_rl_231 ;
	7'h5d :
		TR_60 = RG_rl_231 ;
	7'h5e :
		TR_60 = RG_rl_231 ;
	7'h5f :
		TR_60 = RG_rl_231 ;
	7'h60 :
		TR_60 = RG_rl_231 ;
	7'h61 :
		TR_60 = RG_rl_231 ;
	7'h62 :
		TR_60 = RG_rl_231 ;
	7'h63 :
		TR_60 = RG_rl_231 ;
	7'h64 :
		TR_60 = RG_rl_231 ;
	7'h65 :
		TR_60 = RG_rl_231 ;
	7'h66 :
		TR_60 = RG_rl_231 ;
	7'h67 :
		TR_60 = RG_rl_231 ;
	7'h68 :
		TR_60 = RG_rl_231 ;
	7'h69 :
		TR_60 = RG_rl_231 ;
	7'h6a :
		TR_60 = RG_rl_231 ;
	7'h6b :
		TR_60 = RG_rl_231 ;
	7'h6c :
		TR_60 = RG_rl_231 ;
	7'h6d :
		TR_60 = RG_rl_231 ;
	7'h6e :
		TR_60 = RG_rl_231 ;
	7'h6f :
		TR_60 = RG_rl_231 ;
	7'h70 :
		TR_60 = RG_rl_231 ;
	7'h71 :
		TR_60 = RG_rl_231 ;
	7'h72 :
		TR_60 = RG_rl_231 ;
	7'h73 :
		TR_60 = RG_rl_231 ;
	7'h74 :
		TR_60 = RG_rl_231 ;
	7'h75 :
		TR_60 = RG_rl_231 ;
	7'h76 :
		TR_60 = RG_rl_231 ;
	7'h77 :
		TR_60 = RG_rl_231 ;
	7'h78 :
		TR_60 = RG_rl_231 ;
	7'h79 :
		TR_60 = RG_rl_231 ;
	7'h7a :
		TR_60 = RG_rl_231 ;
	7'h7b :
		TR_60 = RG_rl_231 ;
	7'h7c :
		TR_60 = RG_rl_231 ;
	7'h7d :
		TR_60 = RG_rl_231 ;
	7'h7e :
		TR_60 = RG_rl_231 ;
	7'h7f :
		TR_60 = RG_rl_231 ;
	default :
		TR_60 = 9'hx ;
	endcase
always @ ( RG_rl_232 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_61 = RG_rl_232 ;
	7'h01 :
		TR_61 = RG_rl_232 ;
	7'h02 :
		TR_61 = RG_rl_232 ;
	7'h03 :
		TR_61 = RG_rl_232 ;
	7'h04 :
		TR_61 = RG_rl_232 ;
	7'h05 :
		TR_61 = RG_rl_232 ;
	7'h06 :
		TR_61 = RG_rl_232 ;
	7'h07 :
		TR_61 = RG_rl_232 ;
	7'h08 :
		TR_61 = RG_rl_232 ;
	7'h09 :
		TR_61 = RG_rl_232 ;
	7'h0a :
		TR_61 = RG_rl_232 ;
	7'h0b :
		TR_61 = RG_rl_232 ;
	7'h0c :
		TR_61 = RG_rl_232 ;
	7'h0d :
		TR_61 = RG_rl_232 ;
	7'h0e :
		TR_61 = RG_rl_232 ;
	7'h0f :
		TR_61 = RG_rl_232 ;
	7'h10 :
		TR_61 = RG_rl_232 ;
	7'h11 :
		TR_61 = RG_rl_232 ;
	7'h12 :
		TR_61 = RG_rl_232 ;
	7'h13 :
		TR_61 = RG_rl_232 ;
	7'h14 :
		TR_61 = RG_rl_232 ;
	7'h15 :
		TR_61 = RG_rl_232 ;
	7'h16 :
		TR_61 = RG_rl_232 ;
	7'h17 :
		TR_61 = RG_rl_232 ;
	7'h18 :
		TR_61 = RG_rl_232 ;
	7'h19 :
		TR_61 = RG_rl_232 ;
	7'h1a :
		TR_61 = RG_rl_232 ;
	7'h1b :
		TR_61 = RG_rl_232 ;
	7'h1c :
		TR_61 = RG_rl_232 ;
	7'h1d :
		TR_61 = RG_rl_232 ;
	7'h1e :
		TR_61 = RG_rl_232 ;
	7'h1f :
		TR_61 = RG_rl_232 ;
	7'h20 :
		TR_61 = RG_rl_232 ;
	7'h21 :
		TR_61 = RG_rl_232 ;
	7'h22 :
		TR_61 = RG_rl_232 ;
	7'h23 :
		TR_61 = RG_rl_232 ;
	7'h24 :
		TR_61 = RG_rl_232 ;
	7'h25 :
		TR_61 = RG_rl_232 ;
	7'h26 :
		TR_61 = RG_rl_232 ;
	7'h27 :
		TR_61 = RG_rl_232 ;
	7'h28 :
		TR_61 = RG_rl_232 ;
	7'h29 :
		TR_61 = RG_rl_232 ;
	7'h2a :
		TR_61 = RG_rl_232 ;
	7'h2b :
		TR_61 = RG_rl_232 ;
	7'h2c :
		TR_61 = RG_rl_232 ;
	7'h2d :
		TR_61 = RG_rl_232 ;
	7'h2e :
		TR_61 = RG_rl_232 ;
	7'h2f :
		TR_61 = RG_rl_232 ;
	7'h30 :
		TR_61 = RG_rl_232 ;
	7'h31 :
		TR_61 = 9'h000 ;	// line#=../rle.cpp:68
	7'h32 :
		TR_61 = RG_rl_232 ;
	7'h33 :
		TR_61 = RG_rl_232 ;
	7'h34 :
		TR_61 = RG_rl_232 ;
	7'h35 :
		TR_61 = RG_rl_232 ;
	7'h36 :
		TR_61 = RG_rl_232 ;
	7'h37 :
		TR_61 = RG_rl_232 ;
	7'h38 :
		TR_61 = RG_rl_232 ;
	7'h39 :
		TR_61 = RG_rl_232 ;
	7'h3a :
		TR_61 = RG_rl_232 ;
	7'h3b :
		TR_61 = RG_rl_232 ;
	7'h3c :
		TR_61 = RG_rl_232 ;
	7'h3d :
		TR_61 = RG_rl_232 ;
	7'h3e :
		TR_61 = RG_rl_232 ;
	7'h3f :
		TR_61 = RG_rl_232 ;
	7'h40 :
		TR_61 = RG_rl_232 ;
	7'h41 :
		TR_61 = RG_rl_232 ;
	7'h42 :
		TR_61 = RG_rl_232 ;
	7'h43 :
		TR_61 = RG_rl_232 ;
	7'h44 :
		TR_61 = RG_rl_232 ;
	7'h45 :
		TR_61 = RG_rl_232 ;
	7'h46 :
		TR_61 = RG_rl_232 ;
	7'h47 :
		TR_61 = RG_rl_232 ;
	7'h48 :
		TR_61 = RG_rl_232 ;
	7'h49 :
		TR_61 = RG_rl_232 ;
	7'h4a :
		TR_61 = RG_rl_232 ;
	7'h4b :
		TR_61 = RG_rl_232 ;
	7'h4c :
		TR_61 = RG_rl_232 ;
	7'h4d :
		TR_61 = RG_rl_232 ;
	7'h4e :
		TR_61 = RG_rl_232 ;
	7'h4f :
		TR_61 = RG_rl_232 ;
	7'h50 :
		TR_61 = RG_rl_232 ;
	7'h51 :
		TR_61 = RG_rl_232 ;
	7'h52 :
		TR_61 = RG_rl_232 ;
	7'h53 :
		TR_61 = RG_rl_232 ;
	7'h54 :
		TR_61 = RG_rl_232 ;
	7'h55 :
		TR_61 = RG_rl_232 ;
	7'h56 :
		TR_61 = RG_rl_232 ;
	7'h57 :
		TR_61 = RG_rl_232 ;
	7'h58 :
		TR_61 = RG_rl_232 ;
	7'h59 :
		TR_61 = RG_rl_232 ;
	7'h5a :
		TR_61 = RG_rl_232 ;
	7'h5b :
		TR_61 = RG_rl_232 ;
	7'h5c :
		TR_61 = RG_rl_232 ;
	7'h5d :
		TR_61 = RG_rl_232 ;
	7'h5e :
		TR_61 = RG_rl_232 ;
	7'h5f :
		TR_61 = RG_rl_232 ;
	7'h60 :
		TR_61 = RG_rl_232 ;
	7'h61 :
		TR_61 = RG_rl_232 ;
	7'h62 :
		TR_61 = RG_rl_232 ;
	7'h63 :
		TR_61 = RG_rl_232 ;
	7'h64 :
		TR_61 = RG_rl_232 ;
	7'h65 :
		TR_61 = RG_rl_232 ;
	7'h66 :
		TR_61 = RG_rl_232 ;
	7'h67 :
		TR_61 = RG_rl_232 ;
	7'h68 :
		TR_61 = RG_rl_232 ;
	7'h69 :
		TR_61 = RG_rl_232 ;
	7'h6a :
		TR_61 = RG_rl_232 ;
	7'h6b :
		TR_61 = RG_rl_232 ;
	7'h6c :
		TR_61 = RG_rl_232 ;
	7'h6d :
		TR_61 = RG_rl_232 ;
	7'h6e :
		TR_61 = RG_rl_232 ;
	7'h6f :
		TR_61 = RG_rl_232 ;
	7'h70 :
		TR_61 = RG_rl_232 ;
	7'h71 :
		TR_61 = RG_rl_232 ;
	7'h72 :
		TR_61 = RG_rl_232 ;
	7'h73 :
		TR_61 = RG_rl_232 ;
	7'h74 :
		TR_61 = RG_rl_232 ;
	7'h75 :
		TR_61 = RG_rl_232 ;
	7'h76 :
		TR_61 = RG_rl_232 ;
	7'h77 :
		TR_61 = RG_rl_232 ;
	7'h78 :
		TR_61 = RG_rl_232 ;
	7'h79 :
		TR_61 = RG_rl_232 ;
	7'h7a :
		TR_61 = RG_rl_232 ;
	7'h7b :
		TR_61 = RG_rl_232 ;
	7'h7c :
		TR_61 = RG_rl_232 ;
	7'h7d :
		TR_61 = RG_rl_232 ;
	7'h7e :
		TR_61 = RG_rl_232 ;
	7'h7f :
		TR_61 = RG_rl_232 ;
	default :
		TR_61 = 9'hx ;
	endcase
always @ ( RG_rl_233 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_62 = RG_rl_233 ;
	7'h01 :
		TR_62 = RG_rl_233 ;
	7'h02 :
		TR_62 = RG_rl_233 ;
	7'h03 :
		TR_62 = RG_rl_233 ;
	7'h04 :
		TR_62 = RG_rl_233 ;
	7'h05 :
		TR_62 = RG_rl_233 ;
	7'h06 :
		TR_62 = RG_rl_233 ;
	7'h07 :
		TR_62 = RG_rl_233 ;
	7'h08 :
		TR_62 = RG_rl_233 ;
	7'h09 :
		TR_62 = RG_rl_233 ;
	7'h0a :
		TR_62 = RG_rl_233 ;
	7'h0b :
		TR_62 = RG_rl_233 ;
	7'h0c :
		TR_62 = RG_rl_233 ;
	7'h0d :
		TR_62 = RG_rl_233 ;
	7'h0e :
		TR_62 = RG_rl_233 ;
	7'h0f :
		TR_62 = RG_rl_233 ;
	7'h10 :
		TR_62 = RG_rl_233 ;
	7'h11 :
		TR_62 = RG_rl_233 ;
	7'h12 :
		TR_62 = RG_rl_233 ;
	7'h13 :
		TR_62 = RG_rl_233 ;
	7'h14 :
		TR_62 = RG_rl_233 ;
	7'h15 :
		TR_62 = RG_rl_233 ;
	7'h16 :
		TR_62 = RG_rl_233 ;
	7'h17 :
		TR_62 = RG_rl_233 ;
	7'h18 :
		TR_62 = RG_rl_233 ;
	7'h19 :
		TR_62 = RG_rl_233 ;
	7'h1a :
		TR_62 = RG_rl_233 ;
	7'h1b :
		TR_62 = RG_rl_233 ;
	7'h1c :
		TR_62 = RG_rl_233 ;
	7'h1d :
		TR_62 = RG_rl_233 ;
	7'h1e :
		TR_62 = RG_rl_233 ;
	7'h1f :
		TR_62 = RG_rl_233 ;
	7'h20 :
		TR_62 = RG_rl_233 ;
	7'h21 :
		TR_62 = RG_rl_233 ;
	7'h22 :
		TR_62 = RG_rl_233 ;
	7'h23 :
		TR_62 = RG_rl_233 ;
	7'h24 :
		TR_62 = RG_rl_233 ;
	7'h25 :
		TR_62 = RG_rl_233 ;
	7'h26 :
		TR_62 = RG_rl_233 ;
	7'h27 :
		TR_62 = RG_rl_233 ;
	7'h28 :
		TR_62 = RG_rl_233 ;
	7'h29 :
		TR_62 = RG_rl_233 ;
	7'h2a :
		TR_62 = RG_rl_233 ;
	7'h2b :
		TR_62 = RG_rl_233 ;
	7'h2c :
		TR_62 = RG_rl_233 ;
	7'h2d :
		TR_62 = RG_rl_233 ;
	7'h2e :
		TR_62 = RG_rl_233 ;
	7'h2f :
		TR_62 = RG_rl_233 ;
	7'h30 :
		TR_62 = RG_rl_233 ;
	7'h31 :
		TR_62 = RG_rl_233 ;
	7'h32 :
		TR_62 = 9'h000 ;	// line#=../rle.cpp:68
	7'h33 :
		TR_62 = RG_rl_233 ;
	7'h34 :
		TR_62 = RG_rl_233 ;
	7'h35 :
		TR_62 = RG_rl_233 ;
	7'h36 :
		TR_62 = RG_rl_233 ;
	7'h37 :
		TR_62 = RG_rl_233 ;
	7'h38 :
		TR_62 = RG_rl_233 ;
	7'h39 :
		TR_62 = RG_rl_233 ;
	7'h3a :
		TR_62 = RG_rl_233 ;
	7'h3b :
		TR_62 = RG_rl_233 ;
	7'h3c :
		TR_62 = RG_rl_233 ;
	7'h3d :
		TR_62 = RG_rl_233 ;
	7'h3e :
		TR_62 = RG_rl_233 ;
	7'h3f :
		TR_62 = RG_rl_233 ;
	7'h40 :
		TR_62 = RG_rl_233 ;
	7'h41 :
		TR_62 = RG_rl_233 ;
	7'h42 :
		TR_62 = RG_rl_233 ;
	7'h43 :
		TR_62 = RG_rl_233 ;
	7'h44 :
		TR_62 = RG_rl_233 ;
	7'h45 :
		TR_62 = RG_rl_233 ;
	7'h46 :
		TR_62 = RG_rl_233 ;
	7'h47 :
		TR_62 = RG_rl_233 ;
	7'h48 :
		TR_62 = RG_rl_233 ;
	7'h49 :
		TR_62 = RG_rl_233 ;
	7'h4a :
		TR_62 = RG_rl_233 ;
	7'h4b :
		TR_62 = RG_rl_233 ;
	7'h4c :
		TR_62 = RG_rl_233 ;
	7'h4d :
		TR_62 = RG_rl_233 ;
	7'h4e :
		TR_62 = RG_rl_233 ;
	7'h4f :
		TR_62 = RG_rl_233 ;
	7'h50 :
		TR_62 = RG_rl_233 ;
	7'h51 :
		TR_62 = RG_rl_233 ;
	7'h52 :
		TR_62 = RG_rl_233 ;
	7'h53 :
		TR_62 = RG_rl_233 ;
	7'h54 :
		TR_62 = RG_rl_233 ;
	7'h55 :
		TR_62 = RG_rl_233 ;
	7'h56 :
		TR_62 = RG_rl_233 ;
	7'h57 :
		TR_62 = RG_rl_233 ;
	7'h58 :
		TR_62 = RG_rl_233 ;
	7'h59 :
		TR_62 = RG_rl_233 ;
	7'h5a :
		TR_62 = RG_rl_233 ;
	7'h5b :
		TR_62 = RG_rl_233 ;
	7'h5c :
		TR_62 = RG_rl_233 ;
	7'h5d :
		TR_62 = RG_rl_233 ;
	7'h5e :
		TR_62 = RG_rl_233 ;
	7'h5f :
		TR_62 = RG_rl_233 ;
	7'h60 :
		TR_62 = RG_rl_233 ;
	7'h61 :
		TR_62 = RG_rl_233 ;
	7'h62 :
		TR_62 = RG_rl_233 ;
	7'h63 :
		TR_62 = RG_rl_233 ;
	7'h64 :
		TR_62 = RG_rl_233 ;
	7'h65 :
		TR_62 = RG_rl_233 ;
	7'h66 :
		TR_62 = RG_rl_233 ;
	7'h67 :
		TR_62 = RG_rl_233 ;
	7'h68 :
		TR_62 = RG_rl_233 ;
	7'h69 :
		TR_62 = RG_rl_233 ;
	7'h6a :
		TR_62 = RG_rl_233 ;
	7'h6b :
		TR_62 = RG_rl_233 ;
	7'h6c :
		TR_62 = RG_rl_233 ;
	7'h6d :
		TR_62 = RG_rl_233 ;
	7'h6e :
		TR_62 = RG_rl_233 ;
	7'h6f :
		TR_62 = RG_rl_233 ;
	7'h70 :
		TR_62 = RG_rl_233 ;
	7'h71 :
		TR_62 = RG_rl_233 ;
	7'h72 :
		TR_62 = RG_rl_233 ;
	7'h73 :
		TR_62 = RG_rl_233 ;
	7'h74 :
		TR_62 = RG_rl_233 ;
	7'h75 :
		TR_62 = RG_rl_233 ;
	7'h76 :
		TR_62 = RG_rl_233 ;
	7'h77 :
		TR_62 = RG_rl_233 ;
	7'h78 :
		TR_62 = RG_rl_233 ;
	7'h79 :
		TR_62 = RG_rl_233 ;
	7'h7a :
		TR_62 = RG_rl_233 ;
	7'h7b :
		TR_62 = RG_rl_233 ;
	7'h7c :
		TR_62 = RG_rl_233 ;
	7'h7d :
		TR_62 = RG_rl_233 ;
	7'h7e :
		TR_62 = RG_rl_233 ;
	7'h7f :
		TR_62 = RG_rl_233 ;
	default :
		TR_62 = 9'hx ;
	endcase
always @ ( RG_rl_234 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_63 = RG_rl_234 ;
	7'h01 :
		TR_63 = RG_rl_234 ;
	7'h02 :
		TR_63 = RG_rl_234 ;
	7'h03 :
		TR_63 = RG_rl_234 ;
	7'h04 :
		TR_63 = RG_rl_234 ;
	7'h05 :
		TR_63 = RG_rl_234 ;
	7'h06 :
		TR_63 = RG_rl_234 ;
	7'h07 :
		TR_63 = RG_rl_234 ;
	7'h08 :
		TR_63 = RG_rl_234 ;
	7'h09 :
		TR_63 = RG_rl_234 ;
	7'h0a :
		TR_63 = RG_rl_234 ;
	7'h0b :
		TR_63 = RG_rl_234 ;
	7'h0c :
		TR_63 = RG_rl_234 ;
	7'h0d :
		TR_63 = RG_rl_234 ;
	7'h0e :
		TR_63 = RG_rl_234 ;
	7'h0f :
		TR_63 = RG_rl_234 ;
	7'h10 :
		TR_63 = RG_rl_234 ;
	7'h11 :
		TR_63 = RG_rl_234 ;
	7'h12 :
		TR_63 = RG_rl_234 ;
	7'h13 :
		TR_63 = RG_rl_234 ;
	7'h14 :
		TR_63 = RG_rl_234 ;
	7'h15 :
		TR_63 = RG_rl_234 ;
	7'h16 :
		TR_63 = RG_rl_234 ;
	7'h17 :
		TR_63 = RG_rl_234 ;
	7'h18 :
		TR_63 = RG_rl_234 ;
	7'h19 :
		TR_63 = RG_rl_234 ;
	7'h1a :
		TR_63 = RG_rl_234 ;
	7'h1b :
		TR_63 = RG_rl_234 ;
	7'h1c :
		TR_63 = RG_rl_234 ;
	7'h1d :
		TR_63 = RG_rl_234 ;
	7'h1e :
		TR_63 = RG_rl_234 ;
	7'h1f :
		TR_63 = RG_rl_234 ;
	7'h20 :
		TR_63 = RG_rl_234 ;
	7'h21 :
		TR_63 = RG_rl_234 ;
	7'h22 :
		TR_63 = RG_rl_234 ;
	7'h23 :
		TR_63 = RG_rl_234 ;
	7'h24 :
		TR_63 = RG_rl_234 ;
	7'h25 :
		TR_63 = RG_rl_234 ;
	7'h26 :
		TR_63 = RG_rl_234 ;
	7'h27 :
		TR_63 = RG_rl_234 ;
	7'h28 :
		TR_63 = RG_rl_234 ;
	7'h29 :
		TR_63 = RG_rl_234 ;
	7'h2a :
		TR_63 = RG_rl_234 ;
	7'h2b :
		TR_63 = RG_rl_234 ;
	7'h2c :
		TR_63 = RG_rl_234 ;
	7'h2d :
		TR_63 = RG_rl_234 ;
	7'h2e :
		TR_63 = RG_rl_234 ;
	7'h2f :
		TR_63 = RG_rl_234 ;
	7'h30 :
		TR_63 = RG_rl_234 ;
	7'h31 :
		TR_63 = RG_rl_234 ;
	7'h32 :
		TR_63 = RG_rl_234 ;
	7'h33 :
		TR_63 = 9'h000 ;	// line#=../rle.cpp:68
	7'h34 :
		TR_63 = RG_rl_234 ;
	7'h35 :
		TR_63 = RG_rl_234 ;
	7'h36 :
		TR_63 = RG_rl_234 ;
	7'h37 :
		TR_63 = RG_rl_234 ;
	7'h38 :
		TR_63 = RG_rl_234 ;
	7'h39 :
		TR_63 = RG_rl_234 ;
	7'h3a :
		TR_63 = RG_rl_234 ;
	7'h3b :
		TR_63 = RG_rl_234 ;
	7'h3c :
		TR_63 = RG_rl_234 ;
	7'h3d :
		TR_63 = RG_rl_234 ;
	7'h3e :
		TR_63 = RG_rl_234 ;
	7'h3f :
		TR_63 = RG_rl_234 ;
	7'h40 :
		TR_63 = RG_rl_234 ;
	7'h41 :
		TR_63 = RG_rl_234 ;
	7'h42 :
		TR_63 = RG_rl_234 ;
	7'h43 :
		TR_63 = RG_rl_234 ;
	7'h44 :
		TR_63 = RG_rl_234 ;
	7'h45 :
		TR_63 = RG_rl_234 ;
	7'h46 :
		TR_63 = RG_rl_234 ;
	7'h47 :
		TR_63 = RG_rl_234 ;
	7'h48 :
		TR_63 = RG_rl_234 ;
	7'h49 :
		TR_63 = RG_rl_234 ;
	7'h4a :
		TR_63 = RG_rl_234 ;
	7'h4b :
		TR_63 = RG_rl_234 ;
	7'h4c :
		TR_63 = RG_rl_234 ;
	7'h4d :
		TR_63 = RG_rl_234 ;
	7'h4e :
		TR_63 = RG_rl_234 ;
	7'h4f :
		TR_63 = RG_rl_234 ;
	7'h50 :
		TR_63 = RG_rl_234 ;
	7'h51 :
		TR_63 = RG_rl_234 ;
	7'h52 :
		TR_63 = RG_rl_234 ;
	7'h53 :
		TR_63 = RG_rl_234 ;
	7'h54 :
		TR_63 = RG_rl_234 ;
	7'h55 :
		TR_63 = RG_rl_234 ;
	7'h56 :
		TR_63 = RG_rl_234 ;
	7'h57 :
		TR_63 = RG_rl_234 ;
	7'h58 :
		TR_63 = RG_rl_234 ;
	7'h59 :
		TR_63 = RG_rl_234 ;
	7'h5a :
		TR_63 = RG_rl_234 ;
	7'h5b :
		TR_63 = RG_rl_234 ;
	7'h5c :
		TR_63 = RG_rl_234 ;
	7'h5d :
		TR_63 = RG_rl_234 ;
	7'h5e :
		TR_63 = RG_rl_234 ;
	7'h5f :
		TR_63 = RG_rl_234 ;
	7'h60 :
		TR_63 = RG_rl_234 ;
	7'h61 :
		TR_63 = RG_rl_234 ;
	7'h62 :
		TR_63 = RG_rl_234 ;
	7'h63 :
		TR_63 = RG_rl_234 ;
	7'h64 :
		TR_63 = RG_rl_234 ;
	7'h65 :
		TR_63 = RG_rl_234 ;
	7'h66 :
		TR_63 = RG_rl_234 ;
	7'h67 :
		TR_63 = RG_rl_234 ;
	7'h68 :
		TR_63 = RG_rl_234 ;
	7'h69 :
		TR_63 = RG_rl_234 ;
	7'h6a :
		TR_63 = RG_rl_234 ;
	7'h6b :
		TR_63 = RG_rl_234 ;
	7'h6c :
		TR_63 = RG_rl_234 ;
	7'h6d :
		TR_63 = RG_rl_234 ;
	7'h6e :
		TR_63 = RG_rl_234 ;
	7'h6f :
		TR_63 = RG_rl_234 ;
	7'h70 :
		TR_63 = RG_rl_234 ;
	7'h71 :
		TR_63 = RG_rl_234 ;
	7'h72 :
		TR_63 = RG_rl_234 ;
	7'h73 :
		TR_63 = RG_rl_234 ;
	7'h74 :
		TR_63 = RG_rl_234 ;
	7'h75 :
		TR_63 = RG_rl_234 ;
	7'h76 :
		TR_63 = RG_rl_234 ;
	7'h77 :
		TR_63 = RG_rl_234 ;
	7'h78 :
		TR_63 = RG_rl_234 ;
	7'h79 :
		TR_63 = RG_rl_234 ;
	7'h7a :
		TR_63 = RG_rl_234 ;
	7'h7b :
		TR_63 = RG_rl_234 ;
	7'h7c :
		TR_63 = RG_rl_234 ;
	7'h7d :
		TR_63 = RG_rl_234 ;
	7'h7e :
		TR_63 = RG_rl_234 ;
	7'h7f :
		TR_63 = RG_rl_234 ;
	default :
		TR_63 = 9'hx ;
	endcase
always @ ( RG_rl_235 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_64 = RG_rl_235 ;
	7'h01 :
		TR_64 = RG_rl_235 ;
	7'h02 :
		TR_64 = RG_rl_235 ;
	7'h03 :
		TR_64 = RG_rl_235 ;
	7'h04 :
		TR_64 = RG_rl_235 ;
	7'h05 :
		TR_64 = RG_rl_235 ;
	7'h06 :
		TR_64 = RG_rl_235 ;
	7'h07 :
		TR_64 = RG_rl_235 ;
	7'h08 :
		TR_64 = RG_rl_235 ;
	7'h09 :
		TR_64 = RG_rl_235 ;
	7'h0a :
		TR_64 = RG_rl_235 ;
	7'h0b :
		TR_64 = RG_rl_235 ;
	7'h0c :
		TR_64 = RG_rl_235 ;
	7'h0d :
		TR_64 = RG_rl_235 ;
	7'h0e :
		TR_64 = RG_rl_235 ;
	7'h0f :
		TR_64 = RG_rl_235 ;
	7'h10 :
		TR_64 = RG_rl_235 ;
	7'h11 :
		TR_64 = RG_rl_235 ;
	7'h12 :
		TR_64 = RG_rl_235 ;
	7'h13 :
		TR_64 = RG_rl_235 ;
	7'h14 :
		TR_64 = RG_rl_235 ;
	7'h15 :
		TR_64 = RG_rl_235 ;
	7'h16 :
		TR_64 = RG_rl_235 ;
	7'h17 :
		TR_64 = RG_rl_235 ;
	7'h18 :
		TR_64 = RG_rl_235 ;
	7'h19 :
		TR_64 = RG_rl_235 ;
	7'h1a :
		TR_64 = RG_rl_235 ;
	7'h1b :
		TR_64 = RG_rl_235 ;
	7'h1c :
		TR_64 = RG_rl_235 ;
	7'h1d :
		TR_64 = RG_rl_235 ;
	7'h1e :
		TR_64 = RG_rl_235 ;
	7'h1f :
		TR_64 = RG_rl_235 ;
	7'h20 :
		TR_64 = RG_rl_235 ;
	7'h21 :
		TR_64 = RG_rl_235 ;
	7'h22 :
		TR_64 = RG_rl_235 ;
	7'h23 :
		TR_64 = RG_rl_235 ;
	7'h24 :
		TR_64 = RG_rl_235 ;
	7'h25 :
		TR_64 = RG_rl_235 ;
	7'h26 :
		TR_64 = RG_rl_235 ;
	7'h27 :
		TR_64 = RG_rl_235 ;
	7'h28 :
		TR_64 = RG_rl_235 ;
	7'h29 :
		TR_64 = RG_rl_235 ;
	7'h2a :
		TR_64 = RG_rl_235 ;
	7'h2b :
		TR_64 = RG_rl_235 ;
	7'h2c :
		TR_64 = RG_rl_235 ;
	7'h2d :
		TR_64 = RG_rl_235 ;
	7'h2e :
		TR_64 = RG_rl_235 ;
	7'h2f :
		TR_64 = RG_rl_235 ;
	7'h30 :
		TR_64 = RG_rl_235 ;
	7'h31 :
		TR_64 = RG_rl_235 ;
	7'h32 :
		TR_64 = RG_rl_235 ;
	7'h33 :
		TR_64 = RG_rl_235 ;
	7'h34 :
		TR_64 = 9'h000 ;	// line#=../rle.cpp:68
	7'h35 :
		TR_64 = RG_rl_235 ;
	7'h36 :
		TR_64 = RG_rl_235 ;
	7'h37 :
		TR_64 = RG_rl_235 ;
	7'h38 :
		TR_64 = RG_rl_235 ;
	7'h39 :
		TR_64 = RG_rl_235 ;
	7'h3a :
		TR_64 = RG_rl_235 ;
	7'h3b :
		TR_64 = RG_rl_235 ;
	7'h3c :
		TR_64 = RG_rl_235 ;
	7'h3d :
		TR_64 = RG_rl_235 ;
	7'h3e :
		TR_64 = RG_rl_235 ;
	7'h3f :
		TR_64 = RG_rl_235 ;
	7'h40 :
		TR_64 = RG_rl_235 ;
	7'h41 :
		TR_64 = RG_rl_235 ;
	7'h42 :
		TR_64 = RG_rl_235 ;
	7'h43 :
		TR_64 = RG_rl_235 ;
	7'h44 :
		TR_64 = RG_rl_235 ;
	7'h45 :
		TR_64 = RG_rl_235 ;
	7'h46 :
		TR_64 = RG_rl_235 ;
	7'h47 :
		TR_64 = RG_rl_235 ;
	7'h48 :
		TR_64 = RG_rl_235 ;
	7'h49 :
		TR_64 = RG_rl_235 ;
	7'h4a :
		TR_64 = RG_rl_235 ;
	7'h4b :
		TR_64 = RG_rl_235 ;
	7'h4c :
		TR_64 = RG_rl_235 ;
	7'h4d :
		TR_64 = RG_rl_235 ;
	7'h4e :
		TR_64 = RG_rl_235 ;
	7'h4f :
		TR_64 = RG_rl_235 ;
	7'h50 :
		TR_64 = RG_rl_235 ;
	7'h51 :
		TR_64 = RG_rl_235 ;
	7'h52 :
		TR_64 = RG_rl_235 ;
	7'h53 :
		TR_64 = RG_rl_235 ;
	7'h54 :
		TR_64 = RG_rl_235 ;
	7'h55 :
		TR_64 = RG_rl_235 ;
	7'h56 :
		TR_64 = RG_rl_235 ;
	7'h57 :
		TR_64 = RG_rl_235 ;
	7'h58 :
		TR_64 = RG_rl_235 ;
	7'h59 :
		TR_64 = RG_rl_235 ;
	7'h5a :
		TR_64 = RG_rl_235 ;
	7'h5b :
		TR_64 = RG_rl_235 ;
	7'h5c :
		TR_64 = RG_rl_235 ;
	7'h5d :
		TR_64 = RG_rl_235 ;
	7'h5e :
		TR_64 = RG_rl_235 ;
	7'h5f :
		TR_64 = RG_rl_235 ;
	7'h60 :
		TR_64 = RG_rl_235 ;
	7'h61 :
		TR_64 = RG_rl_235 ;
	7'h62 :
		TR_64 = RG_rl_235 ;
	7'h63 :
		TR_64 = RG_rl_235 ;
	7'h64 :
		TR_64 = RG_rl_235 ;
	7'h65 :
		TR_64 = RG_rl_235 ;
	7'h66 :
		TR_64 = RG_rl_235 ;
	7'h67 :
		TR_64 = RG_rl_235 ;
	7'h68 :
		TR_64 = RG_rl_235 ;
	7'h69 :
		TR_64 = RG_rl_235 ;
	7'h6a :
		TR_64 = RG_rl_235 ;
	7'h6b :
		TR_64 = RG_rl_235 ;
	7'h6c :
		TR_64 = RG_rl_235 ;
	7'h6d :
		TR_64 = RG_rl_235 ;
	7'h6e :
		TR_64 = RG_rl_235 ;
	7'h6f :
		TR_64 = RG_rl_235 ;
	7'h70 :
		TR_64 = RG_rl_235 ;
	7'h71 :
		TR_64 = RG_rl_235 ;
	7'h72 :
		TR_64 = RG_rl_235 ;
	7'h73 :
		TR_64 = RG_rl_235 ;
	7'h74 :
		TR_64 = RG_rl_235 ;
	7'h75 :
		TR_64 = RG_rl_235 ;
	7'h76 :
		TR_64 = RG_rl_235 ;
	7'h77 :
		TR_64 = RG_rl_235 ;
	7'h78 :
		TR_64 = RG_rl_235 ;
	7'h79 :
		TR_64 = RG_rl_235 ;
	7'h7a :
		TR_64 = RG_rl_235 ;
	7'h7b :
		TR_64 = RG_rl_235 ;
	7'h7c :
		TR_64 = RG_rl_235 ;
	7'h7d :
		TR_64 = RG_rl_235 ;
	7'h7e :
		TR_64 = RG_rl_235 ;
	7'h7f :
		TR_64 = RG_rl_235 ;
	default :
		TR_64 = 9'hx ;
	endcase
always @ ( RG_rl_236 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_65 = RG_rl_236 ;
	7'h01 :
		TR_65 = RG_rl_236 ;
	7'h02 :
		TR_65 = RG_rl_236 ;
	7'h03 :
		TR_65 = RG_rl_236 ;
	7'h04 :
		TR_65 = RG_rl_236 ;
	7'h05 :
		TR_65 = RG_rl_236 ;
	7'h06 :
		TR_65 = RG_rl_236 ;
	7'h07 :
		TR_65 = RG_rl_236 ;
	7'h08 :
		TR_65 = RG_rl_236 ;
	7'h09 :
		TR_65 = RG_rl_236 ;
	7'h0a :
		TR_65 = RG_rl_236 ;
	7'h0b :
		TR_65 = RG_rl_236 ;
	7'h0c :
		TR_65 = RG_rl_236 ;
	7'h0d :
		TR_65 = RG_rl_236 ;
	7'h0e :
		TR_65 = RG_rl_236 ;
	7'h0f :
		TR_65 = RG_rl_236 ;
	7'h10 :
		TR_65 = RG_rl_236 ;
	7'h11 :
		TR_65 = RG_rl_236 ;
	7'h12 :
		TR_65 = RG_rl_236 ;
	7'h13 :
		TR_65 = RG_rl_236 ;
	7'h14 :
		TR_65 = RG_rl_236 ;
	7'h15 :
		TR_65 = RG_rl_236 ;
	7'h16 :
		TR_65 = RG_rl_236 ;
	7'h17 :
		TR_65 = RG_rl_236 ;
	7'h18 :
		TR_65 = RG_rl_236 ;
	7'h19 :
		TR_65 = RG_rl_236 ;
	7'h1a :
		TR_65 = RG_rl_236 ;
	7'h1b :
		TR_65 = RG_rl_236 ;
	7'h1c :
		TR_65 = RG_rl_236 ;
	7'h1d :
		TR_65 = RG_rl_236 ;
	7'h1e :
		TR_65 = RG_rl_236 ;
	7'h1f :
		TR_65 = RG_rl_236 ;
	7'h20 :
		TR_65 = RG_rl_236 ;
	7'h21 :
		TR_65 = RG_rl_236 ;
	7'h22 :
		TR_65 = RG_rl_236 ;
	7'h23 :
		TR_65 = RG_rl_236 ;
	7'h24 :
		TR_65 = RG_rl_236 ;
	7'h25 :
		TR_65 = RG_rl_236 ;
	7'h26 :
		TR_65 = RG_rl_236 ;
	7'h27 :
		TR_65 = RG_rl_236 ;
	7'h28 :
		TR_65 = RG_rl_236 ;
	7'h29 :
		TR_65 = RG_rl_236 ;
	7'h2a :
		TR_65 = RG_rl_236 ;
	7'h2b :
		TR_65 = RG_rl_236 ;
	7'h2c :
		TR_65 = RG_rl_236 ;
	7'h2d :
		TR_65 = RG_rl_236 ;
	7'h2e :
		TR_65 = RG_rl_236 ;
	7'h2f :
		TR_65 = RG_rl_236 ;
	7'h30 :
		TR_65 = RG_rl_236 ;
	7'h31 :
		TR_65 = RG_rl_236 ;
	7'h32 :
		TR_65 = RG_rl_236 ;
	7'h33 :
		TR_65 = RG_rl_236 ;
	7'h34 :
		TR_65 = RG_rl_236 ;
	7'h35 :
		TR_65 = 9'h000 ;	// line#=../rle.cpp:68
	7'h36 :
		TR_65 = RG_rl_236 ;
	7'h37 :
		TR_65 = RG_rl_236 ;
	7'h38 :
		TR_65 = RG_rl_236 ;
	7'h39 :
		TR_65 = RG_rl_236 ;
	7'h3a :
		TR_65 = RG_rl_236 ;
	7'h3b :
		TR_65 = RG_rl_236 ;
	7'h3c :
		TR_65 = RG_rl_236 ;
	7'h3d :
		TR_65 = RG_rl_236 ;
	7'h3e :
		TR_65 = RG_rl_236 ;
	7'h3f :
		TR_65 = RG_rl_236 ;
	7'h40 :
		TR_65 = RG_rl_236 ;
	7'h41 :
		TR_65 = RG_rl_236 ;
	7'h42 :
		TR_65 = RG_rl_236 ;
	7'h43 :
		TR_65 = RG_rl_236 ;
	7'h44 :
		TR_65 = RG_rl_236 ;
	7'h45 :
		TR_65 = RG_rl_236 ;
	7'h46 :
		TR_65 = RG_rl_236 ;
	7'h47 :
		TR_65 = RG_rl_236 ;
	7'h48 :
		TR_65 = RG_rl_236 ;
	7'h49 :
		TR_65 = RG_rl_236 ;
	7'h4a :
		TR_65 = RG_rl_236 ;
	7'h4b :
		TR_65 = RG_rl_236 ;
	7'h4c :
		TR_65 = RG_rl_236 ;
	7'h4d :
		TR_65 = RG_rl_236 ;
	7'h4e :
		TR_65 = RG_rl_236 ;
	7'h4f :
		TR_65 = RG_rl_236 ;
	7'h50 :
		TR_65 = RG_rl_236 ;
	7'h51 :
		TR_65 = RG_rl_236 ;
	7'h52 :
		TR_65 = RG_rl_236 ;
	7'h53 :
		TR_65 = RG_rl_236 ;
	7'h54 :
		TR_65 = RG_rl_236 ;
	7'h55 :
		TR_65 = RG_rl_236 ;
	7'h56 :
		TR_65 = RG_rl_236 ;
	7'h57 :
		TR_65 = RG_rl_236 ;
	7'h58 :
		TR_65 = RG_rl_236 ;
	7'h59 :
		TR_65 = RG_rl_236 ;
	7'h5a :
		TR_65 = RG_rl_236 ;
	7'h5b :
		TR_65 = RG_rl_236 ;
	7'h5c :
		TR_65 = RG_rl_236 ;
	7'h5d :
		TR_65 = RG_rl_236 ;
	7'h5e :
		TR_65 = RG_rl_236 ;
	7'h5f :
		TR_65 = RG_rl_236 ;
	7'h60 :
		TR_65 = RG_rl_236 ;
	7'h61 :
		TR_65 = RG_rl_236 ;
	7'h62 :
		TR_65 = RG_rl_236 ;
	7'h63 :
		TR_65 = RG_rl_236 ;
	7'h64 :
		TR_65 = RG_rl_236 ;
	7'h65 :
		TR_65 = RG_rl_236 ;
	7'h66 :
		TR_65 = RG_rl_236 ;
	7'h67 :
		TR_65 = RG_rl_236 ;
	7'h68 :
		TR_65 = RG_rl_236 ;
	7'h69 :
		TR_65 = RG_rl_236 ;
	7'h6a :
		TR_65 = RG_rl_236 ;
	7'h6b :
		TR_65 = RG_rl_236 ;
	7'h6c :
		TR_65 = RG_rl_236 ;
	7'h6d :
		TR_65 = RG_rl_236 ;
	7'h6e :
		TR_65 = RG_rl_236 ;
	7'h6f :
		TR_65 = RG_rl_236 ;
	7'h70 :
		TR_65 = RG_rl_236 ;
	7'h71 :
		TR_65 = RG_rl_236 ;
	7'h72 :
		TR_65 = RG_rl_236 ;
	7'h73 :
		TR_65 = RG_rl_236 ;
	7'h74 :
		TR_65 = RG_rl_236 ;
	7'h75 :
		TR_65 = RG_rl_236 ;
	7'h76 :
		TR_65 = RG_rl_236 ;
	7'h77 :
		TR_65 = RG_rl_236 ;
	7'h78 :
		TR_65 = RG_rl_236 ;
	7'h79 :
		TR_65 = RG_rl_236 ;
	7'h7a :
		TR_65 = RG_rl_236 ;
	7'h7b :
		TR_65 = RG_rl_236 ;
	7'h7c :
		TR_65 = RG_rl_236 ;
	7'h7d :
		TR_65 = RG_rl_236 ;
	7'h7e :
		TR_65 = RG_rl_236 ;
	7'h7f :
		TR_65 = RG_rl_236 ;
	default :
		TR_65 = 9'hx ;
	endcase
always @ ( RG_rl_237 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_66 = RG_rl_237 ;
	7'h01 :
		TR_66 = RG_rl_237 ;
	7'h02 :
		TR_66 = RG_rl_237 ;
	7'h03 :
		TR_66 = RG_rl_237 ;
	7'h04 :
		TR_66 = RG_rl_237 ;
	7'h05 :
		TR_66 = RG_rl_237 ;
	7'h06 :
		TR_66 = RG_rl_237 ;
	7'h07 :
		TR_66 = RG_rl_237 ;
	7'h08 :
		TR_66 = RG_rl_237 ;
	7'h09 :
		TR_66 = RG_rl_237 ;
	7'h0a :
		TR_66 = RG_rl_237 ;
	7'h0b :
		TR_66 = RG_rl_237 ;
	7'h0c :
		TR_66 = RG_rl_237 ;
	7'h0d :
		TR_66 = RG_rl_237 ;
	7'h0e :
		TR_66 = RG_rl_237 ;
	7'h0f :
		TR_66 = RG_rl_237 ;
	7'h10 :
		TR_66 = RG_rl_237 ;
	7'h11 :
		TR_66 = RG_rl_237 ;
	7'h12 :
		TR_66 = RG_rl_237 ;
	7'h13 :
		TR_66 = RG_rl_237 ;
	7'h14 :
		TR_66 = RG_rl_237 ;
	7'h15 :
		TR_66 = RG_rl_237 ;
	7'h16 :
		TR_66 = RG_rl_237 ;
	7'h17 :
		TR_66 = RG_rl_237 ;
	7'h18 :
		TR_66 = RG_rl_237 ;
	7'h19 :
		TR_66 = RG_rl_237 ;
	7'h1a :
		TR_66 = RG_rl_237 ;
	7'h1b :
		TR_66 = RG_rl_237 ;
	7'h1c :
		TR_66 = RG_rl_237 ;
	7'h1d :
		TR_66 = RG_rl_237 ;
	7'h1e :
		TR_66 = RG_rl_237 ;
	7'h1f :
		TR_66 = RG_rl_237 ;
	7'h20 :
		TR_66 = RG_rl_237 ;
	7'h21 :
		TR_66 = RG_rl_237 ;
	7'h22 :
		TR_66 = RG_rl_237 ;
	7'h23 :
		TR_66 = RG_rl_237 ;
	7'h24 :
		TR_66 = RG_rl_237 ;
	7'h25 :
		TR_66 = RG_rl_237 ;
	7'h26 :
		TR_66 = RG_rl_237 ;
	7'h27 :
		TR_66 = RG_rl_237 ;
	7'h28 :
		TR_66 = RG_rl_237 ;
	7'h29 :
		TR_66 = RG_rl_237 ;
	7'h2a :
		TR_66 = RG_rl_237 ;
	7'h2b :
		TR_66 = RG_rl_237 ;
	7'h2c :
		TR_66 = RG_rl_237 ;
	7'h2d :
		TR_66 = RG_rl_237 ;
	7'h2e :
		TR_66 = RG_rl_237 ;
	7'h2f :
		TR_66 = RG_rl_237 ;
	7'h30 :
		TR_66 = RG_rl_237 ;
	7'h31 :
		TR_66 = RG_rl_237 ;
	7'h32 :
		TR_66 = RG_rl_237 ;
	7'h33 :
		TR_66 = RG_rl_237 ;
	7'h34 :
		TR_66 = RG_rl_237 ;
	7'h35 :
		TR_66 = RG_rl_237 ;
	7'h36 :
		TR_66 = 9'h000 ;	// line#=../rle.cpp:68
	7'h37 :
		TR_66 = RG_rl_237 ;
	7'h38 :
		TR_66 = RG_rl_237 ;
	7'h39 :
		TR_66 = RG_rl_237 ;
	7'h3a :
		TR_66 = RG_rl_237 ;
	7'h3b :
		TR_66 = RG_rl_237 ;
	7'h3c :
		TR_66 = RG_rl_237 ;
	7'h3d :
		TR_66 = RG_rl_237 ;
	7'h3e :
		TR_66 = RG_rl_237 ;
	7'h3f :
		TR_66 = RG_rl_237 ;
	7'h40 :
		TR_66 = RG_rl_237 ;
	7'h41 :
		TR_66 = RG_rl_237 ;
	7'h42 :
		TR_66 = RG_rl_237 ;
	7'h43 :
		TR_66 = RG_rl_237 ;
	7'h44 :
		TR_66 = RG_rl_237 ;
	7'h45 :
		TR_66 = RG_rl_237 ;
	7'h46 :
		TR_66 = RG_rl_237 ;
	7'h47 :
		TR_66 = RG_rl_237 ;
	7'h48 :
		TR_66 = RG_rl_237 ;
	7'h49 :
		TR_66 = RG_rl_237 ;
	7'h4a :
		TR_66 = RG_rl_237 ;
	7'h4b :
		TR_66 = RG_rl_237 ;
	7'h4c :
		TR_66 = RG_rl_237 ;
	7'h4d :
		TR_66 = RG_rl_237 ;
	7'h4e :
		TR_66 = RG_rl_237 ;
	7'h4f :
		TR_66 = RG_rl_237 ;
	7'h50 :
		TR_66 = RG_rl_237 ;
	7'h51 :
		TR_66 = RG_rl_237 ;
	7'h52 :
		TR_66 = RG_rl_237 ;
	7'h53 :
		TR_66 = RG_rl_237 ;
	7'h54 :
		TR_66 = RG_rl_237 ;
	7'h55 :
		TR_66 = RG_rl_237 ;
	7'h56 :
		TR_66 = RG_rl_237 ;
	7'h57 :
		TR_66 = RG_rl_237 ;
	7'h58 :
		TR_66 = RG_rl_237 ;
	7'h59 :
		TR_66 = RG_rl_237 ;
	7'h5a :
		TR_66 = RG_rl_237 ;
	7'h5b :
		TR_66 = RG_rl_237 ;
	7'h5c :
		TR_66 = RG_rl_237 ;
	7'h5d :
		TR_66 = RG_rl_237 ;
	7'h5e :
		TR_66 = RG_rl_237 ;
	7'h5f :
		TR_66 = RG_rl_237 ;
	7'h60 :
		TR_66 = RG_rl_237 ;
	7'h61 :
		TR_66 = RG_rl_237 ;
	7'h62 :
		TR_66 = RG_rl_237 ;
	7'h63 :
		TR_66 = RG_rl_237 ;
	7'h64 :
		TR_66 = RG_rl_237 ;
	7'h65 :
		TR_66 = RG_rl_237 ;
	7'h66 :
		TR_66 = RG_rl_237 ;
	7'h67 :
		TR_66 = RG_rl_237 ;
	7'h68 :
		TR_66 = RG_rl_237 ;
	7'h69 :
		TR_66 = RG_rl_237 ;
	7'h6a :
		TR_66 = RG_rl_237 ;
	7'h6b :
		TR_66 = RG_rl_237 ;
	7'h6c :
		TR_66 = RG_rl_237 ;
	7'h6d :
		TR_66 = RG_rl_237 ;
	7'h6e :
		TR_66 = RG_rl_237 ;
	7'h6f :
		TR_66 = RG_rl_237 ;
	7'h70 :
		TR_66 = RG_rl_237 ;
	7'h71 :
		TR_66 = RG_rl_237 ;
	7'h72 :
		TR_66 = RG_rl_237 ;
	7'h73 :
		TR_66 = RG_rl_237 ;
	7'h74 :
		TR_66 = RG_rl_237 ;
	7'h75 :
		TR_66 = RG_rl_237 ;
	7'h76 :
		TR_66 = RG_rl_237 ;
	7'h77 :
		TR_66 = RG_rl_237 ;
	7'h78 :
		TR_66 = RG_rl_237 ;
	7'h79 :
		TR_66 = RG_rl_237 ;
	7'h7a :
		TR_66 = RG_rl_237 ;
	7'h7b :
		TR_66 = RG_rl_237 ;
	7'h7c :
		TR_66 = RG_rl_237 ;
	7'h7d :
		TR_66 = RG_rl_237 ;
	7'h7e :
		TR_66 = RG_rl_237 ;
	7'h7f :
		TR_66 = RG_rl_237 ;
	default :
		TR_66 = 9'hx ;
	endcase
always @ ( RG_rl_238 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_67 = RG_rl_238 ;
	7'h01 :
		TR_67 = RG_rl_238 ;
	7'h02 :
		TR_67 = RG_rl_238 ;
	7'h03 :
		TR_67 = RG_rl_238 ;
	7'h04 :
		TR_67 = RG_rl_238 ;
	7'h05 :
		TR_67 = RG_rl_238 ;
	7'h06 :
		TR_67 = RG_rl_238 ;
	7'h07 :
		TR_67 = RG_rl_238 ;
	7'h08 :
		TR_67 = RG_rl_238 ;
	7'h09 :
		TR_67 = RG_rl_238 ;
	7'h0a :
		TR_67 = RG_rl_238 ;
	7'h0b :
		TR_67 = RG_rl_238 ;
	7'h0c :
		TR_67 = RG_rl_238 ;
	7'h0d :
		TR_67 = RG_rl_238 ;
	7'h0e :
		TR_67 = RG_rl_238 ;
	7'h0f :
		TR_67 = RG_rl_238 ;
	7'h10 :
		TR_67 = RG_rl_238 ;
	7'h11 :
		TR_67 = RG_rl_238 ;
	7'h12 :
		TR_67 = RG_rl_238 ;
	7'h13 :
		TR_67 = RG_rl_238 ;
	7'h14 :
		TR_67 = RG_rl_238 ;
	7'h15 :
		TR_67 = RG_rl_238 ;
	7'h16 :
		TR_67 = RG_rl_238 ;
	7'h17 :
		TR_67 = RG_rl_238 ;
	7'h18 :
		TR_67 = RG_rl_238 ;
	7'h19 :
		TR_67 = RG_rl_238 ;
	7'h1a :
		TR_67 = RG_rl_238 ;
	7'h1b :
		TR_67 = RG_rl_238 ;
	7'h1c :
		TR_67 = RG_rl_238 ;
	7'h1d :
		TR_67 = RG_rl_238 ;
	7'h1e :
		TR_67 = RG_rl_238 ;
	7'h1f :
		TR_67 = RG_rl_238 ;
	7'h20 :
		TR_67 = RG_rl_238 ;
	7'h21 :
		TR_67 = RG_rl_238 ;
	7'h22 :
		TR_67 = RG_rl_238 ;
	7'h23 :
		TR_67 = RG_rl_238 ;
	7'h24 :
		TR_67 = RG_rl_238 ;
	7'h25 :
		TR_67 = RG_rl_238 ;
	7'h26 :
		TR_67 = RG_rl_238 ;
	7'h27 :
		TR_67 = RG_rl_238 ;
	7'h28 :
		TR_67 = RG_rl_238 ;
	7'h29 :
		TR_67 = RG_rl_238 ;
	7'h2a :
		TR_67 = RG_rl_238 ;
	7'h2b :
		TR_67 = RG_rl_238 ;
	7'h2c :
		TR_67 = RG_rl_238 ;
	7'h2d :
		TR_67 = RG_rl_238 ;
	7'h2e :
		TR_67 = RG_rl_238 ;
	7'h2f :
		TR_67 = RG_rl_238 ;
	7'h30 :
		TR_67 = RG_rl_238 ;
	7'h31 :
		TR_67 = RG_rl_238 ;
	7'h32 :
		TR_67 = RG_rl_238 ;
	7'h33 :
		TR_67 = RG_rl_238 ;
	7'h34 :
		TR_67 = RG_rl_238 ;
	7'h35 :
		TR_67 = RG_rl_238 ;
	7'h36 :
		TR_67 = RG_rl_238 ;
	7'h37 :
		TR_67 = 9'h000 ;	// line#=../rle.cpp:68
	7'h38 :
		TR_67 = RG_rl_238 ;
	7'h39 :
		TR_67 = RG_rl_238 ;
	7'h3a :
		TR_67 = RG_rl_238 ;
	7'h3b :
		TR_67 = RG_rl_238 ;
	7'h3c :
		TR_67 = RG_rl_238 ;
	7'h3d :
		TR_67 = RG_rl_238 ;
	7'h3e :
		TR_67 = RG_rl_238 ;
	7'h3f :
		TR_67 = RG_rl_238 ;
	7'h40 :
		TR_67 = RG_rl_238 ;
	7'h41 :
		TR_67 = RG_rl_238 ;
	7'h42 :
		TR_67 = RG_rl_238 ;
	7'h43 :
		TR_67 = RG_rl_238 ;
	7'h44 :
		TR_67 = RG_rl_238 ;
	7'h45 :
		TR_67 = RG_rl_238 ;
	7'h46 :
		TR_67 = RG_rl_238 ;
	7'h47 :
		TR_67 = RG_rl_238 ;
	7'h48 :
		TR_67 = RG_rl_238 ;
	7'h49 :
		TR_67 = RG_rl_238 ;
	7'h4a :
		TR_67 = RG_rl_238 ;
	7'h4b :
		TR_67 = RG_rl_238 ;
	7'h4c :
		TR_67 = RG_rl_238 ;
	7'h4d :
		TR_67 = RG_rl_238 ;
	7'h4e :
		TR_67 = RG_rl_238 ;
	7'h4f :
		TR_67 = RG_rl_238 ;
	7'h50 :
		TR_67 = RG_rl_238 ;
	7'h51 :
		TR_67 = RG_rl_238 ;
	7'h52 :
		TR_67 = RG_rl_238 ;
	7'h53 :
		TR_67 = RG_rl_238 ;
	7'h54 :
		TR_67 = RG_rl_238 ;
	7'h55 :
		TR_67 = RG_rl_238 ;
	7'h56 :
		TR_67 = RG_rl_238 ;
	7'h57 :
		TR_67 = RG_rl_238 ;
	7'h58 :
		TR_67 = RG_rl_238 ;
	7'h59 :
		TR_67 = RG_rl_238 ;
	7'h5a :
		TR_67 = RG_rl_238 ;
	7'h5b :
		TR_67 = RG_rl_238 ;
	7'h5c :
		TR_67 = RG_rl_238 ;
	7'h5d :
		TR_67 = RG_rl_238 ;
	7'h5e :
		TR_67 = RG_rl_238 ;
	7'h5f :
		TR_67 = RG_rl_238 ;
	7'h60 :
		TR_67 = RG_rl_238 ;
	7'h61 :
		TR_67 = RG_rl_238 ;
	7'h62 :
		TR_67 = RG_rl_238 ;
	7'h63 :
		TR_67 = RG_rl_238 ;
	7'h64 :
		TR_67 = RG_rl_238 ;
	7'h65 :
		TR_67 = RG_rl_238 ;
	7'h66 :
		TR_67 = RG_rl_238 ;
	7'h67 :
		TR_67 = RG_rl_238 ;
	7'h68 :
		TR_67 = RG_rl_238 ;
	7'h69 :
		TR_67 = RG_rl_238 ;
	7'h6a :
		TR_67 = RG_rl_238 ;
	7'h6b :
		TR_67 = RG_rl_238 ;
	7'h6c :
		TR_67 = RG_rl_238 ;
	7'h6d :
		TR_67 = RG_rl_238 ;
	7'h6e :
		TR_67 = RG_rl_238 ;
	7'h6f :
		TR_67 = RG_rl_238 ;
	7'h70 :
		TR_67 = RG_rl_238 ;
	7'h71 :
		TR_67 = RG_rl_238 ;
	7'h72 :
		TR_67 = RG_rl_238 ;
	7'h73 :
		TR_67 = RG_rl_238 ;
	7'h74 :
		TR_67 = RG_rl_238 ;
	7'h75 :
		TR_67 = RG_rl_238 ;
	7'h76 :
		TR_67 = RG_rl_238 ;
	7'h77 :
		TR_67 = RG_rl_238 ;
	7'h78 :
		TR_67 = RG_rl_238 ;
	7'h79 :
		TR_67 = RG_rl_238 ;
	7'h7a :
		TR_67 = RG_rl_238 ;
	7'h7b :
		TR_67 = RG_rl_238 ;
	7'h7c :
		TR_67 = RG_rl_238 ;
	7'h7d :
		TR_67 = RG_rl_238 ;
	7'h7e :
		TR_67 = RG_rl_238 ;
	7'h7f :
		TR_67 = RG_rl_238 ;
	default :
		TR_67 = 9'hx ;
	endcase
always @ ( RG_rl_239 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_68 = RG_rl_239 ;
	7'h01 :
		TR_68 = RG_rl_239 ;
	7'h02 :
		TR_68 = RG_rl_239 ;
	7'h03 :
		TR_68 = RG_rl_239 ;
	7'h04 :
		TR_68 = RG_rl_239 ;
	7'h05 :
		TR_68 = RG_rl_239 ;
	7'h06 :
		TR_68 = RG_rl_239 ;
	7'h07 :
		TR_68 = RG_rl_239 ;
	7'h08 :
		TR_68 = RG_rl_239 ;
	7'h09 :
		TR_68 = RG_rl_239 ;
	7'h0a :
		TR_68 = RG_rl_239 ;
	7'h0b :
		TR_68 = RG_rl_239 ;
	7'h0c :
		TR_68 = RG_rl_239 ;
	7'h0d :
		TR_68 = RG_rl_239 ;
	7'h0e :
		TR_68 = RG_rl_239 ;
	7'h0f :
		TR_68 = RG_rl_239 ;
	7'h10 :
		TR_68 = RG_rl_239 ;
	7'h11 :
		TR_68 = RG_rl_239 ;
	7'h12 :
		TR_68 = RG_rl_239 ;
	7'h13 :
		TR_68 = RG_rl_239 ;
	7'h14 :
		TR_68 = RG_rl_239 ;
	7'h15 :
		TR_68 = RG_rl_239 ;
	7'h16 :
		TR_68 = RG_rl_239 ;
	7'h17 :
		TR_68 = RG_rl_239 ;
	7'h18 :
		TR_68 = RG_rl_239 ;
	7'h19 :
		TR_68 = RG_rl_239 ;
	7'h1a :
		TR_68 = RG_rl_239 ;
	7'h1b :
		TR_68 = RG_rl_239 ;
	7'h1c :
		TR_68 = RG_rl_239 ;
	7'h1d :
		TR_68 = RG_rl_239 ;
	7'h1e :
		TR_68 = RG_rl_239 ;
	7'h1f :
		TR_68 = RG_rl_239 ;
	7'h20 :
		TR_68 = RG_rl_239 ;
	7'h21 :
		TR_68 = RG_rl_239 ;
	7'h22 :
		TR_68 = RG_rl_239 ;
	7'h23 :
		TR_68 = RG_rl_239 ;
	7'h24 :
		TR_68 = RG_rl_239 ;
	7'h25 :
		TR_68 = RG_rl_239 ;
	7'h26 :
		TR_68 = RG_rl_239 ;
	7'h27 :
		TR_68 = RG_rl_239 ;
	7'h28 :
		TR_68 = RG_rl_239 ;
	7'h29 :
		TR_68 = RG_rl_239 ;
	7'h2a :
		TR_68 = RG_rl_239 ;
	7'h2b :
		TR_68 = RG_rl_239 ;
	7'h2c :
		TR_68 = RG_rl_239 ;
	7'h2d :
		TR_68 = RG_rl_239 ;
	7'h2e :
		TR_68 = RG_rl_239 ;
	7'h2f :
		TR_68 = RG_rl_239 ;
	7'h30 :
		TR_68 = RG_rl_239 ;
	7'h31 :
		TR_68 = RG_rl_239 ;
	7'h32 :
		TR_68 = RG_rl_239 ;
	7'h33 :
		TR_68 = RG_rl_239 ;
	7'h34 :
		TR_68 = RG_rl_239 ;
	7'h35 :
		TR_68 = RG_rl_239 ;
	7'h36 :
		TR_68 = RG_rl_239 ;
	7'h37 :
		TR_68 = RG_rl_239 ;
	7'h38 :
		TR_68 = 9'h000 ;	// line#=../rle.cpp:68
	7'h39 :
		TR_68 = RG_rl_239 ;
	7'h3a :
		TR_68 = RG_rl_239 ;
	7'h3b :
		TR_68 = RG_rl_239 ;
	7'h3c :
		TR_68 = RG_rl_239 ;
	7'h3d :
		TR_68 = RG_rl_239 ;
	7'h3e :
		TR_68 = RG_rl_239 ;
	7'h3f :
		TR_68 = RG_rl_239 ;
	7'h40 :
		TR_68 = RG_rl_239 ;
	7'h41 :
		TR_68 = RG_rl_239 ;
	7'h42 :
		TR_68 = RG_rl_239 ;
	7'h43 :
		TR_68 = RG_rl_239 ;
	7'h44 :
		TR_68 = RG_rl_239 ;
	7'h45 :
		TR_68 = RG_rl_239 ;
	7'h46 :
		TR_68 = RG_rl_239 ;
	7'h47 :
		TR_68 = RG_rl_239 ;
	7'h48 :
		TR_68 = RG_rl_239 ;
	7'h49 :
		TR_68 = RG_rl_239 ;
	7'h4a :
		TR_68 = RG_rl_239 ;
	7'h4b :
		TR_68 = RG_rl_239 ;
	7'h4c :
		TR_68 = RG_rl_239 ;
	7'h4d :
		TR_68 = RG_rl_239 ;
	7'h4e :
		TR_68 = RG_rl_239 ;
	7'h4f :
		TR_68 = RG_rl_239 ;
	7'h50 :
		TR_68 = RG_rl_239 ;
	7'h51 :
		TR_68 = RG_rl_239 ;
	7'h52 :
		TR_68 = RG_rl_239 ;
	7'h53 :
		TR_68 = RG_rl_239 ;
	7'h54 :
		TR_68 = RG_rl_239 ;
	7'h55 :
		TR_68 = RG_rl_239 ;
	7'h56 :
		TR_68 = RG_rl_239 ;
	7'h57 :
		TR_68 = RG_rl_239 ;
	7'h58 :
		TR_68 = RG_rl_239 ;
	7'h59 :
		TR_68 = RG_rl_239 ;
	7'h5a :
		TR_68 = RG_rl_239 ;
	7'h5b :
		TR_68 = RG_rl_239 ;
	7'h5c :
		TR_68 = RG_rl_239 ;
	7'h5d :
		TR_68 = RG_rl_239 ;
	7'h5e :
		TR_68 = RG_rl_239 ;
	7'h5f :
		TR_68 = RG_rl_239 ;
	7'h60 :
		TR_68 = RG_rl_239 ;
	7'h61 :
		TR_68 = RG_rl_239 ;
	7'h62 :
		TR_68 = RG_rl_239 ;
	7'h63 :
		TR_68 = RG_rl_239 ;
	7'h64 :
		TR_68 = RG_rl_239 ;
	7'h65 :
		TR_68 = RG_rl_239 ;
	7'h66 :
		TR_68 = RG_rl_239 ;
	7'h67 :
		TR_68 = RG_rl_239 ;
	7'h68 :
		TR_68 = RG_rl_239 ;
	7'h69 :
		TR_68 = RG_rl_239 ;
	7'h6a :
		TR_68 = RG_rl_239 ;
	7'h6b :
		TR_68 = RG_rl_239 ;
	7'h6c :
		TR_68 = RG_rl_239 ;
	7'h6d :
		TR_68 = RG_rl_239 ;
	7'h6e :
		TR_68 = RG_rl_239 ;
	7'h6f :
		TR_68 = RG_rl_239 ;
	7'h70 :
		TR_68 = RG_rl_239 ;
	7'h71 :
		TR_68 = RG_rl_239 ;
	7'h72 :
		TR_68 = RG_rl_239 ;
	7'h73 :
		TR_68 = RG_rl_239 ;
	7'h74 :
		TR_68 = RG_rl_239 ;
	7'h75 :
		TR_68 = RG_rl_239 ;
	7'h76 :
		TR_68 = RG_rl_239 ;
	7'h77 :
		TR_68 = RG_rl_239 ;
	7'h78 :
		TR_68 = RG_rl_239 ;
	7'h79 :
		TR_68 = RG_rl_239 ;
	7'h7a :
		TR_68 = RG_rl_239 ;
	7'h7b :
		TR_68 = RG_rl_239 ;
	7'h7c :
		TR_68 = RG_rl_239 ;
	7'h7d :
		TR_68 = RG_rl_239 ;
	7'h7e :
		TR_68 = RG_rl_239 ;
	7'h7f :
		TR_68 = RG_rl_239 ;
	default :
		TR_68 = 9'hx ;
	endcase
always @ ( RG_rl_240 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_69 = RG_rl_240 ;
	7'h01 :
		TR_69 = RG_rl_240 ;
	7'h02 :
		TR_69 = RG_rl_240 ;
	7'h03 :
		TR_69 = RG_rl_240 ;
	7'h04 :
		TR_69 = RG_rl_240 ;
	7'h05 :
		TR_69 = RG_rl_240 ;
	7'h06 :
		TR_69 = RG_rl_240 ;
	7'h07 :
		TR_69 = RG_rl_240 ;
	7'h08 :
		TR_69 = RG_rl_240 ;
	7'h09 :
		TR_69 = RG_rl_240 ;
	7'h0a :
		TR_69 = RG_rl_240 ;
	7'h0b :
		TR_69 = RG_rl_240 ;
	7'h0c :
		TR_69 = RG_rl_240 ;
	7'h0d :
		TR_69 = RG_rl_240 ;
	7'h0e :
		TR_69 = RG_rl_240 ;
	7'h0f :
		TR_69 = RG_rl_240 ;
	7'h10 :
		TR_69 = RG_rl_240 ;
	7'h11 :
		TR_69 = RG_rl_240 ;
	7'h12 :
		TR_69 = RG_rl_240 ;
	7'h13 :
		TR_69 = RG_rl_240 ;
	7'h14 :
		TR_69 = RG_rl_240 ;
	7'h15 :
		TR_69 = RG_rl_240 ;
	7'h16 :
		TR_69 = RG_rl_240 ;
	7'h17 :
		TR_69 = RG_rl_240 ;
	7'h18 :
		TR_69 = RG_rl_240 ;
	7'h19 :
		TR_69 = RG_rl_240 ;
	7'h1a :
		TR_69 = RG_rl_240 ;
	7'h1b :
		TR_69 = RG_rl_240 ;
	7'h1c :
		TR_69 = RG_rl_240 ;
	7'h1d :
		TR_69 = RG_rl_240 ;
	7'h1e :
		TR_69 = RG_rl_240 ;
	7'h1f :
		TR_69 = RG_rl_240 ;
	7'h20 :
		TR_69 = RG_rl_240 ;
	7'h21 :
		TR_69 = RG_rl_240 ;
	7'h22 :
		TR_69 = RG_rl_240 ;
	7'h23 :
		TR_69 = RG_rl_240 ;
	7'h24 :
		TR_69 = RG_rl_240 ;
	7'h25 :
		TR_69 = RG_rl_240 ;
	7'h26 :
		TR_69 = RG_rl_240 ;
	7'h27 :
		TR_69 = RG_rl_240 ;
	7'h28 :
		TR_69 = RG_rl_240 ;
	7'h29 :
		TR_69 = RG_rl_240 ;
	7'h2a :
		TR_69 = RG_rl_240 ;
	7'h2b :
		TR_69 = RG_rl_240 ;
	7'h2c :
		TR_69 = RG_rl_240 ;
	7'h2d :
		TR_69 = RG_rl_240 ;
	7'h2e :
		TR_69 = RG_rl_240 ;
	7'h2f :
		TR_69 = RG_rl_240 ;
	7'h30 :
		TR_69 = RG_rl_240 ;
	7'h31 :
		TR_69 = RG_rl_240 ;
	7'h32 :
		TR_69 = RG_rl_240 ;
	7'h33 :
		TR_69 = RG_rl_240 ;
	7'h34 :
		TR_69 = RG_rl_240 ;
	7'h35 :
		TR_69 = RG_rl_240 ;
	7'h36 :
		TR_69 = RG_rl_240 ;
	7'h37 :
		TR_69 = RG_rl_240 ;
	7'h38 :
		TR_69 = RG_rl_240 ;
	7'h39 :
		TR_69 = 9'h000 ;	// line#=../rle.cpp:68
	7'h3a :
		TR_69 = RG_rl_240 ;
	7'h3b :
		TR_69 = RG_rl_240 ;
	7'h3c :
		TR_69 = RG_rl_240 ;
	7'h3d :
		TR_69 = RG_rl_240 ;
	7'h3e :
		TR_69 = RG_rl_240 ;
	7'h3f :
		TR_69 = RG_rl_240 ;
	7'h40 :
		TR_69 = RG_rl_240 ;
	7'h41 :
		TR_69 = RG_rl_240 ;
	7'h42 :
		TR_69 = RG_rl_240 ;
	7'h43 :
		TR_69 = RG_rl_240 ;
	7'h44 :
		TR_69 = RG_rl_240 ;
	7'h45 :
		TR_69 = RG_rl_240 ;
	7'h46 :
		TR_69 = RG_rl_240 ;
	7'h47 :
		TR_69 = RG_rl_240 ;
	7'h48 :
		TR_69 = RG_rl_240 ;
	7'h49 :
		TR_69 = RG_rl_240 ;
	7'h4a :
		TR_69 = RG_rl_240 ;
	7'h4b :
		TR_69 = RG_rl_240 ;
	7'h4c :
		TR_69 = RG_rl_240 ;
	7'h4d :
		TR_69 = RG_rl_240 ;
	7'h4e :
		TR_69 = RG_rl_240 ;
	7'h4f :
		TR_69 = RG_rl_240 ;
	7'h50 :
		TR_69 = RG_rl_240 ;
	7'h51 :
		TR_69 = RG_rl_240 ;
	7'h52 :
		TR_69 = RG_rl_240 ;
	7'h53 :
		TR_69 = RG_rl_240 ;
	7'h54 :
		TR_69 = RG_rl_240 ;
	7'h55 :
		TR_69 = RG_rl_240 ;
	7'h56 :
		TR_69 = RG_rl_240 ;
	7'h57 :
		TR_69 = RG_rl_240 ;
	7'h58 :
		TR_69 = RG_rl_240 ;
	7'h59 :
		TR_69 = RG_rl_240 ;
	7'h5a :
		TR_69 = RG_rl_240 ;
	7'h5b :
		TR_69 = RG_rl_240 ;
	7'h5c :
		TR_69 = RG_rl_240 ;
	7'h5d :
		TR_69 = RG_rl_240 ;
	7'h5e :
		TR_69 = RG_rl_240 ;
	7'h5f :
		TR_69 = RG_rl_240 ;
	7'h60 :
		TR_69 = RG_rl_240 ;
	7'h61 :
		TR_69 = RG_rl_240 ;
	7'h62 :
		TR_69 = RG_rl_240 ;
	7'h63 :
		TR_69 = RG_rl_240 ;
	7'h64 :
		TR_69 = RG_rl_240 ;
	7'h65 :
		TR_69 = RG_rl_240 ;
	7'h66 :
		TR_69 = RG_rl_240 ;
	7'h67 :
		TR_69 = RG_rl_240 ;
	7'h68 :
		TR_69 = RG_rl_240 ;
	7'h69 :
		TR_69 = RG_rl_240 ;
	7'h6a :
		TR_69 = RG_rl_240 ;
	7'h6b :
		TR_69 = RG_rl_240 ;
	7'h6c :
		TR_69 = RG_rl_240 ;
	7'h6d :
		TR_69 = RG_rl_240 ;
	7'h6e :
		TR_69 = RG_rl_240 ;
	7'h6f :
		TR_69 = RG_rl_240 ;
	7'h70 :
		TR_69 = RG_rl_240 ;
	7'h71 :
		TR_69 = RG_rl_240 ;
	7'h72 :
		TR_69 = RG_rl_240 ;
	7'h73 :
		TR_69 = RG_rl_240 ;
	7'h74 :
		TR_69 = RG_rl_240 ;
	7'h75 :
		TR_69 = RG_rl_240 ;
	7'h76 :
		TR_69 = RG_rl_240 ;
	7'h77 :
		TR_69 = RG_rl_240 ;
	7'h78 :
		TR_69 = RG_rl_240 ;
	7'h79 :
		TR_69 = RG_rl_240 ;
	7'h7a :
		TR_69 = RG_rl_240 ;
	7'h7b :
		TR_69 = RG_rl_240 ;
	7'h7c :
		TR_69 = RG_rl_240 ;
	7'h7d :
		TR_69 = RG_rl_240 ;
	7'h7e :
		TR_69 = RG_rl_240 ;
	7'h7f :
		TR_69 = RG_rl_240 ;
	default :
		TR_69 = 9'hx ;
	endcase
always @ ( RG_rl_241 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_70 = RG_rl_241 ;
	7'h01 :
		TR_70 = RG_rl_241 ;
	7'h02 :
		TR_70 = RG_rl_241 ;
	7'h03 :
		TR_70 = RG_rl_241 ;
	7'h04 :
		TR_70 = RG_rl_241 ;
	7'h05 :
		TR_70 = RG_rl_241 ;
	7'h06 :
		TR_70 = RG_rl_241 ;
	7'h07 :
		TR_70 = RG_rl_241 ;
	7'h08 :
		TR_70 = RG_rl_241 ;
	7'h09 :
		TR_70 = RG_rl_241 ;
	7'h0a :
		TR_70 = RG_rl_241 ;
	7'h0b :
		TR_70 = RG_rl_241 ;
	7'h0c :
		TR_70 = RG_rl_241 ;
	7'h0d :
		TR_70 = RG_rl_241 ;
	7'h0e :
		TR_70 = RG_rl_241 ;
	7'h0f :
		TR_70 = RG_rl_241 ;
	7'h10 :
		TR_70 = RG_rl_241 ;
	7'h11 :
		TR_70 = RG_rl_241 ;
	7'h12 :
		TR_70 = RG_rl_241 ;
	7'h13 :
		TR_70 = RG_rl_241 ;
	7'h14 :
		TR_70 = RG_rl_241 ;
	7'h15 :
		TR_70 = RG_rl_241 ;
	7'h16 :
		TR_70 = RG_rl_241 ;
	7'h17 :
		TR_70 = RG_rl_241 ;
	7'h18 :
		TR_70 = RG_rl_241 ;
	7'h19 :
		TR_70 = RG_rl_241 ;
	7'h1a :
		TR_70 = RG_rl_241 ;
	7'h1b :
		TR_70 = RG_rl_241 ;
	7'h1c :
		TR_70 = RG_rl_241 ;
	7'h1d :
		TR_70 = RG_rl_241 ;
	7'h1e :
		TR_70 = RG_rl_241 ;
	7'h1f :
		TR_70 = RG_rl_241 ;
	7'h20 :
		TR_70 = RG_rl_241 ;
	7'h21 :
		TR_70 = RG_rl_241 ;
	7'h22 :
		TR_70 = RG_rl_241 ;
	7'h23 :
		TR_70 = RG_rl_241 ;
	7'h24 :
		TR_70 = RG_rl_241 ;
	7'h25 :
		TR_70 = RG_rl_241 ;
	7'h26 :
		TR_70 = RG_rl_241 ;
	7'h27 :
		TR_70 = RG_rl_241 ;
	7'h28 :
		TR_70 = RG_rl_241 ;
	7'h29 :
		TR_70 = RG_rl_241 ;
	7'h2a :
		TR_70 = RG_rl_241 ;
	7'h2b :
		TR_70 = RG_rl_241 ;
	7'h2c :
		TR_70 = RG_rl_241 ;
	7'h2d :
		TR_70 = RG_rl_241 ;
	7'h2e :
		TR_70 = RG_rl_241 ;
	7'h2f :
		TR_70 = RG_rl_241 ;
	7'h30 :
		TR_70 = RG_rl_241 ;
	7'h31 :
		TR_70 = RG_rl_241 ;
	7'h32 :
		TR_70 = RG_rl_241 ;
	7'h33 :
		TR_70 = RG_rl_241 ;
	7'h34 :
		TR_70 = RG_rl_241 ;
	7'h35 :
		TR_70 = RG_rl_241 ;
	7'h36 :
		TR_70 = RG_rl_241 ;
	7'h37 :
		TR_70 = RG_rl_241 ;
	7'h38 :
		TR_70 = RG_rl_241 ;
	7'h39 :
		TR_70 = RG_rl_241 ;
	7'h3a :
		TR_70 = 9'h000 ;	// line#=../rle.cpp:68
	7'h3b :
		TR_70 = RG_rl_241 ;
	7'h3c :
		TR_70 = RG_rl_241 ;
	7'h3d :
		TR_70 = RG_rl_241 ;
	7'h3e :
		TR_70 = RG_rl_241 ;
	7'h3f :
		TR_70 = RG_rl_241 ;
	7'h40 :
		TR_70 = RG_rl_241 ;
	7'h41 :
		TR_70 = RG_rl_241 ;
	7'h42 :
		TR_70 = RG_rl_241 ;
	7'h43 :
		TR_70 = RG_rl_241 ;
	7'h44 :
		TR_70 = RG_rl_241 ;
	7'h45 :
		TR_70 = RG_rl_241 ;
	7'h46 :
		TR_70 = RG_rl_241 ;
	7'h47 :
		TR_70 = RG_rl_241 ;
	7'h48 :
		TR_70 = RG_rl_241 ;
	7'h49 :
		TR_70 = RG_rl_241 ;
	7'h4a :
		TR_70 = RG_rl_241 ;
	7'h4b :
		TR_70 = RG_rl_241 ;
	7'h4c :
		TR_70 = RG_rl_241 ;
	7'h4d :
		TR_70 = RG_rl_241 ;
	7'h4e :
		TR_70 = RG_rl_241 ;
	7'h4f :
		TR_70 = RG_rl_241 ;
	7'h50 :
		TR_70 = RG_rl_241 ;
	7'h51 :
		TR_70 = RG_rl_241 ;
	7'h52 :
		TR_70 = RG_rl_241 ;
	7'h53 :
		TR_70 = RG_rl_241 ;
	7'h54 :
		TR_70 = RG_rl_241 ;
	7'h55 :
		TR_70 = RG_rl_241 ;
	7'h56 :
		TR_70 = RG_rl_241 ;
	7'h57 :
		TR_70 = RG_rl_241 ;
	7'h58 :
		TR_70 = RG_rl_241 ;
	7'h59 :
		TR_70 = RG_rl_241 ;
	7'h5a :
		TR_70 = RG_rl_241 ;
	7'h5b :
		TR_70 = RG_rl_241 ;
	7'h5c :
		TR_70 = RG_rl_241 ;
	7'h5d :
		TR_70 = RG_rl_241 ;
	7'h5e :
		TR_70 = RG_rl_241 ;
	7'h5f :
		TR_70 = RG_rl_241 ;
	7'h60 :
		TR_70 = RG_rl_241 ;
	7'h61 :
		TR_70 = RG_rl_241 ;
	7'h62 :
		TR_70 = RG_rl_241 ;
	7'h63 :
		TR_70 = RG_rl_241 ;
	7'h64 :
		TR_70 = RG_rl_241 ;
	7'h65 :
		TR_70 = RG_rl_241 ;
	7'h66 :
		TR_70 = RG_rl_241 ;
	7'h67 :
		TR_70 = RG_rl_241 ;
	7'h68 :
		TR_70 = RG_rl_241 ;
	7'h69 :
		TR_70 = RG_rl_241 ;
	7'h6a :
		TR_70 = RG_rl_241 ;
	7'h6b :
		TR_70 = RG_rl_241 ;
	7'h6c :
		TR_70 = RG_rl_241 ;
	7'h6d :
		TR_70 = RG_rl_241 ;
	7'h6e :
		TR_70 = RG_rl_241 ;
	7'h6f :
		TR_70 = RG_rl_241 ;
	7'h70 :
		TR_70 = RG_rl_241 ;
	7'h71 :
		TR_70 = RG_rl_241 ;
	7'h72 :
		TR_70 = RG_rl_241 ;
	7'h73 :
		TR_70 = RG_rl_241 ;
	7'h74 :
		TR_70 = RG_rl_241 ;
	7'h75 :
		TR_70 = RG_rl_241 ;
	7'h76 :
		TR_70 = RG_rl_241 ;
	7'h77 :
		TR_70 = RG_rl_241 ;
	7'h78 :
		TR_70 = RG_rl_241 ;
	7'h79 :
		TR_70 = RG_rl_241 ;
	7'h7a :
		TR_70 = RG_rl_241 ;
	7'h7b :
		TR_70 = RG_rl_241 ;
	7'h7c :
		TR_70 = RG_rl_241 ;
	7'h7d :
		TR_70 = RG_rl_241 ;
	7'h7e :
		TR_70 = RG_rl_241 ;
	7'h7f :
		TR_70 = RG_rl_241 ;
	default :
		TR_70 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_71 = RG_quantized_block_rl ;
	7'h01 :
		TR_71 = RG_quantized_block_rl ;
	7'h02 :
		TR_71 = RG_quantized_block_rl ;
	7'h03 :
		TR_71 = RG_quantized_block_rl ;
	7'h04 :
		TR_71 = RG_quantized_block_rl ;
	7'h05 :
		TR_71 = RG_quantized_block_rl ;
	7'h06 :
		TR_71 = RG_quantized_block_rl ;
	7'h07 :
		TR_71 = RG_quantized_block_rl ;
	7'h08 :
		TR_71 = RG_quantized_block_rl ;
	7'h09 :
		TR_71 = RG_quantized_block_rl ;
	7'h0a :
		TR_71 = RG_quantized_block_rl ;
	7'h0b :
		TR_71 = RG_quantized_block_rl ;
	7'h0c :
		TR_71 = RG_quantized_block_rl ;
	7'h0d :
		TR_71 = RG_quantized_block_rl ;
	7'h0e :
		TR_71 = RG_quantized_block_rl ;
	7'h0f :
		TR_71 = RG_quantized_block_rl ;
	7'h10 :
		TR_71 = RG_quantized_block_rl ;
	7'h11 :
		TR_71 = RG_quantized_block_rl ;
	7'h12 :
		TR_71 = RG_quantized_block_rl ;
	7'h13 :
		TR_71 = RG_quantized_block_rl ;
	7'h14 :
		TR_71 = RG_quantized_block_rl ;
	7'h15 :
		TR_71 = RG_quantized_block_rl ;
	7'h16 :
		TR_71 = RG_quantized_block_rl ;
	7'h17 :
		TR_71 = RG_quantized_block_rl ;
	7'h18 :
		TR_71 = RG_quantized_block_rl ;
	7'h19 :
		TR_71 = RG_quantized_block_rl ;
	7'h1a :
		TR_71 = RG_quantized_block_rl ;
	7'h1b :
		TR_71 = RG_quantized_block_rl ;
	7'h1c :
		TR_71 = RG_quantized_block_rl ;
	7'h1d :
		TR_71 = RG_quantized_block_rl ;
	7'h1e :
		TR_71 = RG_quantized_block_rl ;
	7'h1f :
		TR_71 = RG_quantized_block_rl ;
	7'h20 :
		TR_71 = RG_quantized_block_rl ;
	7'h21 :
		TR_71 = RG_quantized_block_rl ;
	7'h22 :
		TR_71 = RG_quantized_block_rl ;
	7'h23 :
		TR_71 = RG_quantized_block_rl ;
	7'h24 :
		TR_71 = RG_quantized_block_rl ;
	7'h25 :
		TR_71 = RG_quantized_block_rl ;
	7'h26 :
		TR_71 = RG_quantized_block_rl ;
	7'h27 :
		TR_71 = RG_quantized_block_rl ;
	7'h28 :
		TR_71 = RG_quantized_block_rl ;
	7'h29 :
		TR_71 = RG_quantized_block_rl ;
	7'h2a :
		TR_71 = RG_quantized_block_rl ;
	7'h2b :
		TR_71 = RG_quantized_block_rl ;
	7'h2c :
		TR_71 = RG_quantized_block_rl ;
	7'h2d :
		TR_71 = RG_quantized_block_rl ;
	7'h2e :
		TR_71 = RG_quantized_block_rl ;
	7'h2f :
		TR_71 = RG_quantized_block_rl ;
	7'h30 :
		TR_71 = RG_quantized_block_rl ;
	7'h31 :
		TR_71 = RG_quantized_block_rl ;
	7'h32 :
		TR_71 = RG_quantized_block_rl ;
	7'h33 :
		TR_71 = RG_quantized_block_rl ;
	7'h34 :
		TR_71 = RG_quantized_block_rl ;
	7'h35 :
		TR_71 = RG_quantized_block_rl ;
	7'h36 :
		TR_71 = RG_quantized_block_rl ;
	7'h37 :
		TR_71 = RG_quantized_block_rl ;
	7'h38 :
		TR_71 = RG_quantized_block_rl ;
	7'h39 :
		TR_71 = RG_quantized_block_rl ;
	7'h3a :
		TR_71 = RG_quantized_block_rl ;
	7'h3b :
		TR_71 = 9'h000 ;	// line#=../rle.cpp:68
	7'h3c :
		TR_71 = RG_quantized_block_rl ;
	7'h3d :
		TR_71 = RG_quantized_block_rl ;
	7'h3e :
		TR_71 = RG_quantized_block_rl ;
	7'h3f :
		TR_71 = RG_quantized_block_rl ;
	7'h40 :
		TR_71 = RG_quantized_block_rl ;
	7'h41 :
		TR_71 = RG_quantized_block_rl ;
	7'h42 :
		TR_71 = RG_quantized_block_rl ;
	7'h43 :
		TR_71 = RG_quantized_block_rl ;
	7'h44 :
		TR_71 = RG_quantized_block_rl ;
	7'h45 :
		TR_71 = RG_quantized_block_rl ;
	7'h46 :
		TR_71 = RG_quantized_block_rl ;
	7'h47 :
		TR_71 = RG_quantized_block_rl ;
	7'h48 :
		TR_71 = RG_quantized_block_rl ;
	7'h49 :
		TR_71 = RG_quantized_block_rl ;
	7'h4a :
		TR_71 = RG_quantized_block_rl ;
	7'h4b :
		TR_71 = RG_quantized_block_rl ;
	7'h4c :
		TR_71 = RG_quantized_block_rl ;
	7'h4d :
		TR_71 = RG_quantized_block_rl ;
	7'h4e :
		TR_71 = RG_quantized_block_rl ;
	7'h4f :
		TR_71 = RG_quantized_block_rl ;
	7'h50 :
		TR_71 = RG_quantized_block_rl ;
	7'h51 :
		TR_71 = RG_quantized_block_rl ;
	7'h52 :
		TR_71 = RG_quantized_block_rl ;
	7'h53 :
		TR_71 = RG_quantized_block_rl ;
	7'h54 :
		TR_71 = RG_quantized_block_rl ;
	7'h55 :
		TR_71 = RG_quantized_block_rl ;
	7'h56 :
		TR_71 = RG_quantized_block_rl ;
	7'h57 :
		TR_71 = RG_quantized_block_rl ;
	7'h58 :
		TR_71 = RG_quantized_block_rl ;
	7'h59 :
		TR_71 = RG_quantized_block_rl ;
	7'h5a :
		TR_71 = RG_quantized_block_rl ;
	7'h5b :
		TR_71 = RG_quantized_block_rl ;
	7'h5c :
		TR_71 = RG_quantized_block_rl ;
	7'h5d :
		TR_71 = RG_quantized_block_rl ;
	7'h5e :
		TR_71 = RG_quantized_block_rl ;
	7'h5f :
		TR_71 = RG_quantized_block_rl ;
	7'h60 :
		TR_71 = RG_quantized_block_rl ;
	7'h61 :
		TR_71 = RG_quantized_block_rl ;
	7'h62 :
		TR_71 = RG_quantized_block_rl ;
	7'h63 :
		TR_71 = RG_quantized_block_rl ;
	7'h64 :
		TR_71 = RG_quantized_block_rl ;
	7'h65 :
		TR_71 = RG_quantized_block_rl ;
	7'h66 :
		TR_71 = RG_quantized_block_rl ;
	7'h67 :
		TR_71 = RG_quantized_block_rl ;
	7'h68 :
		TR_71 = RG_quantized_block_rl ;
	7'h69 :
		TR_71 = RG_quantized_block_rl ;
	7'h6a :
		TR_71 = RG_quantized_block_rl ;
	7'h6b :
		TR_71 = RG_quantized_block_rl ;
	7'h6c :
		TR_71 = RG_quantized_block_rl ;
	7'h6d :
		TR_71 = RG_quantized_block_rl ;
	7'h6e :
		TR_71 = RG_quantized_block_rl ;
	7'h6f :
		TR_71 = RG_quantized_block_rl ;
	7'h70 :
		TR_71 = RG_quantized_block_rl ;
	7'h71 :
		TR_71 = RG_quantized_block_rl ;
	7'h72 :
		TR_71 = RG_quantized_block_rl ;
	7'h73 :
		TR_71 = RG_quantized_block_rl ;
	7'h74 :
		TR_71 = RG_quantized_block_rl ;
	7'h75 :
		TR_71 = RG_quantized_block_rl ;
	7'h76 :
		TR_71 = RG_quantized_block_rl ;
	7'h77 :
		TR_71 = RG_quantized_block_rl ;
	7'h78 :
		TR_71 = RG_quantized_block_rl ;
	7'h79 :
		TR_71 = RG_quantized_block_rl ;
	7'h7a :
		TR_71 = RG_quantized_block_rl ;
	7'h7b :
		TR_71 = RG_quantized_block_rl ;
	7'h7c :
		TR_71 = RG_quantized_block_rl ;
	7'h7d :
		TR_71 = RG_quantized_block_rl ;
	7'h7e :
		TR_71 = RG_quantized_block_rl ;
	7'h7f :
		TR_71 = RG_quantized_block_rl ;
	default :
		TR_71 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_1 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h01 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h02 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h03 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h04 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h05 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h06 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h07 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h08 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h09 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h0a :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h0b :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h0c :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h0d :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h0e :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h0f :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h10 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h11 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h12 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h13 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h14 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h15 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h16 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h17 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h18 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h19 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h1a :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h1b :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h1c :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h1d :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h1e :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h1f :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h20 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h21 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h22 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h23 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h24 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h25 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h26 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h27 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h28 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h29 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h2a :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h2b :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h2c :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h2d :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h2e :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h2f :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h30 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h31 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h32 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h33 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h34 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h35 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h36 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h37 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h38 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h39 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h3a :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h3b :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h3c :
		TR_72 = 9'h000 ;	// line#=../rle.cpp:68
	7'h3d :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h3e :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h3f :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h40 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h41 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h42 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h43 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h44 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h45 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h46 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h47 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h48 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h49 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h4a :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h4b :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h4c :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h4d :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h4e :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h4f :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h50 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h51 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h52 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h53 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h54 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h55 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h56 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h57 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h58 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h59 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h5a :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h5b :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h5c :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h5d :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h5e :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h5f :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h60 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h61 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h62 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h63 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h64 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h65 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h66 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h67 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h68 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h69 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h6a :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h6b :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h6c :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h6d :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h6e :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h6f :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h70 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h71 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h72 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h73 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h74 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h75 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h76 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h77 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h78 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h79 :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h7a :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h7b :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h7c :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h7d :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h7e :
		TR_72 = RG_quantized_block_rl_1 ;
	7'h7f :
		TR_72 = RG_quantized_block_rl_1 ;
	default :
		TR_72 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_2 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h01 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h02 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h03 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h04 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h05 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h06 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h07 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h08 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h09 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h0a :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h0b :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h0c :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h0d :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h0e :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h0f :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h10 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h11 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h12 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h13 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h14 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h15 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h16 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h17 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h18 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h19 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h1a :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h1b :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h1c :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h1d :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h1e :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h1f :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h20 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h21 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h22 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h23 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h24 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h25 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h26 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h27 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h28 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h29 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h2a :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h2b :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h2c :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h2d :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h2e :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h2f :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h30 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h31 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h32 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h33 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h34 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h35 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h36 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h37 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h38 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h39 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h3a :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h3b :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h3c :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h3d :
		TR_73 = 9'h000 ;	// line#=../rle.cpp:68
	7'h3e :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h3f :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h40 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h41 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h42 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h43 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h44 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h45 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h46 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h47 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h48 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h49 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h4a :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h4b :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h4c :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h4d :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h4e :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h4f :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h50 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h51 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h52 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h53 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h54 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h55 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h56 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h57 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h58 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h59 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h5a :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h5b :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h5c :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h5d :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h5e :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h5f :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h60 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h61 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h62 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h63 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h64 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h65 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h66 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h67 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h68 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h69 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h6a :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h6b :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h6c :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h6d :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h6e :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h6f :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h70 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h71 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h72 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h73 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h74 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h75 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h76 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h77 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h78 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h79 :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h7a :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h7b :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h7c :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h7d :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h7e :
		TR_73 = RG_quantized_block_rl_2 ;
	7'h7f :
		TR_73 = RG_quantized_block_rl_2 ;
	default :
		TR_73 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_3 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h01 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h02 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h03 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h04 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h05 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h06 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h07 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h08 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h09 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h0a :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h0b :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h0c :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h0d :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h0e :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h0f :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h10 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h11 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h12 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h13 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h14 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h15 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h16 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h17 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h18 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h19 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h1a :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h1b :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h1c :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h1d :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h1e :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h1f :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h20 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h21 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h22 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h23 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h24 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h25 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h26 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h27 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h28 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h29 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h2a :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h2b :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h2c :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h2d :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h2e :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h2f :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h30 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h31 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h32 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h33 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h34 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h35 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h36 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h37 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h38 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h39 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h3a :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h3b :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h3c :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h3d :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h3e :
		TR_74 = 9'h000 ;	// line#=../rle.cpp:68
	7'h3f :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h40 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h41 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h42 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h43 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h44 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h45 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h46 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h47 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h48 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h49 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h4a :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h4b :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h4c :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h4d :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h4e :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h4f :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h50 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h51 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h52 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h53 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h54 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h55 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h56 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h57 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h58 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h59 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h5a :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h5b :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h5c :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h5d :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h5e :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h5f :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h60 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h61 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h62 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h63 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h64 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h65 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h66 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h67 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h68 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h69 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h6a :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h6b :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h6c :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h6d :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h6e :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h6f :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h70 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h71 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h72 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h73 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h74 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h75 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h76 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h77 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h78 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h79 :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h7a :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h7b :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h7c :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h7d :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h7e :
		TR_74 = RG_quantized_block_rl_3 ;
	7'h7f :
		TR_74 = RG_quantized_block_rl_3 ;
	default :
		TR_74 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_4 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h01 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h02 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h03 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h04 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h05 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h06 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h07 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h08 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h09 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h0a :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h0b :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h0c :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h0d :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h0e :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h0f :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h10 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h11 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h12 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h13 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h14 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h15 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h16 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h17 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h18 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h19 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h1a :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h1b :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h1c :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h1d :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h1e :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h1f :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h20 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h21 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h22 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h23 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h24 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h25 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h26 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h27 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h28 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h29 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h2a :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h2b :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h2c :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h2d :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h2e :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h2f :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h30 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h31 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h32 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h33 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h34 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h35 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h36 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h37 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h38 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h39 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h3a :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h3b :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h3c :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h3d :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h3e :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h3f :
		TR_75 = 9'h000 ;	// line#=../rle.cpp:68
	7'h40 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h41 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h42 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h43 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h44 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h45 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h46 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h47 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h48 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h49 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h4a :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h4b :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h4c :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h4d :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h4e :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h4f :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h50 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h51 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h52 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h53 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h54 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h55 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h56 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h57 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h58 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h59 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h5a :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h5b :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h5c :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h5d :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h5e :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h5f :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h60 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h61 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h62 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h63 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h64 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h65 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h66 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h67 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h68 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h69 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h6a :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h6b :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h6c :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h6d :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h6e :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h6f :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h70 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h71 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h72 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h73 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h74 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h75 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h76 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h77 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h78 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h79 :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h7a :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h7b :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h7c :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h7d :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h7e :
		TR_75 = RG_quantized_block_rl_4 ;
	7'h7f :
		TR_75 = RG_quantized_block_rl_4 ;
	default :
		TR_75 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_5 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h01 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h02 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h03 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h04 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h05 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h06 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h07 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h08 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h09 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h0a :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h0b :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h0c :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h0d :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h0e :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h0f :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h10 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h11 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h12 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h13 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h14 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h15 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h16 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h17 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h18 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h19 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h1a :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h1b :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h1c :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h1d :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h1e :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h1f :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h20 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h21 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h22 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h23 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h24 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h25 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h26 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h27 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h28 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h29 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h2a :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h2b :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h2c :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h2d :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h2e :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h2f :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h30 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h31 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h32 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h33 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h34 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h35 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h36 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h37 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h38 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h39 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h3a :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h3b :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h3c :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h3d :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h3e :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h3f :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h40 :
		TR_76 = 9'h000 ;	// line#=../rle.cpp:68
	7'h41 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h42 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h43 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h44 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h45 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h46 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h47 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h48 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h49 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h4a :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h4b :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h4c :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h4d :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h4e :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h4f :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h50 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h51 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h52 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h53 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h54 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h55 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h56 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h57 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h58 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h59 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h5a :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h5b :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h5c :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h5d :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h5e :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h5f :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h60 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h61 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h62 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h63 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h64 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h65 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h66 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h67 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h68 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h69 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h6a :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h6b :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h6c :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h6d :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h6e :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h6f :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h70 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h71 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h72 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h73 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h74 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h75 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h76 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h77 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h78 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h79 :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h7a :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h7b :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h7c :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h7d :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h7e :
		TR_76 = RG_quantized_block_rl_5 ;
	7'h7f :
		TR_76 = RG_quantized_block_rl_5 ;
	default :
		TR_76 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_6 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h01 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h02 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h03 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h04 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h05 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h06 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h07 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h08 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h09 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h0a :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h0b :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h0c :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h0d :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h0e :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h0f :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h10 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h11 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h12 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h13 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h14 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h15 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h16 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h17 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h18 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h19 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h1a :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h1b :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h1c :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h1d :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h1e :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h1f :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h20 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h21 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h22 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h23 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h24 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h25 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h26 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h27 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h28 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h29 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h2a :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h2b :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h2c :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h2d :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h2e :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h2f :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h30 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h31 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h32 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h33 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h34 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h35 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h36 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h37 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h38 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h39 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h3a :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h3b :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h3c :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h3d :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h3e :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h3f :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h40 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h41 :
		TR_77 = 9'h000 ;	// line#=../rle.cpp:68
	7'h42 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h43 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h44 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h45 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h46 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h47 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h48 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h49 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h4a :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h4b :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h4c :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h4d :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h4e :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h4f :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h50 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h51 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h52 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h53 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h54 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h55 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h56 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h57 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h58 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h59 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h5a :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h5b :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h5c :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h5d :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h5e :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h5f :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h60 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h61 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h62 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h63 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h64 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h65 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h66 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h67 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h68 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h69 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h6a :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h6b :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h6c :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h6d :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h6e :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h6f :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h70 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h71 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h72 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h73 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h74 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h75 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h76 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h77 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h78 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h79 :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h7a :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h7b :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h7c :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h7d :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h7e :
		TR_77 = RG_quantized_block_rl_6 ;
	7'h7f :
		TR_77 = RG_quantized_block_rl_6 ;
	default :
		TR_77 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_7 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h01 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h02 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h03 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h04 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h05 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h06 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h07 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h08 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h09 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h0a :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h0b :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h0c :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h0d :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h0e :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h0f :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h10 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h11 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h12 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h13 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h14 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h15 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h16 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h17 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h18 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h19 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h1a :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h1b :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h1c :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h1d :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h1e :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h1f :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h20 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h21 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h22 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h23 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h24 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h25 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h26 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h27 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h28 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h29 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h2a :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h2b :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h2c :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h2d :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h2e :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h2f :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h30 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h31 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h32 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h33 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h34 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h35 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h36 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h37 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h38 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h39 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h3a :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h3b :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h3c :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h3d :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h3e :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h3f :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h40 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h41 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h42 :
		TR_78 = 9'h000 ;	// line#=../rle.cpp:68
	7'h43 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h44 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h45 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h46 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h47 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h48 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h49 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h4a :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h4b :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h4c :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h4d :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h4e :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h4f :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h50 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h51 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h52 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h53 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h54 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h55 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h56 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h57 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h58 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h59 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h5a :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h5b :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h5c :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h5d :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h5e :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h5f :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h60 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h61 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h62 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h63 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h64 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h65 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h66 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h67 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h68 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h69 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h6a :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h6b :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h6c :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h6d :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h6e :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h6f :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h70 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h71 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h72 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h73 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h74 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h75 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h76 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h77 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h78 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h79 :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h7a :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h7b :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h7c :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h7d :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h7e :
		TR_78 = RG_quantized_block_rl_7 ;
	7'h7f :
		TR_78 = RG_quantized_block_rl_7 ;
	default :
		TR_78 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_8 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h01 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h02 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h03 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h04 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h05 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h06 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h07 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h08 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h09 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h0a :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h0b :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h0c :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h0d :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h0e :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h0f :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h10 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h11 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h12 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h13 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h14 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h15 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h16 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h17 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h18 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h19 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h1a :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h1b :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h1c :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h1d :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h1e :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h1f :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h20 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h21 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h22 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h23 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h24 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h25 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h26 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h27 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h28 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h29 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h2a :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h2b :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h2c :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h2d :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h2e :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h2f :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h30 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h31 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h32 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h33 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h34 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h35 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h36 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h37 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h38 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h39 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h3a :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h3b :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h3c :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h3d :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h3e :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h3f :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h40 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h41 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h42 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h43 :
		TR_79 = 9'h000 ;	// line#=../rle.cpp:68
	7'h44 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h45 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h46 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h47 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h48 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h49 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h4a :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h4b :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h4c :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h4d :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h4e :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h4f :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h50 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h51 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h52 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h53 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h54 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h55 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h56 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h57 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h58 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h59 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h5a :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h5b :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h5c :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h5d :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h5e :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h5f :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h60 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h61 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h62 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h63 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h64 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h65 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h66 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h67 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h68 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h69 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h6a :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h6b :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h6c :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h6d :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h6e :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h6f :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h70 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h71 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h72 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h73 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h74 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h75 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h76 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h77 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h78 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h79 :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h7a :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h7b :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h7c :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h7d :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h7e :
		TR_79 = RG_quantized_block_rl_8 ;
	7'h7f :
		TR_79 = RG_quantized_block_rl_8 ;
	default :
		TR_79 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_9 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h01 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h02 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h03 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h04 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h05 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h06 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h07 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h08 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h09 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h0a :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h0b :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h0c :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h0d :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h0e :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h0f :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h10 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h11 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h12 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h13 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h14 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h15 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h16 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h17 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h18 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h19 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h1a :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h1b :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h1c :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h1d :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h1e :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h1f :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h20 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h21 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h22 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h23 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h24 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h25 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h26 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h27 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h28 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h29 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h2a :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h2b :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h2c :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h2d :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h2e :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h2f :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h30 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h31 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h32 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h33 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h34 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h35 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h36 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h37 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h38 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h39 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h3a :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h3b :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h3c :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h3d :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h3e :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h3f :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h40 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h41 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h42 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h43 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h44 :
		TR_80 = 9'h000 ;	// line#=../rle.cpp:68
	7'h45 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h46 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h47 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h48 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h49 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h4a :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h4b :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h4c :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h4d :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h4e :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h4f :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h50 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h51 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h52 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h53 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h54 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h55 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h56 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h57 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h58 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h59 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h5a :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h5b :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h5c :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h5d :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h5e :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h5f :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h60 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h61 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h62 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h63 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h64 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h65 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h66 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h67 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h68 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h69 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h6a :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h6b :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h6c :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h6d :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h6e :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h6f :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h70 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h71 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h72 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h73 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h74 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h75 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h76 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h77 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h78 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h79 :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h7a :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h7b :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h7c :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h7d :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h7e :
		TR_80 = RG_quantized_block_rl_9 ;
	7'h7f :
		TR_80 = RG_quantized_block_rl_9 ;
	default :
		TR_80 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_10 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h01 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h02 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h03 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h04 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h05 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h06 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h07 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h08 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h09 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h0a :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h0b :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h0c :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h0d :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h0e :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h0f :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h10 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h11 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h12 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h13 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h14 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h15 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h16 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h17 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h18 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h19 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h1a :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h1b :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h1c :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h1d :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h1e :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h1f :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h20 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h21 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h22 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h23 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h24 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h25 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h26 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h27 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h28 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h29 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h2a :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h2b :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h2c :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h2d :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h2e :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h2f :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h30 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h31 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h32 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h33 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h34 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h35 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h36 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h37 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h38 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h39 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h3a :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h3b :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h3c :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h3d :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h3e :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h3f :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h40 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h41 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h42 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h43 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h44 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h45 :
		TR_81 = 9'h000 ;	// line#=../rle.cpp:68
	7'h46 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h47 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h48 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h49 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h4a :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h4b :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h4c :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h4d :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h4e :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h4f :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h50 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h51 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h52 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h53 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h54 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h55 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h56 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h57 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h58 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h59 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h5a :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h5b :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h5c :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h5d :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h5e :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h5f :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h60 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h61 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h62 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h63 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h64 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h65 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h66 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h67 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h68 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h69 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h6a :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h6b :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h6c :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h6d :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h6e :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h6f :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h70 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h71 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h72 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h73 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h74 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h75 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h76 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h77 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h78 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h79 :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h7a :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h7b :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h7c :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h7d :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h7e :
		TR_81 = RG_quantized_block_rl_10 ;
	7'h7f :
		TR_81 = RG_quantized_block_rl_10 ;
	default :
		TR_81 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_11 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h01 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h02 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h03 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h04 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h05 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h06 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h07 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h08 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h09 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h0a :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h0b :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h0c :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h0d :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h0e :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h0f :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h10 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h11 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h12 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h13 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h14 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h15 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h16 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h17 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h18 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h19 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h1a :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h1b :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h1c :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h1d :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h1e :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h1f :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h20 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h21 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h22 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h23 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h24 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h25 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h26 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h27 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h28 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h29 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h2a :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h2b :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h2c :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h2d :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h2e :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h2f :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h30 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h31 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h32 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h33 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h34 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h35 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h36 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h37 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h38 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h39 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h3a :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h3b :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h3c :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h3d :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h3e :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h3f :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h40 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h41 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h42 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h43 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h44 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h45 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h46 :
		TR_82 = 9'h000 ;	// line#=../rle.cpp:68
	7'h47 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h48 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h49 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h4a :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h4b :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h4c :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h4d :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h4e :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h4f :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h50 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h51 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h52 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h53 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h54 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h55 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h56 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h57 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h58 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h59 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h5a :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h5b :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h5c :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h5d :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h5e :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h5f :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h60 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h61 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h62 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h63 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h64 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h65 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h66 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h67 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h68 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h69 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h6a :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h6b :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h6c :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h6d :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h6e :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h6f :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h70 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h71 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h72 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h73 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h74 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h75 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h76 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h77 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h78 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h79 :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h7a :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h7b :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h7c :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h7d :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h7e :
		TR_82 = RG_quantized_block_rl_11 ;
	7'h7f :
		TR_82 = RG_quantized_block_rl_11 ;
	default :
		TR_82 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_12 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h01 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h02 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h03 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h04 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h05 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h06 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h07 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h08 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h09 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h0a :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h0b :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h0c :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h0d :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h0e :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h0f :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h10 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h11 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h12 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h13 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h14 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h15 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h16 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h17 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h18 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h19 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h1a :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h1b :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h1c :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h1d :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h1e :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h1f :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h20 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h21 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h22 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h23 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h24 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h25 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h26 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h27 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h28 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h29 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h2a :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h2b :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h2c :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h2d :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h2e :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h2f :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h30 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h31 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h32 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h33 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h34 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h35 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h36 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h37 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h38 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h39 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h3a :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h3b :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h3c :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h3d :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h3e :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h3f :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h40 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h41 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h42 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h43 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h44 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h45 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h46 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h47 :
		TR_83 = 9'h000 ;	// line#=../rle.cpp:68
	7'h48 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h49 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h4a :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h4b :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h4c :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h4d :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h4e :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h4f :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h50 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h51 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h52 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h53 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h54 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h55 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h56 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h57 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h58 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h59 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h5a :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h5b :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h5c :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h5d :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h5e :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h5f :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h60 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h61 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h62 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h63 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h64 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h65 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h66 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h67 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h68 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h69 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h6a :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h6b :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h6c :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h6d :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h6e :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h6f :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h70 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h71 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h72 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h73 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h74 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h75 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h76 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h77 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h78 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h79 :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h7a :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h7b :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h7c :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h7d :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h7e :
		TR_83 = RG_quantized_block_rl_12 ;
	7'h7f :
		TR_83 = RG_quantized_block_rl_12 ;
	default :
		TR_83 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_13 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h01 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h02 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h03 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h04 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h05 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h06 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h07 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h08 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h09 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h0a :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h0b :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h0c :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h0d :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h0e :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h0f :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h10 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h11 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h12 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h13 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h14 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h15 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h16 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h17 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h18 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h19 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h1a :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h1b :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h1c :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h1d :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h1e :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h1f :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h20 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h21 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h22 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h23 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h24 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h25 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h26 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h27 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h28 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h29 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h2a :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h2b :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h2c :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h2d :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h2e :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h2f :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h30 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h31 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h32 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h33 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h34 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h35 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h36 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h37 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h38 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h39 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h3a :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h3b :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h3c :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h3d :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h3e :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h3f :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h40 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h41 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h42 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h43 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h44 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h45 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h46 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h47 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h48 :
		TR_84 = 9'h000 ;	// line#=../rle.cpp:68
	7'h49 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h4a :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h4b :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h4c :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h4d :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h4e :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h4f :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h50 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h51 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h52 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h53 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h54 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h55 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h56 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h57 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h58 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h59 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h5a :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h5b :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h5c :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h5d :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h5e :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h5f :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h60 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h61 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h62 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h63 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h64 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h65 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h66 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h67 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h68 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h69 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h6a :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h6b :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h6c :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h6d :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h6e :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h6f :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h70 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h71 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h72 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h73 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h74 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h75 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h76 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h77 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h78 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h79 :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h7a :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h7b :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h7c :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h7d :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h7e :
		TR_84 = RG_quantized_block_rl_13 ;
	7'h7f :
		TR_84 = RG_quantized_block_rl_13 ;
	default :
		TR_84 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_14 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h01 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h02 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h03 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h04 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h05 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h06 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h07 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h08 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h09 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h0a :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h0b :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h0c :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h0d :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h0e :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h0f :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h10 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h11 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h12 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h13 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h14 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h15 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h16 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h17 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h18 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h19 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h1a :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h1b :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h1c :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h1d :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h1e :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h1f :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h20 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h21 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h22 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h23 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h24 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h25 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h26 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h27 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h28 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h29 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h2a :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h2b :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h2c :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h2d :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h2e :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h2f :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h30 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h31 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h32 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h33 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h34 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h35 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h36 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h37 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h38 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h39 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h3a :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h3b :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h3c :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h3d :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h3e :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h3f :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h40 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h41 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h42 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h43 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h44 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h45 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h46 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h47 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h48 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h49 :
		TR_85 = 9'h000 ;	// line#=../rle.cpp:68
	7'h4a :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h4b :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h4c :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h4d :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h4e :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h4f :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h50 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h51 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h52 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h53 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h54 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h55 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h56 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h57 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h58 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h59 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h5a :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h5b :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h5c :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h5d :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h5e :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h5f :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h60 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h61 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h62 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h63 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h64 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h65 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h66 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h67 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h68 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h69 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h6a :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h6b :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h6c :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h6d :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h6e :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h6f :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h70 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h71 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h72 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h73 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h74 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h75 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h76 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h77 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h78 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h79 :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h7a :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h7b :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h7c :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h7d :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h7e :
		TR_85 = RG_quantized_block_rl_14 ;
	7'h7f :
		TR_85 = RG_quantized_block_rl_14 ;
	default :
		TR_85 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_15 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h01 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h02 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h03 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h04 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h05 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h06 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h07 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h08 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h09 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h0a :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h0b :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h0c :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h0d :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h0e :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h0f :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h10 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h11 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h12 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h13 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h14 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h15 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h16 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h17 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h18 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h19 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h1a :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h1b :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h1c :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h1d :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h1e :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h1f :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h20 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h21 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h22 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h23 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h24 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h25 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h26 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h27 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h28 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h29 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h2a :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h2b :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h2c :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h2d :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h2e :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h2f :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h30 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h31 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h32 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h33 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h34 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h35 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h36 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h37 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h38 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h39 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h3a :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h3b :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h3c :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h3d :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h3e :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h3f :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h40 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h41 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h42 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h43 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h44 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h45 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h46 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h47 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h48 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h49 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h4a :
		TR_86 = 9'h000 ;	// line#=../rle.cpp:68
	7'h4b :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h4c :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h4d :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h4e :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h4f :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h50 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h51 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h52 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h53 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h54 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h55 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h56 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h57 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h58 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h59 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h5a :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h5b :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h5c :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h5d :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h5e :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h5f :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h60 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h61 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h62 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h63 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h64 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h65 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h66 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h67 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h68 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h69 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h6a :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h6b :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h6c :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h6d :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h6e :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h6f :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h70 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h71 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h72 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h73 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h74 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h75 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h76 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h77 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h78 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h79 :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h7a :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h7b :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h7c :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h7d :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h7e :
		TR_86 = RG_quantized_block_rl_15 ;
	7'h7f :
		TR_86 = RG_quantized_block_rl_15 ;
	default :
		TR_86 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_16 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h01 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h02 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h03 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h04 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h05 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h06 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h07 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h08 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h09 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h0a :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h0b :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h0c :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h0d :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h0e :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h0f :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h10 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h11 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h12 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h13 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h14 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h15 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h16 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h17 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h18 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h19 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h1a :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h1b :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h1c :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h1d :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h1e :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h1f :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h20 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h21 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h22 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h23 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h24 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h25 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h26 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h27 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h28 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h29 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h2a :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h2b :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h2c :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h2d :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h2e :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h2f :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h30 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h31 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h32 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h33 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h34 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h35 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h36 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h37 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h38 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h39 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h3a :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h3b :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h3c :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h3d :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h3e :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h3f :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h40 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h41 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h42 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h43 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h44 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h45 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h46 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h47 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h48 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h49 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h4a :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h4b :
		TR_87 = 9'h000 ;	// line#=../rle.cpp:68
	7'h4c :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h4d :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h4e :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h4f :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h50 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h51 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h52 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h53 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h54 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h55 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h56 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h57 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h58 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h59 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h5a :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h5b :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h5c :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h5d :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h5e :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h5f :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h60 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h61 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h62 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h63 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h64 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h65 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h66 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h67 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h68 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h69 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h6a :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h6b :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h6c :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h6d :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h6e :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h6f :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h70 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h71 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h72 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h73 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h74 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h75 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h76 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h77 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h78 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h79 :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h7a :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h7b :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h7c :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h7d :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h7e :
		TR_87 = RG_quantized_block_rl_16 ;
	7'h7f :
		TR_87 = RG_quantized_block_rl_16 ;
	default :
		TR_87 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_17 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h01 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h02 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h03 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h04 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h05 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h06 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h07 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h08 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h09 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h0a :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h0b :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h0c :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h0d :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h0e :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h0f :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h10 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h11 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h12 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h13 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h14 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h15 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h16 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h17 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h18 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h19 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h1a :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h1b :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h1c :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h1d :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h1e :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h1f :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h20 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h21 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h22 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h23 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h24 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h25 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h26 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h27 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h28 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h29 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h2a :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h2b :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h2c :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h2d :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h2e :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h2f :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h30 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h31 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h32 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h33 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h34 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h35 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h36 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h37 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h38 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h39 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h3a :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h3b :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h3c :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h3d :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h3e :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h3f :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h40 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h41 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h42 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h43 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h44 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h45 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h46 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h47 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h48 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h49 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h4a :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h4b :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h4c :
		TR_88 = 9'h000 ;	// line#=../rle.cpp:68
	7'h4d :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h4e :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h4f :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h50 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h51 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h52 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h53 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h54 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h55 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h56 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h57 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h58 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h59 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h5a :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h5b :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h5c :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h5d :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h5e :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h5f :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h60 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h61 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h62 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h63 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h64 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h65 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h66 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h67 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h68 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h69 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h6a :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h6b :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h6c :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h6d :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h6e :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h6f :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h70 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h71 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h72 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h73 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h74 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h75 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h76 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h77 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h78 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h79 :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h7a :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h7b :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h7c :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h7d :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h7e :
		TR_88 = RG_quantized_block_rl_17 ;
	7'h7f :
		TR_88 = RG_quantized_block_rl_17 ;
	default :
		TR_88 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_18 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h01 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h02 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h03 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h04 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h05 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h06 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h07 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h08 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h09 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h0a :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h0b :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h0c :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h0d :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h0e :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h0f :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h10 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h11 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h12 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h13 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h14 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h15 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h16 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h17 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h18 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h19 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h1a :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h1b :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h1c :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h1d :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h1e :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h1f :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h20 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h21 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h22 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h23 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h24 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h25 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h26 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h27 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h28 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h29 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h2a :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h2b :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h2c :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h2d :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h2e :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h2f :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h30 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h31 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h32 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h33 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h34 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h35 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h36 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h37 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h38 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h39 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h3a :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h3b :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h3c :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h3d :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h3e :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h3f :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h40 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h41 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h42 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h43 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h44 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h45 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h46 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h47 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h48 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h49 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h4a :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h4b :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h4c :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h4d :
		TR_89 = 9'h000 ;	// line#=../rle.cpp:68
	7'h4e :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h4f :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h50 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h51 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h52 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h53 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h54 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h55 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h56 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h57 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h58 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h59 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h5a :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h5b :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h5c :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h5d :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h5e :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h5f :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h60 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h61 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h62 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h63 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h64 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h65 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h66 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h67 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h68 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h69 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h6a :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h6b :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h6c :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h6d :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h6e :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h6f :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h70 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h71 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h72 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h73 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h74 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h75 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h76 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h77 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h78 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h79 :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h7a :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h7b :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h7c :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h7d :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h7e :
		TR_89 = RG_quantized_block_rl_18 ;
	7'h7f :
		TR_89 = RG_quantized_block_rl_18 ;
	default :
		TR_89 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_19 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h01 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h02 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h03 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h04 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h05 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h06 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h07 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h08 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h09 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h0a :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h0b :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h0c :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h0d :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h0e :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h0f :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h10 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h11 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h12 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h13 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h14 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h15 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h16 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h17 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h18 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h19 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h1a :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h1b :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h1c :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h1d :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h1e :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h1f :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h20 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h21 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h22 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h23 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h24 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h25 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h26 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h27 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h28 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h29 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h2a :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h2b :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h2c :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h2d :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h2e :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h2f :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h30 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h31 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h32 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h33 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h34 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h35 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h36 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h37 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h38 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h39 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h3a :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h3b :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h3c :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h3d :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h3e :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h3f :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h40 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h41 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h42 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h43 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h44 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h45 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h46 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h47 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h48 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h49 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h4a :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h4b :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h4c :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h4d :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h4e :
		TR_90 = 9'h000 ;	// line#=../rle.cpp:68
	7'h4f :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h50 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h51 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h52 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h53 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h54 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h55 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h56 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h57 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h58 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h59 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h5a :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h5b :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h5c :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h5d :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h5e :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h5f :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h60 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h61 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h62 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h63 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h64 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h65 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h66 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h67 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h68 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h69 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h6a :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h6b :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h6c :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h6d :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h6e :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h6f :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h70 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h71 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h72 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h73 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h74 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h75 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h76 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h77 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h78 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h79 :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h7a :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h7b :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h7c :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h7d :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h7e :
		TR_90 = RG_quantized_block_rl_19 ;
	7'h7f :
		TR_90 = RG_quantized_block_rl_19 ;
	default :
		TR_90 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_20 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h01 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h02 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h03 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h04 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h05 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h06 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h07 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h08 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h09 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h0a :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h0b :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h0c :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h0d :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h0e :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h0f :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h10 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h11 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h12 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h13 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h14 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h15 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h16 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h17 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h18 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h19 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h1a :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h1b :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h1c :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h1d :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h1e :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h1f :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h20 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h21 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h22 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h23 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h24 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h25 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h26 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h27 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h28 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h29 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h2a :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h2b :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h2c :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h2d :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h2e :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h2f :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h30 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h31 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h32 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h33 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h34 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h35 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h36 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h37 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h38 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h39 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h3a :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h3b :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h3c :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h3d :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h3e :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h3f :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h40 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h41 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h42 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h43 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h44 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h45 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h46 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h47 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h48 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h49 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h4a :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h4b :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h4c :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h4d :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h4e :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h4f :
		TR_91 = 9'h000 ;	// line#=../rle.cpp:68
	7'h50 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h51 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h52 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h53 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h54 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h55 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h56 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h57 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h58 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h59 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h5a :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h5b :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h5c :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h5d :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h5e :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h5f :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h60 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h61 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h62 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h63 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h64 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h65 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h66 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h67 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h68 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h69 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h6a :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h6b :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h6c :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h6d :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h6e :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h6f :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h70 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h71 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h72 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h73 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h74 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h75 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h76 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h77 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h78 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h79 :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h7a :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h7b :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h7c :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h7d :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h7e :
		TR_91 = RG_quantized_block_rl_20 ;
	7'h7f :
		TR_91 = RG_quantized_block_rl_20 ;
	default :
		TR_91 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_21 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h01 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h02 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h03 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h04 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h05 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h06 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h07 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h08 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h09 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h0a :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h0b :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h0c :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h0d :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h0e :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h0f :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h10 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h11 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h12 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h13 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h14 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h15 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h16 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h17 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h18 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h19 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h1a :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h1b :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h1c :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h1d :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h1e :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h1f :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h20 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h21 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h22 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h23 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h24 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h25 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h26 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h27 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h28 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h29 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h2a :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h2b :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h2c :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h2d :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h2e :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h2f :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h30 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h31 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h32 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h33 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h34 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h35 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h36 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h37 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h38 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h39 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h3a :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h3b :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h3c :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h3d :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h3e :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h3f :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h40 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h41 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h42 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h43 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h44 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h45 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h46 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h47 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h48 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h49 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h4a :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h4b :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h4c :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h4d :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h4e :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h4f :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h50 :
		TR_92 = 9'h000 ;	// line#=../rle.cpp:68
	7'h51 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h52 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h53 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h54 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h55 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h56 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h57 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h58 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h59 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h5a :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h5b :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h5c :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h5d :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h5e :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h5f :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h60 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h61 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h62 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h63 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h64 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h65 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h66 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h67 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h68 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h69 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h6a :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h6b :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h6c :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h6d :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h6e :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h6f :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h70 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h71 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h72 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h73 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h74 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h75 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h76 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h77 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h78 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h79 :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h7a :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h7b :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h7c :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h7d :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h7e :
		TR_92 = RG_quantized_block_rl_21 ;
	7'h7f :
		TR_92 = RG_quantized_block_rl_21 ;
	default :
		TR_92 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_22 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h01 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h02 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h03 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h04 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h05 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h06 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h07 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h08 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h09 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h0a :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h0b :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h0c :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h0d :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h0e :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h0f :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h10 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h11 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h12 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h13 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h14 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h15 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h16 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h17 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h18 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h19 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h1a :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h1b :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h1c :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h1d :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h1e :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h1f :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h20 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h21 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h22 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h23 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h24 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h25 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h26 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h27 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h28 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h29 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h2a :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h2b :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h2c :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h2d :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h2e :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h2f :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h30 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h31 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h32 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h33 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h34 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h35 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h36 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h37 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h38 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h39 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h3a :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h3b :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h3c :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h3d :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h3e :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h3f :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h40 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h41 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h42 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h43 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h44 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h45 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h46 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h47 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h48 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h49 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h4a :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h4b :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h4c :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h4d :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h4e :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h4f :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h50 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h51 :
		TR_93 = 9'h000 ;	// line#=../rle.cpp:68
	7'h52 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h53 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h54 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h55 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h56 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h57 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h58 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h59 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h5a :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h5b :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h5c :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h5d :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h5e :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h5f :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h60 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h61 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h62 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h63 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h64 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h65 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h66 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h67 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h68 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h69 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h6a :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h6b :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h6c :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h6d :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h6e :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h6f :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h70 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h71 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h72 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h73 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h74 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h75 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h76 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h77 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h78 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h79 :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h7a :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h7b :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h7c :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h7d :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h7e :
		TR_93 = RG_quantized_block_rl_22 ;
	7'h7f :
		TR_93 = RG_quantized_block_rl_22 ;
	default :
		TR_93 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_23 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h01 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h02 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h03 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h04 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h05 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h06 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h07 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h08 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h09 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h0a :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h0b :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h0c :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h0d :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h0e :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h0f :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h10 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h11 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h12 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h13 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h14 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h15 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h16 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h17 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h18 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h19 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h1a :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h1b :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h1c :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h1d :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h1e :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h1f :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h20 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h21 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h22 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h23 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h24 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h25 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h26 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h27 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h28 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h29 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h2a :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h2b :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h2c :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h2d :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h2e :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h2f :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h30 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h31 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h32 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h33 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h34 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h35 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h36 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h37 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h38 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h39 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h3a :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h3b :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h3c :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h3d :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h3e :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h3f :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h40 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h41 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h42 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h43 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h44 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h45 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h46 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h47 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h48 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h49 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h4a :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h4b :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h4c :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h4d :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h4e :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h4f :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h50 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h51 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h52 :
		TR_94 = 9'h000 ;	// line#=../rle.cpp:68
	7'h53 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h54 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h55 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h56 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h57 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h58 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h59 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h5a :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h5b :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h5c :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h5d :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h5e :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h5f :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h60 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h61 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h62 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h63 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h64 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h65 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h66 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h67 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h68 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h69 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h6a :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h6b :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h6c :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h6d :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h6e :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h6f :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h70 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h71 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h72 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h73 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h74 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h75 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h76 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h77 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h78 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h79 :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h7a :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h7b :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h7c :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h7d :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h7e :
		TR_94 = RG_quantized_block_rl_23 ;
	7'h7f :
		TR_94 = RG_quantized_block_rl_23 ;
	default :
		TR_94 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_24 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h01 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h02 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h03 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h04 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h05 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h06 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h07 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h08 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h09 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h0a :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h0b :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h0c :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h0d :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h0e :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h0f :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h10 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h11 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h12 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h13 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h14 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h15 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h16 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h17 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h18 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h19 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h1a :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h1b :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h1c :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h1d :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h1e :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h1f :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h20 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h21 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h22 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h23 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h24 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h25 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h26 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h27 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h28 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h29 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h2a :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h2b :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h2c :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h2d :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h2e :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h2f :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h30 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h31 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h32 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h33 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h34 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h35 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h36 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h37 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h38 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h39 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h3a :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h3b :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h3c :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h3d :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h3e :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h3f :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h40 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h41 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h42 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h43 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h44 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h45 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h46 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h47 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h48 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h49 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h4a :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h4b :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h4c :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h4d :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h4e :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h4f :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h50 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h51 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h52 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h53 :
		TR_95 = 9'h000 ;	// line#=../rle.cpp:68
	7'h54 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h55 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h56 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h57 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h58 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h59 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h5a :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h5b :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h5c :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h5d :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h5e :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h5f :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h60 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h61 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h62 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h63 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h64 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h65 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h66 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h67 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h68 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h69 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h6a :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h6b :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h6c :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h6d :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h6e :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h6f :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h70 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h71 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h72 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h73 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h74 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h75 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h76 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h77 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h78 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h79 :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h7a :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h7b :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h7c :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h7d :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h7e :
		TR_95 = RG_quantized_block_rl_24 ;
	7'h7f :
		TR_95 = RG_quantized_block_rl_24 ;
	default :
		TR_95 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_25 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h01 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h02 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h03 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h04 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h05 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h06 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h07 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h08 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h09 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h0a :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h0b :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h0c :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h0d :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h0e :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h0f :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h10 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h11 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h12 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h13 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h14 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h15 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h16 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h17 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h18 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h19 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h1a :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h1b :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h1c :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h1d :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h1e :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h1f :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h20 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h21 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h22 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h23 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h24 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h25 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h26 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h27 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h28 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h29 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h2a :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h2b :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h2c :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h2d :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h2e :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h2f :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h30 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h31 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h32 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h33 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h34 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h35 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h36 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h37 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h38 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h39 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h3a :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h3b :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h3c :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h3d :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h3e :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h3f :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h40 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h41 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h42 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h43 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h44 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h45 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h46 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h47 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h48 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h49 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h4a :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h4b :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h4c :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h4d :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h4e :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h4f :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h50 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h51 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h52 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h53 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h54 :
		TR_96 = 9'h000 ;	// line#=../rle.cpp:68
	7'h55 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h56 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h57 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h58 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h59 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h5a :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h5b :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h5c :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h5d :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h5e :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h5f :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h60 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h61 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h62 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h63 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h64 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h65 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h66 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h67 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h68 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h69 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h6a :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h6b :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h6c :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h6d :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h6e :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h6f :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h70 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h71 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h72 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h73 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h74 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h75 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h76 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h77 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h78 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h79 :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h7a :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h7b :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h7c :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h7d :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h7e :
		TR_96 = RG_quantized_block_rl_25 ;
	7'h7f :
		TR_96 = RG_quantized_block_rl_25 ;
	default :
		TR_96 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_26 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h01 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h02 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h03 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h04 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h05 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h06 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h07 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h08 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h09 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h0a :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h0b :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h0c :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h0d :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h0e :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h0f :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h10 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h11 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h12 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h13 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h14 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h15 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h16 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h17 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h18 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h19 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h1a :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h1b :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h1c :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h1d :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h1e :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h1f :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h20 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h21 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h22 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h23 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h24 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h25 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h26 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h27 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h28 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h29 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h2a :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h2b :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h2c :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h2d :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h2e :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h2f :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h30 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h31 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h32 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h33 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h34 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h35 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h36 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h37 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h38 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h39 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h3a :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h3b :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h3c :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h3d :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h3e :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h3f :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h40 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h41 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h42 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h43 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h44 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h45 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h46 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h47 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h48 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h49 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h4a :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h4b :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h4c :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h4d :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h4e :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h4f :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h50 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h51 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h52 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h53 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h54 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h55 :
		TR_97 = 9'h000 ;	// line#=../rle.cpp:68
	7'h56 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h57 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h58 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h59 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h5a :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h5b :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h5c :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h5d :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h5e :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h5f :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h60 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h61 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h62 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h63 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h64 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h65 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h66 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h67 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h68 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h69 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h6a :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h6b :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h6c :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h6d :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h6e :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h6f :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h70 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h71 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h72 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h73 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h74 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h75 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h76 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h77 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h78 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h79 :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h7a :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h7b :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h7c :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h7d :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h7e :
		TR_97 = RG_quantized_block_rl_26 ;
	7'h7f :
		TR_97 = RG_quantized_block_rl_26 ;
	default :
		TR_97 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_27 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h01 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h02 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h03 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h04 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h05 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h06 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h07 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h08 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h09 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h0a :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h0b :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h0c :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h0d :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h0e :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h0f :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h10 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h11 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h12 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h13 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h14 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h15 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h16 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h17 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h18 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h19 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h1a :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h1b :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h1c :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h1d :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h1e :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h1f :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h20 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h21 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h22 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h23 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h24 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h25 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h26 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h27 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h28 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h29 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h2a :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h2b :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h2c :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h2d :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h2e :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h2f :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h30 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h31 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h32 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h33 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h34 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h35 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h36 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h37 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h38 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h39 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h3a :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h3b :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h3c :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h3d :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h3e :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h3f :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h40 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h41 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h42 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h43 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h44 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h45 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h46 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h47 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h48 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h49 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h4a :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h4b :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h4c :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h4d :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h4e :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h4f :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h50 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h51 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h52 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h53 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h54 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h55 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h56 :
		TR_98 = 9'h000 ;	// line#=../rle.cpp:68
	7'h57 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h58 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h59 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h5a :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h5b :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h5c :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h5d :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h5e :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h5f :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h60 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h61 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h62 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h63 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h64 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h65 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h66 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h67 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h68 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h69 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h6a :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h6b :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h6c :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h6d :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h6e :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h6f :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h70 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h71 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h72 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h73 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h74 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h75 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h76 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h77 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h78 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h79 :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h7a :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h7b :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h7c :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h7d :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h7e :
		TR_98 = RG_quantized_block_rl_27 ;
	7'h7f :
		TR_98 = RG_quantized_block_rl_27 ;
	default :
		TR_98 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_28 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h01 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h02 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h03 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h04 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h05 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h06 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h07 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h08 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h09 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h0a :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h0b :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h0c :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h0d :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h0e :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h0f :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h10 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h11 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h12 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h13 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h14 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h15 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h16 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h17 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h18 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h19 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h1a :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h1b :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h1c :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h1d :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h1e :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h1f :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h20 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h21 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h22 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h23 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h24 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h25 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h26 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h27 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h28 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h29 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h2a :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h2b :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h2c :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h2d :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h2e :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h2f :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h30 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h31 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h32 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h33 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h34 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h35 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h36 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h37 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h38 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h39 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h3a :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h3b :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h3c :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h3d :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h3e :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h3f :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h40 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h41 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h42 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h43 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h44 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h45 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h46 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h47 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h48 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h49 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h4a :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h4b :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h4c :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h4d :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h4e :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h4f :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h50 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h51 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h52 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h53 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h54 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h55 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h56 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h57 :
		TR_99 = 9'h000 ;	// line#=../rle.cpp:68
	7'h58 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h59 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h5a :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h5b :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h5c :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h5d :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h5e :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h5f :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h60 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h61 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h62 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h63 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h64 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h65 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h66 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h67 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h68 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h69 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h6a :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h6b :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h6c :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h6d :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h6e :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h6f :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h70 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h71 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h72 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h73 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h74 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h75 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h76 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h77 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h78 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h79 :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h7a :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h7b :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h7c :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h7d :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h7e :
		TR_99 = RG_quantized_block_rl_28 ;
	7'h7f :
		TR_99 = RG_quantized_block_rl_28 ;
	default :
		TR_99 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_29 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h01 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h02 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h03 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h04 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h05 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h06 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h07 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h08 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h09 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h0a :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h0b :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h0c :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h0d :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h0e :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h0f :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h10 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h11 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h12 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h13 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h14 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h15 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h16 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h17 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h18 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h19 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h1a :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h1b :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h1c :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h1d :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h1e :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h1f :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h20 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h21 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h22 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h23 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h24 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h25 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h26 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h27 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h28 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h29 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h2a :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h2b :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h2c :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h2d :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h2e :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h2f :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h30 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h31 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h32 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h33 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h34 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h35 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h36 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h37 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h38 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h39 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h3a :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h3b :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h3c :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h3d :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h3e :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h3f :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h40 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h41 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h42 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h43 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h44 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h45 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h46 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h47 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h48 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h49 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h4a :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h4b :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h4c :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h4d :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h4e :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h4f :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h50 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h51 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h52 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h53 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h54 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h55 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h56 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h57 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h58 :
		TR_100 = 9'h000 ;	// line#=../rle.cpp:68
	7'h59 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h5a :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h5b :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h5c :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h5d :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h5e :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h5f :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h60 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h61 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h62 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h63 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h64 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h65 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h66 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h67 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h68 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h69 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h6a :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h6b :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h6c :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h6d :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h6e :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h6f :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h70 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h71 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h72 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h73 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h74 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h75 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h76 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h77 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h78 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h79 :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h7a :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h7b :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h7c :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h7d :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h7e :
		TR_100 = RG_quantized_block_rl_29 ;
	7'h7f :
		TR_100 = RG_quantized_block_rl_29 ;
	default :
		TR_100 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_30 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h01 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h02 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h03 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h04 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h05 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h06 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h07 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h08 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h09 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h0a :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h0b :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h0c :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h0d :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h0e :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h0f :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h10 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h11 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h12 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h13 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h14 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h15 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h16 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h17 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h18 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h19 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h1a :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h1b :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h1c :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h1d :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h1e :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h1f :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h20 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h21 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h22 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h23 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h24 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h25 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h26 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h27 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h28 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h29 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h2a :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h2b :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h2c :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h2d :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h2e :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h2f :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h30 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h31 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h32 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h33 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h34 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h35 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h36 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h37 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h38 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h39 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h3a :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h3b :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h3c :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h3d :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h3e :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h3f :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h40 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h41 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h42 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h43 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h44 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h45 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h46 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h47 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h48 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h49 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h4a :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h4b :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h4c :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h4d :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h4e :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h4f :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h50 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h51 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h52 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h53 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h54 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h55 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h56 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h57 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h58 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h59 :
		TR_101 = 9'h000 ;	// line#=../rle.cpp:68
	7'h5a :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h5b :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h5c :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h5d :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h5e :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h5f :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h60 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h61 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h62 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h63 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h64 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h65 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h66 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h67 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h68 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h69 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h6a :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h6b :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h6c :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h6d :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h6e :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h6f :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h70 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h71 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h72 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h73 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h74 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h75 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h76 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h77 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h78 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h79 :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h7a :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h7b :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h7c :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h7d :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h7e :
		TR_101 = RG_quantized_block_rl_30 ;
	7'h7f :
		TR_101 = RG_quantized_block_rl_30 ;
	default :
		TR_101 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_31 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h01 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h02 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h03 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h04 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h05 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h06 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h07 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h08 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h09 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h0a :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h0b :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h0c :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h0d :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h0e :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h0f :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h10 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h11 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h12 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h13 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h14 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h15 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h16 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h17 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h18 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h19 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h1a :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h1b :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h1c :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h1d :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h1e :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h1f :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h20 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h21 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h22 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h23 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h24 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h25 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h26 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h27 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h28 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h29 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h2a :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h2b :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h2c :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h2d :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h2e :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h2f :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h30 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h31 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h32 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h33 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h34 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h35 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h36 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h37 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h38 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h39 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h3a :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h3b :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h3c :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h3d :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h3e :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h3f :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h40 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h41 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h42 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h43 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h44 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h45 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h46 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h47 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h48 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h49 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h4a :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h4b :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h4c :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h4d :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h4e :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h4f :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h50 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h51 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h52 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h53 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h54 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h55 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h56 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h57 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h58 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h59 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h5a :
		TR_102 = 9'h000 ;	// line#=../rle.cpp:68
	7'h5b :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h5c :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h5d :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h5e :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h5f :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h60 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h61 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h62 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h63 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h64 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h65 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h66 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h67 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h68 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h69 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h6a :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h6b :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h6c :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h6d :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h6e :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h6f :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h70 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h71 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h72 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h73 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h74 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h75 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h76 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h77 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h78 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h79 :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h7a :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h7b :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h7c :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h7d :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h7e :
		TR_102 = RG_quantized_block_rl_31 ;
	7'h7f :
		TR_102 = RG_quantized_block_rl_31 ;
	default :
		TR_102 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_32 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h01 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h02 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h03 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h04 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h05 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h06 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h07 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h08 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h09 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h0a :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h0b :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h0c :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h0d :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h0e :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h0f :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h10 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h11 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h12 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h13 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h14 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h15 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h16 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h17 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h18 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h19 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h1a :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h1b :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h1c :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h1d :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h1e :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h1f :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h20 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h21 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h22 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h23 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h24 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h25 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h26 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h27 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h28 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h29 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h2a :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h2b :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h2c :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h2d :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h2e :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h2f :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h30 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h31 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h32 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h33 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h34 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h35 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h36 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h37 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h38 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h39 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h3a :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h3b :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h3c :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h3d :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h3e :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h3f :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h40 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h41 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h42 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h43 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h44 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h45 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h46 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h47 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h48 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h49 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h4a :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h4b :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h4c :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h4d :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h4e :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h4f :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h50 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h51 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h52 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h53 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h54 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h55 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h56 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h57 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h58 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h59 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h5a :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h5b :
		TR_103 = 9'h000 ;	// line#=../rle.cpp:68
	7'h5c :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h5d :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h5e :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h5f :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h60 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h61 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h62 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h63 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h64 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h65 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h66 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h67 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h68 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h69 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h6a :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h6b :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h6c :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h6d :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h6e :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h6f :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h70 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h71 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h72 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h73 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h74 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h75 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h76 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h77 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h78 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h79 :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h7a :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h7b :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h7c :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h7d :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h7e :
		TR_103 = RG_quantized_block_rl_32 ;
	7'h7f :
		TR_103 = RG_quantized_block_rl_32 ;
	default :
		TR_103 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_33 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h01 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h02 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h03 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h04 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h05 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h06 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h07 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h08 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h09 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h0a :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h0b :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h0c :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h0d :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h0e :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h0f :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h10 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h11 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h12 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h13 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h14 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h15 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h16 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h17 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h18 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h19 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h1a :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h1b :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h1c :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h1d :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h1e :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h1f :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h20 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h21 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h22 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h23 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h24 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h25 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h26 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h27 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h28 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h29 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h2a :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h2b :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h2c :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h2d :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h2e :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h2f :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h30 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h31 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h32 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h33 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h34 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h35 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h36 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h37 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h38 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h39 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h3a :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h3b :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h3c :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h3d :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h3e :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h3f :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h40 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h41 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h42 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h43 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h44 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h45 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h46 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h47 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h48 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h49 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h4a :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h4b :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h4c :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h4d :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h4e :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h4f :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h50 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h51 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h52 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h53 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h54 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h55 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h56 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h57 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h58 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h59 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h5a :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h5b :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h5c :
		TR_104 = 9'h000 ;	// line#=../rle.cpp:68
	7'h5d :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h5e :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h5f :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h60 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h61 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h62 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h63 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h64 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h65 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h66 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h67 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h68 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h69 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h6a :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h6b :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h6c :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h6d :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h6e :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h6f :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h70 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h71 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h72 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h73 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h74 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h75 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h76 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h77 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h78 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h79 :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h7a :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h7b :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h7c :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h7d :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h7e :
		TR_104 = RG_quantized_block_rl_33 ;
	7'h7f :
		TR_104 = RG_quantized_block_rl_33 ;
	default :
		TR_104 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_34 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h01 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h02 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h03 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h04 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h05 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h06 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h07 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h08 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h09 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h0a :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h0b :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h0c :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h0d :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h0e :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h0f :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h10 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h11 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h12 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h13 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h14 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h15 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h16 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h17 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h18 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h19 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h1a :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h1b :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h1c :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h1d :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h1e :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h1f :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h20 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h21 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h22 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h23 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h24 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h25 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h26 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h27 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h28 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h29 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h2a :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h2b :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h2c :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h2d :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h2e :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h2f :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h30 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h31 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h32 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h33 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h34 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h35 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h36 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h37 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h38 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h39 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h3a :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h3b :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h3c :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h3d :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h3e :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h3f :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h40 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h41 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h42 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h43 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h44 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h45 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h46 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h47 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h48 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h49 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h4a :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h4b :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h4c :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h4d :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h4e :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h4f :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h50 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h51 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h52 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h53 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h54 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h55 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h56 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h57 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h58 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h59 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h5a :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h5b :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h5c :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h5d :
		TR_105 = 9'h000 ;	// line#=../rle.cpp:68
	7'h5e :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h5f :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h60 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h61 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h62 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h63 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h64 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h65 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h66 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h67 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h68 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h69 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h6a :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h6b :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h6c :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h6d :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h6e :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h6f :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h70 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h71 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h72 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h73 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h74 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h75 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h76 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h77 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h78 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h79 :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h7a :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h7b :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h7c :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h7d :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h7e :
		TR_105 = RG_quantized_block_rl_34 ;
	7'h7f :
		TR_105 = RG_quantized_block_rl_34 ;
	default :
		TR_105 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_35 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h01 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h02 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h03 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h04 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h05 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h06 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h07 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h08 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h09 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h0a :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h0b :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h0c :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h0d :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h0e :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h0f :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h10 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h11 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h12 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h13 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h14 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h15 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h16 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h17 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h18 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h19 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h1a :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h1b :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h1c :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h1d :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h1e :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h1f :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h20 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h21 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h22 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h23 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h24 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h25 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h26 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h27 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h28 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h29 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h2a :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h2b :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h2c :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h2d :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h2e :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h2f :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h30 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h31 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h32 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h33 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h34 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h35 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h36 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h37 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h38 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h39 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h3a :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h3b :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h3c :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h3d :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h3e :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h3f :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h40 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h41 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h42 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h43 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h44 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h45 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h46 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h47 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h48 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h49 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h4a :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h4b :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h4c :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h4d :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h4e :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h4f :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h50 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h51 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h52 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h53 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h54 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h55 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h56 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h57 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h58 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h59 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h5a :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h5b :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h5c :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h5d :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h5e :
		TR_106 = 9'h000 ;	// line#=../rle.cpp:68
	7'h5f :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h60 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h61 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h62 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h63 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h64 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h65 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h66 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h67 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h68 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h69 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h6a :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h6b :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h6c :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h6d :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h6e :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h6f :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h70 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h71 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h72 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h73 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h74 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h75 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h76 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h77 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h78 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h79 :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h7a :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h7b :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h7c :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h7d :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h7e :
		TR_106 = RG_quantized_block_rl_35 ;
	7'h7f :
		TR_106 = RG_quantized_block_rl_35 ;
	default :
		TR_106 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_36 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h01 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h02 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h03 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h04 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h05 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h06 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h07 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h08 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h09 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h0a :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h0b :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h0c :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h0d :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h0e :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h0f :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h10 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h11 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h12 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h13 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h14 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h15 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h16 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h17 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h18 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h19 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h1a :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h1b :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h1c :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h1d :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h1e :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h1f :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h20 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h21 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h22 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h23 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h24 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h25 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h26 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h27 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h28 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h29 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h2a :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h2b :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h2c :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h2d :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h2e :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h2f :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h30 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h31 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h32 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h33 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h34 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h35 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h36 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h37 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h38 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h39 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h3a :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h3b :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h3c :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h3d :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h3e :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h3f :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h40 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h41 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h42 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h43 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h44 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h45 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h46 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h47 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h48 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h49 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h4a :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h4b :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h4c :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h4d :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h4e :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h4f :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h50 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h51 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h52 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h53 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h54 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h55 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h56 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h57 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h58 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h59 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h5a :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h5b :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h5c :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h5d :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h5e :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h5f :
		TR_107 = 9'h000 ;	// line#=../rle.cpp:68
	7'h60 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h61 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h62 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h63 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h64 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h65 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h66 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h67 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h68 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h69 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h6a :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h6b :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h6c :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h6d :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h6e :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h6f :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h70 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h71 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h72 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h73 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h74 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h75 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h76 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h77 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h78 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h79 :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h7a :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h7b :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h7c :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h7d :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h7e :
		TR_107 = RG_quantized_block_rl_36 ;
	7'h7f :
		TR_107 = RG_quantized_block_rl_36 ;
	default :
		TR_107 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_37 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h01 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h02 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h03 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h04 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h05 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h06 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h07 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h08 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h09 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h0a :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h0b :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h0c :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h0d :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h0e :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h0f :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h10 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h11 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h12 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h13 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h14 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h15 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h16 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h17 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h18 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h19 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h1a :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h1b :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h1c :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h1d :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h1e :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h1f :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h20 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h21 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h22 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h23 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h24 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h25 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h26 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h27 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h28 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h29 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h2a :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h2b :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h2c :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h2d :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h2e :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h2f :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h30 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h31 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h32 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h33 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h34 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h35 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h36 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h37 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h38 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h39 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h3a :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h3b :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h3c :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h3d :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h3e :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h3f :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h40 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h41 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h42 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h43 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h44 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h45 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h46 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h47 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h48 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h49 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h4a :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h4b :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h4c :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h4d :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h4e :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h4f :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h50 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h51 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h52 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h53 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h54 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h55 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h56 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h57 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h58 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h59 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h5a :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h5b :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h5c :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h5d :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h5e :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h5f :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h60 :
		TR_108 = 9'h000 ;	// line#=../rle.cpp:68
	7'h61 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h62 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h63 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h64 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h65 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h66 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h67 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h68 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h69 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h6a :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h6b :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h6c :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h6d :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h6e :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h6f :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h70 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h71 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h72 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h73 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h74 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h75 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h76 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h77 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h78 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h79 :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h7a :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h7b :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h7c :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h7d :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h7e :
		TR_108 = RG_quantized_block_rl_37 ;
	7'h7f :
		TR_108 = RG_quantized_block_rl_37 ;
	default :
		TR_108 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_38 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h01 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h02 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h03 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h04 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h05 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h06 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h07 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h08 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h09 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h0a :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h0b :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h0c :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h0d :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h0e :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h0f :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h10 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h11 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h12 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h13 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h14 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h15 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h16 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h17 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h18 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h19 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h1a :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h1b :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h1c :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h1d :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h1e :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h1f :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h20 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h21 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h22 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h23 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h24 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h25 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h26 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h27 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h28 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h29 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h2a :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h2b :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h2c :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h2d :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h2e :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h2f :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h30 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h31 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h32 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h33 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h34 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h35 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h36 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h37 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h38 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h39 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h3a :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h3b :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h3c :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h3d :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h3e :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h3f :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h40 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h41 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h42 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h43 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h44 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h45 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h46 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h47 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h48 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h49 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h4a :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h4b :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h4c :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h4d :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h4e :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h4f :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h50 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h51 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h52 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h53 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h54 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h55 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h56 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h57 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h58 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h59 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h5a :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h5b :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h5c :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h5d :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h5e :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h5f :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h60 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h61 :
		TR_109 = 9'h000 ;	// line#=../rle.cpp:68
	7'h62 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h63 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h64 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h65 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h66 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h67 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h68 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h69 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h6a :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h6b :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h6c :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h6d :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h6e :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h6f :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h70 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h71 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h72 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h73 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h74 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h75 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h76 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h77 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h78 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h79 :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h7a :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h7b :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h7c :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h7d :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h7e :
		TR_109 = RG_quantized_block_rl_38 ;
	7'h7f :
		TR_109 = RG_quantized_block_rl_38 ;
	default :
		TR_109 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_39 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h01 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h02 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h03 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h04 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h05 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h06 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h07 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h08 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h09 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h0a :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h0b :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h0c :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h0d :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h0e :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h0f :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h10 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h11 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h12 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h13 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h14 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h15 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h16 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h17 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h18 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h19 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h1a :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h1b :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h1c :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h1d :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h1e :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h1f :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h20 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h21 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h22 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h23 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h24 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h25 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h26 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h27 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h28 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h29 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h2a :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h2b :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h2c :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h2d :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h2e :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h2f :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h30 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h31 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h32 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h33 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h34 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h35 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h36 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h37 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h38 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h39 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h3a :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h3b :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h3c :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h3d :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h3e :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h3f :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h40 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h41 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h42 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h43 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h44 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h45 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h46 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h47 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h48 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h49 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h4a :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h4b :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h4c :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h4d :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h4e :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h4f :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h50 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h51 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h52 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h53 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h54 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h55 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h56 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h57 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h58 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h59 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h5a :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h5b :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h5c :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h5d :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h5e :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h5f :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h60 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h61 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h62 :
		TR_110 = 9'h000 ;	// line#=../rle.cpp:68
	7'h63 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h64 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h65 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h66 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h67 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h68 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h69 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h6a :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h6b :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h6c :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h6d :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h6e :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h6f :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h70 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h71 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h72 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h73 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h74 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h75 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h76 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h77 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h78 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h79 :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h7a :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h7b :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h7c :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h7d :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h7e :
		TR_110 = RG_quantized_block_rl_39 ;
	7'h7f :
		TR_110 = RG_quantized_block_rl_39 ;
	default :
		TR_110 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_40 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h01 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h02 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h03 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h04 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h05 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h06 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h07 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h08 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h09 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h0a :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h0b :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h0c :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h0d :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h0e :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h0f :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h10 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h11 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h12 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h13 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h14 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h15 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h16 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h17 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h18 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h19 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h1a :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h1b :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h1c :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h1d :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h1e :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h1f :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h20 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h21 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h22 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h23 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h24 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h25 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h26 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h27 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h28 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h29 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h2a :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h2b :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h2c :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h2d :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h2e :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h2f :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h30 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h31 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h32 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h33 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h34 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h35 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h36 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h37 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h38 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h39 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h3a :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h3b :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h3c :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h3d :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h3e :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h3f :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h40 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h41 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h42 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h43 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h44 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h45 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h46 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h47 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h48 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h49 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h4a :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h4b :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h4c :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h4d :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h4e :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h4f :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h50 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h51 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h52 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h53 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h54 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h55 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h56 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h57 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h58 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h59 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h5a :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h5b :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h5c :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h5d :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h5e :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h5f :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h60 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h61 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h62 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h63 :
		TR_111 = 9'h000 ;	// line#=../rle.cpp:68
	7'h64 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h65 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h66 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h67 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h68 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h69 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h6a :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h6b :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h6c :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h6d :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h6e :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h6f :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h70 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h71 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h72 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h73 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h74 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h75 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h76 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h77 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h78 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h79 :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h7a :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h7b :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h7c :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h7d :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h7e :
		TR_111 = RG_quantized_block_rl_40 ;
	7'h7f :
		TR_111 = RG_quantized_block_rl_40 ;
	default :
		TR_111 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_41 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h01 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h02 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h03 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h04 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h05 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h06 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h07 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h08 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h09 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h0a :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h0b :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h0c :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h0d :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h0e :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h0f :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h10 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h11 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h12 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h13 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h14 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h15 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h16 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h17 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h18 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h19 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h1a :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h1b :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h1c :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h1d :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h1e :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h1f :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h20 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h21 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h22 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h23 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h24 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h25 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h26 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h27 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h28 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h29 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h2a :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h2b :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h2c :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h2d :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h2e :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h2f :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h30 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h31 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h32 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h33 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h34 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h35 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h36 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h37 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h38 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h39 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h3a :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h3b :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h3c :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h3d :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h3e :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h3f :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h40 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h41 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h42 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h43 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h44 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h45 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h46 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h47 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h48 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h49 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h4a :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h4b :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h4c :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h4d :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h4e :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h4f :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h50 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h51 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h52 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h53 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h54 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h55 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h56 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h57 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h58 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h59 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h5a :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h5b :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h5c :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h5d :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h5e :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h5f :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h60 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h61 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h62 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h63 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h64 :
		TR_112 = 9'h000 ;	// line#=../rle.cpp:68
	7'h65 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h66 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h67 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h68 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h69 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h6a :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h6b :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h6c :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h6d :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h6e :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h6f :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h70 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h71 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h72 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h73 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h74 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h75 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h76 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h77 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h78 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h79 :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h7a :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h7b :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h7c :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h7d :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h7e :
		TR_112 = RG_quantized_block_rl_41 ;
	7'h7f :
		TR_112 = RG_quantized_block_rl_41 ;
	default :
		TR_112 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_42 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h01 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h02 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h03 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h04 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h05 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h06 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h07 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h08 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h09 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h0a :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h0b :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h0c :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h0d :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h0e :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h0f :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h10 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h11 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h12 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h13 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h14 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h15 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h16 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h17 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h18 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h19 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h1a :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h1b :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h1c :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h1d :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h1e :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h1f :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h20 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h21 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h22 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h23 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h24 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h25 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h26 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h27 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h28 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h29 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h2a :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h2b :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h2c :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h2d :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h2e :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h2f :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h30 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h31 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h32 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h33 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h34 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h35 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h36 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h37 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h38 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h39 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h3a :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h3b :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h3c :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h3d :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h3e :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h3f :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h40 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h41 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h42 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h43 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h44 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h45 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h46 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h47 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h48 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h49 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h4a :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h4b :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h4c :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h4d :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h4e :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h4f :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h50 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h51 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h52 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h53 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h54 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h55 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h56 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h57 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h58 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h59 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h5a :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h5b :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h5c :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h5d :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h5e :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h5f :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h60 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h61 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h62 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h63 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h64 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h65 :
		TR_113 = 9'h000 ;	// line#=../rle.cpp:68
	7'h66 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h67 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h68 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h69 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h6a :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h6b :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h6c :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h6d :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h6e :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h6f :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h70 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h71 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h72 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h73 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h74 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h75 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h76 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h77 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h78 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h79 :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h7a :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h7b :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h7c :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h7d :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h7e :
		TR_113 = RG_quantized_block_rl_42 ;
	7'h7f :
		TR_113 = RG_quantized_block_rl_42 ;
	default :
		TR_113 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_43 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h01 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h02 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h03 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h04 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h05 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h06 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h07 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h08 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h09 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h0a :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h0b :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h0c :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h0d :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h0e :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h0f :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h10 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h11 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h12 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h13 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h14 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h15 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h16 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h17 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h18 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h19 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h1a :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h1b :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h1c :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h1d :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h1e :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h1f :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h20 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h21 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h22 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h23 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h24 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h25 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h26 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h27 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h28 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h29 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h2a :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h2b :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h2c :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h2d :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h2e :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h2f :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h30 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h31 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h32 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h33 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h34 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h35 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h36 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h37 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h38 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h39 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h3a :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h3b :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h3c :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h3d :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h3e :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h3f :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h40 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h41 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h42 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h43 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h44 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h45 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h46 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h47 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h48 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h49 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h4a :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h4b :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h4c :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h4d :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h4e :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h4f :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h50 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h51 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h52 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h53 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h54 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h55 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h56 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h57 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h58 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h59 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h5a :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h5b :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h5c :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h5d :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h5e :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h5f :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h60 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h61 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h62 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h63 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h64 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h65 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h66 :
		TR_114 = 9'h000 ;	// line#=../rle.cpp:68
	7'h67 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h68 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h69 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h6a :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h6b :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h6c :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h6d :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h6e :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h6f :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h70 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h71 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h72 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h73 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h74 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h75 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h76 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h77 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h78 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h79 :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h7a :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h7b :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h7c :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h7d :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h7e :
		TR_114 = RG_quantized_block_rl_43 ;
	7'h7f :
		TR_114 = RG_quantized_block_rl_43 ;
	default :
		TR_114 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_44 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h01 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h02 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h03 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h04 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h05 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h06 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h07 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h08 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h09 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h0a :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h0b :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h0c :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h0d :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h0e :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h0f :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h10 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h11 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h12 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h13 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h14 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h15 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h16 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h17 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h18 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h19 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h1a :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h1b :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h1c :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h1d :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h1e :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h1f :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h20 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h21 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h22 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h23 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h24 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h25 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h26 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h27 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h28 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h29 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h2a :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h2b :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h2c :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h2d :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h2e :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h2f :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h30 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h31 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h32 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h33 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h34 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h35 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h36 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h37 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h38 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h39 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h3a :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h3b :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h3c :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h3d :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h3e :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h3f :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h40 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h41 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h42 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h43 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h44 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h45 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h46 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h47 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h48 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h49 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h4a :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h4b :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h4c :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h4d :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h4e :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h4f :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h50 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h51 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h52 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h53 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h54 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h55 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h56 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h57 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h58 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h59 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h5a :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h5b :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h5c :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h5d :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h5e :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h5f :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h60 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h61 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h62 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h63 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h64 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h65 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h66 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h67 :
		TR_115 = 9'h000 ;	// line#=../rle.cpp:68
	7'h68 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h69 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h6a :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h6b :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h6c :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h6d :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h6e :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h6f :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h70 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h71 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h72 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h73 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h74 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h75 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h76 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h77 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h78 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h79 :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h7a :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h7b :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h7c :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h7d :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h7e :
		TR_115 = RG_quantized_block_rl_44 ;
	7'h7f :
		TR_115 = RG_quantized_block_rl_44 ;
	default :
		TR_115 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_45 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h01 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h02 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h03 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h04 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h05 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h06 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h07 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h08 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h09 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h0a :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h0b :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h0c :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h0d :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h0e :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h0f :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h10 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h11 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h12 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h13 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h14 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h15 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h16 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h17 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h18 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h19 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h1a :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h1b :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h1c :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h1d :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h1e :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h1f :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h20 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h21 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h22 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h23 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h24 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h25 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h26 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h27 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h28 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h29 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h2a :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h2b :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h2c :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h2d :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h2e :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h2f :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h30 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h31 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h32 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h33 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h34 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h35 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h36 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h37 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h38 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h39 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h3a :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h3b :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h3c :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h3d :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h3e :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h3f :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h40 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h41 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h42 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h43 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h44 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h45 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h46 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h47 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h48 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h49 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h4a :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h4b :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h4c :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h4d :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h4e :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h4f :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h50 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h51 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h52 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h53 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h54 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h55 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h56 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h57 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h58 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h59 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h5a :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h5b :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h5c :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h5d :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h5e :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h5f :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h60 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h61 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h62 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h63 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h64 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h65 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h66 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h67 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h68 :
		TR_116 = 9'h000 ;	// line#=../rle.cpp:68
	7'h69 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h6a :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h6b :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h6c :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h6d :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h6e :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h6f :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h70 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h71 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h72 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h73 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h74 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h75 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h76 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h77 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h78 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h79 :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h7a :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h7b :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h7c :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h7d :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h7e :
		TR_116 = RG_quantized_block_rl_45 ;
	7'h7f :
		TR_116 = RG_quantized_block_rl_45 ;
	default :
		TR_116 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_46 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h01 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h02 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h03 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h04 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h05 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h06 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h07 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h08 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h09 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h0a :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h0b :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h0c :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h0d :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h0e :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h0f :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h10 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h11 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h12 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h13 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h14 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h15 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h16 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h17 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h18 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h19 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h1a :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h1b :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h1c :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h1d :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h1e :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h1f :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h20 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h21 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h22 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h23 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h24 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h25 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h26 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h27 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h28 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h29 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h2a :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h2b :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h2c :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h2d :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h2e :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h2f :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h30 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h31 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h32 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h33 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h34 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h35 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h36 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h37 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h38 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h39 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h3a :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h3b :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h3c :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h3d :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h3e :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h3f :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h40 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h41 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h42 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h43 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h44 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h45 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h46 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h47 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h48 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h49 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h4a :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h4b :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h4c :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h4d :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h4e :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h4f :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h50 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h51 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h52 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h53 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h54 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h55 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h56 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h57 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h58 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h59 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h5a :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h5b :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h5c :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h5d :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h5e :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h5f :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h60 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h61 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h62 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h63 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h64 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h65 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h66 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h67 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h68 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h69 :
		TR_117 = 9'h000 ;	// line#=../rle.cpp:68
	7'h6a :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h6b :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h6c :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h6d :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h6e :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h6f :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h70 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h71 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h72 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h73 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h74 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h75 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h76 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h77 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h78 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h79 :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h7a :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h7b :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h7c :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h7d :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h7e :
		TR_117 = RG_quantized_block_rl_46 ;
	7'h7f :
		TR_117 = RG_quantized_block_rl_46 ;
	default :
		TR_117 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_47 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h01 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h02 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h03 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h04 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h05 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h06 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h07 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h08 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h09 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h0a :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h0b :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h0c :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h0d :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h0e :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h0f :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h10 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h11 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h12 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h13 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h14 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h15 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h16 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h17 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h18 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h19 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h1a :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h1b :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h1c :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h1d :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h1e :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h1f :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h20 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h21 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h22 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h23 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h24 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h25 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h26 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h27 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h28 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h29 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h2a :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h2b :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h2c :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h2d :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h2e :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h2f :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h30 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h31 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h32 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h33 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h34 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h35 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h36 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h37 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h38 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h39 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h3a :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h3b :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h3c :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h3d :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h3e :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h3f :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h40 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h41 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h42 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h43 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h44 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h45 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h46 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h47 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h48 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h49 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h4a :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h4b :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h4c :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h4d :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h4e :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h4f :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h50 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h51 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h52 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h53 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h54 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h55 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h56 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h57 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h58 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h59 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h5a :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h5b :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h5c :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h5d :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h5e :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h5f :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h60 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h61 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h62 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h63 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h64 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h65 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h66 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h67 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h68 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h69 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h6a :
		TR_118 = 9'h000 ;	// line#=../rle.cpp:68
	7'h6b :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h6c :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h6d :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h6e :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h6f :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h70 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h71 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h72 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h73 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h74 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h75 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h76 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h77 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h78 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h79 :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h7a :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h7b :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h7c :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h7d :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h7e :
		TR_118 = RG_quantized_block_rl_47 ;
	7'h7f :
		TR_118 = RG_quantized_block_rl_47 ;
	default :
		TR_118 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_48 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h01 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h02 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h03 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h04 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h05 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h06 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h07 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h08 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h09 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h0a :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h0b :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h0c :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h0d :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h0e :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h0f :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h10 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h11 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h12 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h13 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h14 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h15 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h16 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h17 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h18 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h19 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h1a :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h1b :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h1c :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h1d :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h1e :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h1f :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h20 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h21 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h22 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h23 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h24 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h25 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h26 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h27 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h28 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h29 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h2a :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h2b :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h2c :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h2d :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h2e :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h2f :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h30 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h31 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h32 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h33 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h34 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h35 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h36 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h37 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h38 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h39 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h3a :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h3b :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h3c :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h3d :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h3e :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h3f :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h40 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h41 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h42 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h43 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h44 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h45 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h46 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h47 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h48 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h49 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h4a :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h4b :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h4c :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h4d :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h4e :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h4f :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h50 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h51 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h52 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h53 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h54 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h55 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h56 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h57 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h58 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h59 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h5a :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h5b :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h5c :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h5d :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h5e :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h5f :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h60 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h61 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h62 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h63 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h64 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h65 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h66 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h67 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h68 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h69 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h6a :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h6b :
		TR_119 = 9'h000 ;	// line#=../rle.cpp:68
	7'h6c :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h6d :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h6e :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h6f :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h70 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h71 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h72 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h73 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h74 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h75 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h76 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h77 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h78 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h79 :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h7a :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h7b :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h7c :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h7d :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h7e :
		TR_119 = RG_quantized_block_rl_48 ;
	7'h7f :
		TR_119 = RG_quantized_block_rl_48 ;
	default :
		TR_119 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_49 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h01 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h02 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h03 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h04 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h05 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h06 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h07 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h08 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h09 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h0a :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h0b :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h0c :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h0d :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h0e :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h0f :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h10 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h11 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h12 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h13 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h14 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h15 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h16 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h17 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h18 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h19 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h1a :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h1b :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h1c :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h1d :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h1e :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h1f :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h20 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h21 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h22 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h23 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h24 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h25 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h26 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h27 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h28 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h29 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h2a :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h2b :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h2c :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h2d :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h2e :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h2f :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h30 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h31 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h32 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h33 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h34 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h35 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h36 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h37 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h38 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h39 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h3a :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h3b :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h3c :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h3d :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h3e :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h3f :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h40 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h41 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h42 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h43 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h44 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h45 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h46 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h47 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h48 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h49 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h4a :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h4b :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h4c :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h4d :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h4e :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h4f :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h50 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h51 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h52 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h53 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h54 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h55 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h56 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h57 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h58 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h59 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h5a :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h5b :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h5c :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h5d :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h5e :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h5f :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h60 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h61 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h62 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h63 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h64 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h65 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h66 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h67 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h68 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h69 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h6a :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h6b :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h6c :
		TR_120 = 9'h000 ;	// line#=../rle.cpp:68
	7'h6d :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h6e :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h6f :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h70 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h71 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h72 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h73 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h74 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h75 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h76 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h77 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h78 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h79 :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h7a :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h7b :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h7c :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h7d :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h7e :
		TR_120 = RG_quantized_block_rl_49 ;
	7'h7f :
		TR_120 = RG_quantized_block_rl_49 ;
	default :
		TR_120 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_50 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h01 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h02 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h03 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h04 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h05 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h06 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h07 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h08 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h09 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h0a :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h0b :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h0c :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h0d :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h0e :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h0f :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h10 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h11 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h12 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h13 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h14 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h15 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h16 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h17 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h18 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h19 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h1a :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h1b :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h1c :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h1d :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h1e :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h1f :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h20 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h21 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h22 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h23 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h24 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h25 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h26 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h27 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h28 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h29 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h2a :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h2b :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h2c :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h2d :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h2e :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h2f :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h30 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h31 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h32 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h33 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h34 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h35 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h36 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h37 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h38 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h39 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h3a :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h3b :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h3c :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h3d :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h3e :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h3f :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h40 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h41 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h42 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h43 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h44 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h45 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h46 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h47 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h48 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h49 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h4a :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h4b :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h4c :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h4d :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h4e :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h4f :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h50 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h51 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h52 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h53 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h54 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h55 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h56 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h57 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h58 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h59 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h5a :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h5b :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h5c :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h5d :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h5e :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h5f :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h60 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h61 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h62 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h63 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h64 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h65 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h66 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h67 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h68 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h69 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h6a :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h6b :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h6c :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h6d :
		TR_121 = 9'h000 ;	// line#=../rle.cpp:68
	7'h6e :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h6f :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h70 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h71 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h72 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h73 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h74 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h75 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h76 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h77 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h78 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h79 :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h7a :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h7b :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h7c :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h7d :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h7e :
		TR_121 = RG_quantized_block_rl_50 ;
	7'h7f :
		TR_121 = RG_quantized_block_rl_50 ;
	default :
		TR_121 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_51 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h01 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h02 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h03 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h04 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h05 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h06 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h07 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h08 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h09 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h0a :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h0b :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h0c :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h0d :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h0e :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h0f :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h10 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h11 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h12 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h13 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h14 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h15 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h16 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h17 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h18 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h19 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h1a :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h1b :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h1c :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h1d :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h1e :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h1f :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h20 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h21 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h22 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h23 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h24 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h25 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h26 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h27 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h28 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h29 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h2a :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h2b :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h2c :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h2d :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h2e :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h2f :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h30 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h31 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h32 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h33 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h34 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h35 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h36 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h37 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h38 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h39 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h3a :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h3b :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h3c :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h3d :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h3e :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h3f :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h40 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h41 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h42 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h43 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h44 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h45 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h46 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h47 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h48 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h49 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h4a :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h4b :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h4c :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h4d :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h4e :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h4f :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h50 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h51 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h52 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h53 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h54 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h55 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h56 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h57 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h58 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h59 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h5a :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h5b :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h5c :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h5d :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h5e :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h5f :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h60 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h61 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h62 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h63 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h64 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h65 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h66 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h67 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h68 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h69 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h6a :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h6b :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h6c :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h6d :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h6e :
		TR_122 = 9'h000 ;	// line#=../rle.cpp:68
	7'h6f :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h70 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h71 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h72 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h73 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h74 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h75 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h76 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h77 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h78 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h79 :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h7a :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h7b :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h7c :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h7d :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h7e :
		TR_122 = RG_quantized_block_rl_51 ;
	7'h7f :
		TR_122 = RG_quantized_block_rl_51 ;
	default :
		TR_122 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_52 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h01 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h02 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h03 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h04 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h05 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h06 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h07 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h08 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h09 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h0a :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h0b :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h0c :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h0d :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h0e :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h0f :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h10 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h11 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h12 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h13 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h14 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h15 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h16 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h17 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h18 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h19 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h1a :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h1b :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h1c :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h1d :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h1e :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h1f :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h20 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h21 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h22 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h23 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h24 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h25 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h26 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h27 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h28 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h29 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h2a :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h2b :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h2c :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h2d :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h2e :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h2f :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h30 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h31 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h32 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h33 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h34 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h35 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h36 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h37 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h38 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h39 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h3a :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h3b :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h3c :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h3d :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h3e :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h3f :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h40 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h41 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h42 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h43 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h44 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h45 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h46 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h47 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h48 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h49 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h4a :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h4b :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h4c :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h4d :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h4e :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h4f :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h50 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h51 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h52 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h53 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h54 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h55 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h56 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h57 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h58 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h59 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h5a :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h5b :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h5c :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h5d :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h5e :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h5f :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h60 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h61 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h62 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h63 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h64 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h65 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h66 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h67 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h68 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h69 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h6a :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h6b :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h6c :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h6d :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h6e :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h6f :
		TR_123 = 9'h000 ;	// line#=../rle.cpp:68
	7'h70 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h71 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h72 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h73 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h74 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h75 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h76 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h77 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h78 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h79 :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h7a :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h7b :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h7c :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h7d :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h7e :
		TR_123 = RG_quantized_block_rl_52 ;
	7'h7f :
		TR_123 = RG_quantized_block_rl_52 ;
	default :
		TR_123 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_53 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h01 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h02 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h03 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h04 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h05 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h06 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h07 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h08 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h09 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h0a :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h0b :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h0c :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h0d :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h0e :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h0f :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h10 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h11 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h12 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h13 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h14 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h15 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h16 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h17 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h18 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h19 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h1a :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h1b :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h1c :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h1d :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h1e :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h1f :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h20 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h21 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h22 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h23 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h24 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h25 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h26 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h27 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h28 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h29 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h2a :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h2b :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h2c :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h2d :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h2e :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h2f :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h30 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h31 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h32 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h33 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h34 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h35 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h36 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h37 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h38 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h39 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h3a :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h3b :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h3c :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h3d :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h3e :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h3f :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h40 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h41 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h42 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h43 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h44 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h45 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h46 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h47 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h48 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h49 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h4a :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h4b :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h4c :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h4d :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h4e :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h4f :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h50 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h51 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h52 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h53 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h54 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h55 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h56 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h57 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h58 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h59 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h5a :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h5b :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h5c :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h5d :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h5e :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h5f :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h60 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h61 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h62 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h63 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h64 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h65 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h66 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h67 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h68 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h69 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h6a :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h6b :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h6c :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h6d :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h6e :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h6f :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h70 :
		TR_124 = 9'h000 ;	// line#=../rle.cpp:68
	7'h71 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h72 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h73 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h74 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h75 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h76 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h77 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h78 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h79 :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h7a :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h7b :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h7c :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h7d :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h7e :
		TR_124 = RG_quantized_block_rl_53 ;
	7'h7f :
		TR_124 = RG_quantized_block_rl_53 ;
	default :
		TR_124 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_54 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h01 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h02 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h03 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h04 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h05 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h06 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h07 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h08 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h09 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h0f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h10 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h11 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h12 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h13 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h14 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h15 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h16 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h17 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h18 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h19 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h1f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h20 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h21 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h22 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h23 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h24 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h25 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h26 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h27 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h28 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h29 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h2f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h30 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h31 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h32 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h33 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h34 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h35 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h36 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h37 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h38 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h39 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h3f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h40 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h41 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h42 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h43 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h44 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h45 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h46 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h47 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h48 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h49 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h4f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h50 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h51 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h52 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h53 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h54 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h55 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h56 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h57 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h58 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h59 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h5f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h60 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h61 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h62 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h63 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h64 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h65 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h66 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h67 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h68 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h69 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h6f :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h70 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h71 :
		TR_125 = 9'h000 ;	// line#=../rle.cpp:68
	7'h72 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h73 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h74 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h75 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h76 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h77 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h78 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h79 :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7a :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7b :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7c :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7d :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7e :
		TR_125 = RG_quantized_block_rl_54 ;
	7'h7f :
		TR_125 = RG_quantized_block_rl_54 ;
	default :
		TR_125 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_55 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h01 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h02 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h03 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h04 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h05 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h06 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h07 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h08 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h09 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h0a :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h0b :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h0c :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h0d :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h0e :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h0f :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h10 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h11 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h12 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h13 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h14 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h15 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h16 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h17 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h18 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h19 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h1a :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h1b :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h1c :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h1d :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h1e :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h1f :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h20 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h21 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h22 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h23 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h24 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h25 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h26 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h27 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h28 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h29 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h2a :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h2b :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h2c :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h2d :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h2e :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h2f :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h30 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h31 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h32 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h33 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h34 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h35 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h36 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h37 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h38 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h39 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h3a :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h3b :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h3c :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h3d :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h3e :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h3f :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h40 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h41 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h42 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h43 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h44 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h45 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h46 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h47 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h48 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h49 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h4a :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h4b :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h4c :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h4d :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h4e :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h4f :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h50 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h51 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h52 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h53 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h54 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h55 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h56 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h57 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h58 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h59 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h5a :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h5b :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h5c :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h5d :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h5e :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h5f :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h60 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h61 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h62 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h63 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h64 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h65 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h66 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h67 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h68 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h69 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h6a :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h6b :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h6c :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h6d :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h6e :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h6f :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h70 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h71 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h72 :
		TR_126 = 9'h000 ;	// line#=../rle.cpp:68
	7'h73 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h74 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h75 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h76 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h77 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h78 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h79 :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h7a :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h7b :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h7c :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h7d :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h7e :
		TR_126 = RG_quantized_block_rl_55 ;
	7'h7f :
		TR_126 = RG_quantized_block_rl_55 ;
	default :
		TR_126 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_56 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h01 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h02 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h03 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h04 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h05 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h06 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h07 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h08 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h09 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h0a :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h0b :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h0c :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h0d :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h0e :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h0f :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h10 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h11 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h12 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h13 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h14 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h15 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h16 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h17 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h18 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h19 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h1a :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h1b :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h1c :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h1d :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h1e :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h1f :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h20 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h21 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h22 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h23 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h24 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h25 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h26 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h27 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h28 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h29 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h2a :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h2b :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h2c :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h2d :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h2e :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h2f :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h30 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h31 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h32 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h33 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h34 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h35 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h36 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h37 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h38 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h39 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h3a :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h3b :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h3c :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h3d :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h3e :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h3f :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h40 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h41 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h42 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h43 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h44 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h45 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h46 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h47 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h48 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h49 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h4a :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h4b :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h4c :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h4d :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h4e :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h4f :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h50 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h51 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h52 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h53 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h54 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h55 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h56 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h57 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h58 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h59 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h5a :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h5b :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h5c :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h5d :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h5e :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h5f :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h60 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h61 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h62 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h63 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h64 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h65 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h66 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h67 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h68 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h69 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h6a :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h6b :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h6c :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h6d :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h6e :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h6f :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h70 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h71 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h72 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h73 :
		TR_127 = 9'h000 ;	// line#=../rle.cpp:68
	7'h74 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h75 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h76 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h77 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h78 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h79 :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h7a :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h7b :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h7c :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h7d :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h7e :
		TR_127 = RG_quantized_block_rl_56 ;
	7'h7f :
		TR_127 = RG_quantized_block_rl_56 ;
	default :
		TR_127 = 9'hx ;
	endcase
always @ ( RG_rl_242 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_128 = RG_rl_242 ;
	7'h01 :
		TR_128 = RG_rl_242 ;
	7'h02 :
		TR_128 = RG_rl_242 ;
	7'h03 :
		TR_128 = RG_rl_242 ;
	7'h04 :
		TR_128 = RG_rl_242 ;
	7'h05 :
		TR_128 = RG_rl_242 ;
	7'h06 :
		TR_128 = RG_rl_242 ;
	7'h07 :
		TR_128 = RG_rl_242 ;
	7'h08 :
		TR_128 = RG_rl_242 ;
	7'h09 :
		TR_128 = RG_rl_242 ;
	7'h0a :
		TR_128 = RG_rl_242 ;
	7'h0b :
		TR_128 = RG_rl_242 ;
	7'h0c :
		TR_128 = RG_rl_242 ;
	7'h0d :
		TR_128 = RG_rl_242 ;
	7'h0e :
		TR_128 = RG_rl_242 ;
	7'h0f :
		TR_128 = RG_rl_242 ;
	7'h10 :
		TR_128 = RG_rl_242 ;
	7'h11 :
		TR_128 = RG_rl_242 ;
	7'h12 :
		TR_128 = RG_rl_242 ;
	7'h13 :
		TR_128 = RG_rl_242 ;
	7'h14 :
		TR_128 = RG_rl_242 ;
	7'h15 :
		TR_128 = RG_rl_242 ;
	7'h16 :
		TR_128 = RG_rl_242 ;
	7'h17 :
		TR_128 = RG_rl_242 ;
	7'h18 :
		TR_128 = RG_rl_242 ;
	7'h19 :
		TR_128 = RG_rl_242 ;
	7'h1a :
		TR_128 = RG_rl_242 ;
	7'h1b :
		TR_128 = RG_rl_242 ;
	7'h1c :
		TR_128 = RG_rl_242 ;
	7'h1d :
		TR_128 = RG_rl_242 ;
	7'h1e :
		TR_128 = RG_rl_242 ;
	7'h1f :
		TR_128 = RG_rl_242 ;
	7'h20 :
		TR_128 = RG_rl_242 ;
	7'h21 :
		TR_128 = RG_rl_242 ;
	7'h22 :
		TR_128 = RG_rl_242 ;
	7'h23 :
		TR_128 = RG_rl_242 ;
	7'h24 :
		TR_128 = RG_rl_242 ;
	7'h25 :
		TR_128 = RG_rl_242 ;
	7'h26 :
		TR_128 = RG_rl_242 ;
	7'h27 :
		TR_128 = RG_rl_242 ;
	7'h28 :
		TR_128 = RG_rl_242 ;
	7'h29 :
		TR_128 = RG_rl_242 ;
	7'h2a :
		TR_128 = RG_rl_242 ;
	7'h2b :
		TR_128 = RG_rl_242 ;
	7'h2c :
		TR_128 = RG_rl_242 ;
	7'h2d :
		TR_128 = RG_rl_242 ;
	7'h2e :
		TR_128 = RG_rl_242 ;
	7'h2f :
		TR_128 = RG_rl_242 ;
	7'h30 :
		TR_128 = RG_rl_242 ;
	7'h31 :
		TR_128 = RG_rl_242 ;
	7'h32 :
		TR_128 = RG_rl_242 ;
	7'h33 :
		TR_128 = RG_rl_242 ;
	7'h34 :
		TR_128 = RG_rl_242 ;
	7'h35 :
		TR_128 = RG_rl_242 ;
	7'h36 :
		TR_128 = RG_rl_242 ;
	7'h37 :
		TR_128 = RG_rl_242 ;
	7'h38 :
		TR_128 = RG_rl_242 ;
	7'h39 :
		TR_128 = RG_rl_242 ;
	7'h3a :
		TR_128 = RG_rl_242 ;
	7'h3b :
		TR_128 = RG_rl_242 ;
	7'h3c :
		TR_128 = RG_rl_242 ;
	7'h3d :
		TR_128 = RG_rl_242 ;
	7'h3e :
		TR_128 = RG_rl_242 ;
	7'h3f :
		TR_128 = RG_rl_242 ;
	7'h40 :
		TR_128 = RG_rl_242 ;
	7'h41 :
		TR_128 = RG_rl_242 ;
	7'h42 :
		TR_128 = RG_rl_242 ;
	7'h43 :
		TR_128 = RG_rl_242 ;
	7'h44 :
		TR_128 = RG_rl_242 ;
	7'h45 :
		TR_128 = RG_rl_242 ;
	7'h46 :
		TR_128 = RG_rl_242 ;
	7'h47 :
		TR_128 = RG_rl_242 ;
	7'h48 :
		TR_128 = RG_rl_242 ;
	7'h49 :
		TR_128 = RG_rl_242 ;
	7'h4a :
		TR_128 = RG_rl_242 ;
	7'h4b :
		TR_128 = RG_rl_242 ;
	7'h4c :
		TR_128 = RG_rl_242 ;
	7'h4d :
		TR_128 = RG_rl_242 ;
	7'h4e :
		TR_128 = RG_rl_242 ;
	7'h4f :
		TR_128 = RG_rl_242 ;
	7'h50 :
		TR_128 = RG_rl_242 ;
	7'h51 :
		TR_128 = RG_rl_242 ;
	7'h52 :
		TR_128 = RG_rl_242 ;
	7'h53 :
		TR_128 = RG_rl_242 ;
	7'h54 :
		TR_128 = RG_rl_242 ;
	7'h55 :
		TR_128 = RG_rl_242 ;
	7'h56 :
		TR_128 = RG_rl_242 ;
	7'h57 :
		TR_128 = RG_rl_242 ;
	7'h58 :
		TR_128 = RG_rl_242 ;
	7'h59 :
		TR_128 = RG_rl_242 ;
	7'h5a :
		TR_128 = RG_rl_242 ;
	7'h5b :
		TR_128 = RG_rl_242 ;
	7'h5c :
		TR_128 = RG_rl_242 ;
	7'h5d :
		TR_128 = RG_rl_242 ;
	7'h5e :
		TR_128 = RG_rl_242 ;
	7'h5f :
		TR_128 = RG_rl_242 ;
	7'h60 :
		TR_128 = RG_rl_242 ;
	7'h61 :
		TR_128 = RG_rl_242 ;
	7'h62 :
		TR_128 = RG_rl_242 ;
	7'h63 :
		TR_128 = RG_rl_242 ;
	7'h64 :
		TR_128 = RG_rl_242 ;
	7'h65 :
		TR_128 = RG_rl_242 ;
	7'h66 :
		TR_128 = RG_rl_242 ;
	7'h67 :
		TR_128 = RG_rl_242 ;
	7'h68 :
		TR_128 = RG_rl_242 ;
	7'h69 :
		TR_128 = RG_rl_242 ;
	7'h6a :
		TR_128 = RG_rl_242 ;
	7'h6b :
		TR_128 = RG_rl_242 ;
	7'h6c :
		TR_128 = RG_rl_242 ;
	7'h6d :
		TR_128 = RG_rl_242 ;
	7'h6e :
		TR_128 = RG_rl_242 ;
	7'h6f :
		TR_128 = RG_rl_242 ;
	7'h70 :
		TR_128 = RG_rl_242 ;
	7'h71 :
		TR_128 = RG_rl_242 ;
	7'h72 :
		TR_128 = RG_rl_242 ;
	7'h73 :
		TR_128 = RG_rl_242 ;
	7'h74 :
		TR_128 = 9'h000 ;	// line#=../rle.cpp:68
	7'h75 :
		TR_128 = RG_rl_242 ;
	7'h76 :
		TR_128 = RG_rl_242 ;
	7'h77 :
		TR_128 = RG_rl_242 ;
	7'h78 :
		TR_128 = RG_rl_242 ;
	7'h79 :
		TR_128 = RG_rl_242 ;
	7'h7a :
		TR_128 = RG_rl_242 ;
	7'h7b :
		TR_128 = RG_rl_242 ;
	7'h7c :
		TR_128 = RG_rl_242 ;
	7'h7d :
		TR_128 = RG_rl_242 ;
	7'h7e :
		TR_128 = RG_rl_242 ;
	7'h7f :
		TR_128 = RG_rl_242 ;
	default :
		TR_128 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_57 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h01 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h02 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h03 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h04 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h05 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h06 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h07 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h08 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h09 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h0a :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h0b :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h0c :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h0d :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h0e :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h0f :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h10 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h11 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h12 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h13 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h14 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h15 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h16 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h17 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h18 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h19 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h1a :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h1b :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h1c :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h1d :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h1e :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h1f :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h20 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h21 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h22 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h23 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h24 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h25 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h26 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h27 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h28 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h29 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h2a :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h2b :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h2c :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h2d :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h2e :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h2f :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h30 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h31 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h32 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h33 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h34 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h35 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h36 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h37 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h38 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h39 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h3a :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h3b :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h3c :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h3d :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h3e :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h3f :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h40 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h41 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h42 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h43 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h44 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h45 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h46 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h47 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h48 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h49 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h4a :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h4b :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h4c :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h4d :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h4e :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h4f :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h50 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h51 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h52 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h53 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h54 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h55 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h56 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h57 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h58 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h59 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h5a :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h5b :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h5c :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h5d :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h5e :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h5f :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h60 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h61 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h62 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h63 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h64 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h65 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h66 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h67 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h68 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h69 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h6a :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h6b :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h6c :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h6d :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h6e :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h6f :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h70 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h71 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h72 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h73 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h74 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h75 :
		TR_129 = 9'h000 ;	// line#=../rle.cpp:68
	7'h76 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h77 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h78 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h79 :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h7a :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h7b :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h7c :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h7d :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h7e :
		TR_129 = RG_quantized_block_rl_57 ;
	7'h7f :
		TR_129 = RG_quantized_block_rl_57 ;
	default :
		TR_129 = 9'hx ;
	endcase
always @ ( RG_rl_243 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_130 = RG_rl_243 ;
	7'h01 :
		TR_130 = RG_rl_243 ;
	7'h02 :
		TR_130 = RG_rl_243 ;
	7'h03 :
		TR_130 = RG_rl_243 ;
	7'h04 :
		TR_130 = RG_rl_243 ;
	7'h05 :
		TR_130 = RG_rl_243 ;
	7'h06 :
		TR_130 = RG_rl_243 ;
	7'h07 :
		TR_130 = RG_rl_243 ;
	7'h08 :
		TR_130 = RG_rl_243 ;
	7'h09 :
		TR_130 = RG_rl_243 ;
	7'h0a :
		TR_130 = RG_rl_243 ;
	7'h0b :
		TR_130 = RG_rl_243 ;
	7'h0c :
		TR_130 = RG_rl_243 ;
	7'h0d :
		TR_130 = RG_rl_243 ;
	7'h0e :
		TR_130 = RG_rl_243 ;
	7'h0f :
		TR_130 = RG_rl_243 ;
	7'h10 :
		TR_130 = RG_rl_243 ;
	7'h11 :
		TR_130 = RG_rl_243 ;
	7'h12 :
		TR_130 = RG_rl_243 ;
	7'h13 :
		TR_130 = RG_rl_243 ;
	7'h14 :
		TR_130 = RG_rl_243 ;
	7'h15 :
		TR_130 = RG_rl_243 ;
	7'h16 :
		TR_130 = RG_rl_243 ;
	7'h17 :
		TR_130 = RG_rl_243 ;
	7'h18 :
		TR_130 = RG_rl_243 ;
	7'h19 :
		TR_130 = RG_rl_243 ;
	7'h1a :
		TR_130 = RG_rl_243 ;
	7'h1b :
		TR_130 = RG_rl_243 ;
	7'h1c :
		TR_130 = RG_rl_243 ;
	7'h1d :
		TR_130 = RG_rl_243 ;
	7'h1e :
		TR_130 = RG_rl_243 ;
	7'h1f :
		TR_130 = RG_rl_243 ;
	7'h20 :
		TR_130 = RG_rl_243 ;
	7'h21 :
		TR_130 = RG_rl_243 ;
	7'h22 :
		TR_130 = RG_rl_243 ;
	7'h23 :
		TR_130 = RG_rl_243 ;
	7'h24 :
		TR_130 = RG_rl_243 ;
	7'h25 :
		TR_130 = RG_rl_243 ;
	7'h26 :
		TR_130 = RG_rl_243 ;
	7'h27 :
		TR_130 = RG_rl_243 ;
	7'h28 :
		TR_130 = RG_rl_243 ;
	7'h29 :
		TR_130 = RG_rl_243 ;
	7'h2a :
		TR_130 = RG_rl_243 ;
	7'h2b :
		TR_130 = RG_rl_243 ;
	7'h2c :
		TR_130 = RG_rl_243 ;
	7'h2d :
		TR_130 = RG_rl_243 ;
	7'h2e :
		TR_130 = RG_rl_243 ;
	7'h2f :
		TR_130 = RG_rl_243 ;
	7'h30 :
		TR_130 = RG_rl_243 ;
	7'h31 :
		TR_130 = RG_rl_243 ;
	7'h32 :
		TR_130 = RG_rl_243 ;
	7'h33 :
		TR_130 = RG_rl_243 ;
	7'h34 :
		TR_130 = RG_rl_243 ;
	7'h35 :
		TR_130 = RG_rl_243 ;
	7'h36 :
		TR_130 = RG_rl_243 ;
	7'h37 :
		TR_130 = RG_rl_243 ;
	7'h38 :
		TR_130 = RG_rl_243 ;
	7'h39 :
		TR_130 = RG_rl_243 ;
	7'h3a :
		TR_130 = RG_rl_243 ;
	7'h3b :
		TR_130 = RG_rl_243 ;
	7'h3c :
		TR_130 = RG_rl_243 ;
	7'h3d :
		TR_130 = RG_rl_243 ;
	7'h3e :
		TR_130 = RG_rl_243 ;
	7'h3f :
		TR_130 = RG_rl_243 ;
	7'h40 :
		TR_130 = RG_rl_243 ;
	7'h41 :
		TR_130 = RG_rl_243 ;
	7'h42 :
		TR_130 = RG_rl_243 ;
	7'h43 :
		TR_130 = RG_rl_243 ;
	7'h44 :
		TR_130 = RG_rl_243 ;
	7'h45 :
		TR_130 = RG_rl_243 ;
	7'h46 :
		TR_130 = RG_rl_243 ;
	7'h47 :
		TR_130 = RG_rl_243 ;
	7'h48 :
		TR_130 = RG_rl_243 ;
	7'h49 :
		TR_130 = RG_rl_243 ;
	7'h4a :
		TR_130 = RG_rl_243 ;
	7'h4b :
		TR_130 = RG_rl_243 ;
	7'h4c :
		TR_130 = RG_rl_243 ;
	7'h4d :
		TR_130 = RG_rl_243 ;
	7'h4e :
		TR_130 = RG_rl_243 ;
	7'h4f :
		TR_130 = RG_rl_243 ;
	7'h50 :
		TR_130 = RG_rl_243 ;
	7'h51 :
		TR_130 = RG_rl_243 ;
	7'h52 :
		TR_130 = RG_rl_243 ;
	7'h53 :
		TR_130 = RG_rl_243 ;
	7'h54 :
		TR_130 = RG_rl_243 ;
	7'h55 :
		TR_130 = RG_rl_243 ;
	7'h56 :
		TR_130 = RG_rl_243 ;
	7'h57 :
		TR_130 = RG_rl_243 ;
	7'h58 :
		TR_130 = RG_rl_243 ;
	7'h59 :
		TR_130 = RG_rl_243 ;
	7'h5a :
		TR_130 = RG_rl_243 ;
	7'h5b :
		TR_130 = RG_rl_243 ;
	7'h5c :
		TR_130 = RG_rl_243 ;
	7'h5d :
		TR_130 = RG_rl_243 ;
	7'h5e :
		TR_130 = RG_rl_243 ;
	7'h5f :
		TR_130 = RG_rl_243 ;
	7'h60 :
		TR_130 = RG_rl_243 ;
	7'h61 :
		TR_130 = RG_rl_243 ;
	7'h62 :
		TR_130 = RG_rl_243 ;
	7'h63 :
		TR_130 = RG_rl_243 ;
	7'h64 :
		TR_130 = RG_rl_243 ;
	7'h65 :
		TR_130 = RG_rl_243 ;
	7'h66 :
		TR_130 = RG_rl_243 ;
	7'h67 :
		TR_130 = RG_rl_243 ;
	7'h68 :
		TR_130 = RG_rl_243 ;
	7'h69 :
		TR_130 = RG_rl_243 ;
	7'h6a :
		TR_130 = RG_rl_243 ;
	7'h6b :
		TR_130 = RG_rl_243 ;
	7'h6c :
		TR_130 = RG_rl_243 ;
	7'h6d :
		TR_130 = RG_rl_243 ;
	7'h6e :
		TR_130 = RG_rl_243 ;
	7'h6f :
		TR_130 = RG_rl_243 ;
	7'h70 :
		TR_130 = RG_rl_243 ;
	7'h71 :
		TR_130 = RG_rl_243 ;
	7'h72 :
		TR_130 = RG_rl_243 ;
	7'h73 :
		TR_130 = RG_rl_243 ;
	7'h74 :
		TR_130 = RG_rl_243 ;
	7'h75 :
		TR_130 = RG_rl_243 ;
	7'h76 :
		TR_130 = 9'h000 ;	// line#=../rle.cpp:68
	7'h77 :
		TR_130 = RG_rl_243 ;
	7'h78 :
		TR_130 = RG_rl_243 ;
	7'h79 :
		TR_130 = RG_rl_243 ;
	7'h7a :
		TR_130 = RG_rl_243 ;
	7'h7b :
		TR_130 = RG_rl_243 ;
	7'h7c :
		TR_130 = RG_rl_243 ;
	7'h7d :
		TR_130 = RG_rl_243 ;
	7'h7e :
		TR_130 = RG_rl_243 ;
	7'h7f :
		TR_130 = RG_rl_243 ;
	default :
		TR_130 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_58 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h01 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h02 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h03 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h04 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h05 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h06 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h07 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h08 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h09 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h0a :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h0b :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h0c :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h0d :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h0e :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h0f :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h10 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h11 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h12 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h13 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h14 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h15 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h16 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h17 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h18 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h19 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h1a :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h1b :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h1c :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h1d :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h1e :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h1f :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h20 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h21 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h22 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h23 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h24 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h25 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h26 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h27 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h28 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h29 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h2a :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h2b :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h2c :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h2d :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h2e :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h2f :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h30 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h31 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h32 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h33 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h34 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h35 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h36 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h37 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h38 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h39 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h3a :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h3b :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h3c :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h3d :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h3e :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h3f :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h40 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h41 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h42 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h43 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h44 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h45 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h46 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h47 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h48 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h49 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h4a :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h4b :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h4c :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h4d :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h4e :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h4f :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h50 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h51 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h52 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h53 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h54 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h55 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h56 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h57 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h58 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h59 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h5a :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h5b :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h5c :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h5d :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h5e :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h5f :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h60 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h61 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h62 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h63 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h64 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h65 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h66 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h67 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h68 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h69 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h6a :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h6b :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h6c :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h6d :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h6e :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h6f :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h70 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h71 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h72 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h73 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h74 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h75 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h76 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h77 :
		TR_131 = 9'h000 ;	// line#=../rle.cpp:68
	7'h78 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h79 :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h7a :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h7b :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h7c :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h7d :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h7e :
		TR_131 = RG_quantized_block_rl_58 ;
	7'h7f :
		TR_131 = RG_quantized_block_rl_58 ;
	default :
		TR_131 = 9'hx ;
	endcase
always @ ( RG_rl_244 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_132 = RG_rl_244 ;
	7'h01 :
		TR_132 = RG_rl_244 ;
	7'h02 :
		TR_132 = RG_rl_244 ;
	7'h03 :
		TR_132 = RG_rl_244 ;
	7'h04 :
		TR_132 = RG_rl_244 ;
	7'h05 :
		TR_132 = RG_rl_244 ;
	7'h06 :
		TR_132 = RG_rl_244 ;
	7'h07 :
		TR_132 = RG_rl_244 ;
	7'h08 :
		TR_132 = RG_rl_244 ;
	7'h09 :
		TR_132 = RG_rl_244 ;
	7'h0a :
		TR_132 = RG_rl_244 ;
	7'h0b :
		TR_132 = RG_rl_244 ;
	7'h0c :
		TR_132 = RG_rl_244 ;
	7'h0d :
		TR_132 = RG_rl_244 ;
	7'h0e :
		TR_132 = RG_rl_244 ;
	7'h0f :
		TR_132 = RG_rl_244 ;
	7'h10 :
		TR_132 = RG_rl_244 ;
	7'h11 :
		TR_132 = RG_rl_244 ;
	7'h12 :
		TR_132 = RG_rl_244 ;
	7'h13 :
		TR_132 = RG_rl_244 ;
	7'h14 :
		TR_132 = RG_rl_244 ;
	7'h15 :
		TR_132 = RG_rl_244 ;
	7'h16 :
		TR_132 = RG_rl_244 ;
	7'h17 :
		TR_132 = RG_rl_244 ;
	7'h18 :
		TR_132 = RG_rl_244 ;
	7'h19 :
		TR_132 = RG_rl_244 ;
	7'h1a :
		TR_132 = RG_rl_244 ;
	7'h1b :
		TR_132 = RG_rl_244 ;
	7'h1c :
		TR_132 = RG_rl_244 ;
	7'h1d :
		TR_132 = RG_rl_244 ;
	7'h1e :
		TR_132 = RG_rl_244 ;
	7'h1f :
		TR_132 = RG_rl_244 ;
	7'h20 :
		TR_132 = RG_rl_244 ;
	7'h21 :
		TR_132 = RG_rl_244 ;
	7'h22 :
		TR_132 = RG_rl_244 ;
	7'h23 :
		TR_132 = RG_rl_244 ;
	7'h24 :
		TR_132 = RG_rl_244 ;
	7'h25 :
		TR_132 = RG_rl_244 ;
	7'h26 :
		TR_132 = RG_rl_244 ;
	7'h27 :
		TR_132 = RG_rl_244 ;
	7'h28 :
		TR_132 = RG_rl_244 ;
	7'h29 :
		TR_132 = RG_rl_244 ;
	7'h2a :
		TR_132 = RG_rl_244 ;
	7'h2b :
		TR_132 = RG_rl_244 ;
	7'h2c :
		TR_132 = RG_rl_244 ;
	7'h2d :
		TR_132 = RG_rl_244 ;
	7'h2e :
		TR_132 = RG_rl_244 ;
	7'h2f :
		TR_132 = RG_rl_244 ;
	7'h30 :
		TR_132 = RG_rl_244 ;
	7'h31 :
		TR_132 = RG_rl_244 ;
	7'h32 :
		TR_132 = RG_rl_244 ;
	7'h33 :
		TR_132 = RG_rl_244 ;
	7'h34 :
		TR_132 = RG_rl_244 ;
	7'h35 :
		TR_132 = RG_rl_244 ;
	7'h36 :
		TR_132 = RG_rl_244 ;
	7'h37 :
		TR_132 = RG_rl_244 ;
	7'h38 :
		TR_132 = RG_rl_244 ;
	7'h39 :
		TR_132 = RG_rl_244 ;
	7'h3a :
		TR_132 = RG_rl_244 ;
	7'h3b :
		TR_132 = RG_rl_244 ;
	7'h3c :
		TR_132 = RG_rl_244 ;
	7'h3d :
		TR_132 = RG_rl_244 ;
	7'h3e :
		TR_132 = RG_rl_244 ;
	7'h3f :
		TR_132 = RG_rl_244 ;
	7'h40 :
		TR_132 = RG_rl_244 ;
	7'h41 :
		TR_132 = RG_rl_244 ;
	7'h42 :
		TR_132 = RG_rl_244 ;
	7'h43 :
		TR_132 = RG_rl_244 ;
	7'h44 :
		TR_132 = RG_rl_244 ;
	7'h45 :
		TR_132 = RG_rl_244 ;
	7'h46 :
		TR_132 = RG_rl_244 ;
	7'h47 :
		TR_132 = RG_rl_244 ;
	7'h48 :
		TR_132 = RG_rl_244 ;
	7'h49 :
		TR_132 = RG_rl_244 ;
	7'h4a :
		TR_132 = RG_rl_244 ;
	7'h4b :
		TR_132 = RG_rl_244 ;
	7'h4c :
		TR_132 = RG_rl_244 ;
	7'h4d :
		TR_132 = RG_rl_244 ;
	7'h4e :
		TR_132 = RG_rl_244 ;
	7'h4f :
		TR_132 = RG_rl_244 ;
	7'h50 :
		TR_132 = RG_rl_244 ;
	7'h51 :
		TR_132 = RG_rl_244 ;
	7'h52 :
		TR_132 = RG_rl_244 ;
	7'h53 :
		TR_132 = RG_rl_244 ;
	7'h54 :
		TR_132 = RG_rl_244 ;
	7'h55 :
		TR_132 = RG_rl_244 ;
	7'h56 :
		TR_132 = RG_rl_244 ;
	7'h57 :
		TR_132 = RG_rl_244 ;
	7'h58 :
		TR_132 = RG_rl_244 ;
	7'h59 :
		TR_132 = RG_rl_244 ;
	7'h5a :
		TR_132 = RG_rl_244 ;
	7'h5b :
		TR_132 = RG_rl_244 ;
	7'h5c :
		TR_132 = RG_rl_244 ;
	7'h5d :
		TR_132 = RG_rl_244 ;
	7'h5e :
		TR_132 = RG_rl_244 ;
	7'h5f :
		TR_132 = RG_rl_244 ;
	7'h60 :
		TR_132 = RG_rl_244 ;
	7'h61 :
		TR_132 = RG_rl_244 ;
	7'h62 :
		TR_132 = RG_rl_244 ;
	7'h63 :
		TR_132 = RG_rl_244 ;
	7'h64 :
		TR_132 = RG_rl_244 ;
	7'h65 :
		TR_132 = RG_rl_244 ;
	7'h66 :
		TR_132 = RG_rl_244 ;
	7'h67 :
		TR_132 = RG_rl_244 ;
	7'h68 :
		TR_132 = RG_rl_244 ;
	7'h69 :
		TR_132 = RG_rl_244 ;
	7'h6a :
		TR_132 = RG_rl_244 ;
	7'h6b :
		TR_132 = RG_rl_244 ;
	7'h6c :
		TR_132 = RG_rl_244 ;
	7'h6d :
		TR_132 = RG_rl_244 ;
	7'h6e :
		TR_132 = RG_rl_244 ;
	7'h6f :
		TR_132 = RG_rl_244 ;
	7'h70 :
		TR_132 = RG_rl_244 ;
	7'h71 :
		TR_132 = RG_rl_244 ;
	7'h72 :
		TR_132 = RG_rl_244 ;
	7'h73 :
		TR_132 = RG_rl_244 ;
	7'h74 :
		TR_132 = RG_rl_244 ;
	7'h75 :
		TR_132 = RG_rl_244 ;
	7'h76 :
		TR_132 = RG_rl_244 ;
	7'h77 :
		TR_132 = RG_rl_244 ;
	7'h78 :
		TR_132 = 9'h000 ;	// line#=../rle.cpp:68
	7'h79 :
		TR_132 = RG_rl_244 ;
	7'h7a :
		TR_132 = RG_rl_244 ;
	7'h7b :
		TR_132 = RG_rl_244 ;
	7'h7c :
		TR_132 = RG_rl_244 ;
	7'h7d :
		TR_132 = RG_rl_244 ;
	7'h7e :
		TR_132 = RG_rl_244 ;
	7'h7f :
		TR_132 = RG_rl_244 ;
	default :
		TR_132 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_59 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h01 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h02 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h03 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h04 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h05 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h06 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h07 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h08 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h09 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h0a :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h0b :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h0c :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h0d :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h0e :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h0f :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h10 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h11 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h12 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h13 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h14 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h15 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h16 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h17 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h18 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h19 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h1a :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h1b :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h1c :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h1d :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h1e :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h1f :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h20 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h21 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h22 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h23 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h24 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h25 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h26 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h27 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h28 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h29 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h2a :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h2b :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h2c :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h2d :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h2e :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h2f :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h30 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h31 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h32 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h33 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h34 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h35 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h36 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h37 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h38 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h39 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h3a :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h3b :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h3c :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h3d :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h3e :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h3f :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h40 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h41 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h42 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h43 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h44 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h45 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h46 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h47 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h48 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h49 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h4a :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h4b :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h4c :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h4d :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h4e :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h4f :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h50 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h51 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h52 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h53 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h54 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h55 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h56 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h57 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h58 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h59 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h5a :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h5b :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h5c :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h5d :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h5e :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h5f :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h60 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h61 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h62 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h63 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h64 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h65 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h66 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h67 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h68 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h69 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h6a :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h6b :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h6c :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h6d :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h6e :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h6f :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h70 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h71 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h72 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h73 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h74 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h75 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h76 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h77 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h78 :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h79 :
		TR_133 = 9'h000 ;	// line#=../rle.cpp:68
	7'h7a :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h7b :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h7c :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h7d :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h7e :
		TR_133 = RG_quantized_block_rl_59 ;
	7'h7f :
		TR_133 = RG_quantized_block_rl_59 ;
	default :
		TR_133 = 9'hx ;
	endcase
always @ ( RG_rl_245 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_134 = RG_rl_245 ;
	7'h01 :
		TR_134 = RG_rl_245 ;
	7'h02 :
		TR_134 = RG_rl_245 ;
	7'h03 :
		TR_134 = RG_rl_245 ;
	7'h04 :
		TR_134 = RG_rl_245 ;
	7'h05 :
		TR_134 = RG_rl_245 ;
	7'h06 :
		TR_134 = RG_rl_245 ;
	7'h07 :
		TR_134 = RG_rl_245 ;
	7'h08 :
		TR_134 = RG_rl_245 ;
	7'h09 :
		TR_134 = RG_rl_245 ;
	7'h0a :
		TR_134 = RG_rl_245 ;
	7'h0b :
		TR_134 = RG_rl_245 ;
	7'h0c :
		TR_134 = RG_rl_245 ;
	7'h0d :
		TR_134 = RG_rl_245 ;
	7'h0e :
		TR_134 = RG_rl_245 ;
	7'h0f :
		TR_134 = RG_rl_245 ;
	7'h10 :
		TR_134 = RG_rl_245 ;
	7'h11 :
		TR_134 = RG_rl_245 ;
	7'h12 :
		TR_134 = RG_rl_245 ;
	7'h13 :
		TR_134 = RG_rl_245 ;
	7'h14 :
		TR_134 = RG_rl_245 ;
	7'h15 :
		TR_134 = RG_rl_245 ;
	7'h16 :
		TR_134 = RG_rl_245 ;
	7'h17 :
		TR_134 = RG_rl_245 ;
	7'h18 :
		TR_134 = RG_rl_245 ;
	7'h19 :
		TR_134 = RG_rl_245 ;
	7'h1a :
		TR_134 = RG_rl_245 ;
	7'h1b :
		TR_134 = RG_rl_245 ;
	7'h1c :
		TR_134 = RG_rl_245 ;
	7'h1d :
		TR_134 = RG_rl_245 ;
	7'h1e :
		TR_134 = RG_rl_245 ;
	7'h1f :
		TR_134 = RG_rl_245 ;
	7'h20 :
		TR_134 = RG_rl_245 ;
	7'h21 :
		TR_134 = RG_rl_245 ;
	7'h22 :
		TR_134 = RG_rl_245 ;
	7'h23 :
		TR_134 = RG_rl_245 ;
	7'h24 :
		TR_134 = RG_rl_245 ;
	7'h25 :
		TR_134 = RG_rl_245 ;
	7'h26 :
		TR_134 = RG_rl_245 ;
	7'h27 :
		TR_134 = RG_rl_245 ;
	7'h28 :
		TR_134 = RG_rl_245 ;
	7'h29 :
		TR_134 = RG_rl_245 ;
	7'h2a :
		TR_134 = RG_rl_245 ;
	7'h2b :
		TR_134 = RG_rl_245 ;
	7'h2c :
		TR_134 = RG_rl_245 ;
	7'h2d :
		TR_134 = RG_rl_245 ;
	7'h2e :
		TR_134 = RG_rl_245 ;
	7'h2f :
		TR_134 = RG_rl_245 ;
	7'h30 :
		TR_134 = RG_rl_245 ;
	7'h31 :
		TR_134 = RG_rl_245 ;
	7'h32 :
		TR_134 = RG_rl_245 ;
	7'h33 :
		TR_134 = RG_rl_245 ;
	7'h34 :
		TR_134 = RG_rl_245 ;
	7'h35 :
		TR_134 = RG_rl_245 ;
	7'h36 :
		TR_134 = RG_rl_245 ;
	7'h37 :
		TR_134 = RG_rl_245 ;
	7'h38 :
		TR_134 = RG_rl_245 ;
	7'h39 :
		TR_134 = RG_rl_245 ;
	7'h3a :
		TR_134 = RG_rl_245 ;
	7'h3b :
		TR_134 = RG_rl_245 ;
	7'h3c :
		TR_134 = RG_rl_245 ;
	7'h3d :
		TR_134 = RG_rl_245 ;
	7'h3e :
		TR_134 = RG_rl_245 ;
	7'h3f :
		TR_134 = RG_rl_245 ;
	7'h40 :
		TR_134 = RG_rl_245 ;
	7'h41 :
		TR_134 = RG_rl_245 ;
	7'h42 :
		TR_134 = RG_rl_245 ;
	7'h43 :
		TR_134 = RG_rl_245 ;
	7'h44 :
		TR_134 = RG_rl_245 ;
	7'h45 :
		TR_134 = RG_rl_245 ;
	7'h46 :
		TR_134 = RG_rl_245 ;
	7'h47 :
		TR_134 = RG_rl_245 ;
	7'h48 :
		TR_134 = RG_rl_245 ;
	7'h49 :
		TR_134 = RG_rl_245 ;
	7'h4a :
		TR_134 = RG_rl_245 ;
	7'h4b :
		TR_134 = RG_rl_245 ;
	7'h4c :
		TR_134 = RG_rl_245 ;
	7'h4d :
		TR_134 = RG_rl_245 ;
	7'h4e :
		TR_134 = RG_rl_245 ;
	7'h4f :
		TR_134 = RG_rl_245 ;
	7'h50 :
		TR_134 = RG_rl_245 ;
	7'h51 :
		TR_134 = RG_rl_245 ;
	7'h52 :
		TR_134 = RG_rl_245 ;
	7'h53 :
		TR_134 = RG_rl_245 ;
	7'h54 :
		TR_134 = RG_rl_245 ;
	7'h55 :
		TR_134 = RG_rl_245 ;
	7'h56 :
		TR_134 = RG_rl_245 ;
	7'h57 :
		TR_134 = RG_rl_245 ;
	7'h58 :
		TR_134 = RG_rl_245 ;
	7'h59 :
		TR_134 = RG_rl_245 ;
	7'h5a :
		TR_134 = RG_rl_245 ;
	7'h5b :
		TR_134 = RG_rl_245 ;
	7'h5c :
		TR_134 = RG_rl_245 ;
	7'h5d :
		TR_134 = RG_rl_245 ;
	7'h5e :
		TR_134 = RG_rl_245 ;
	7'h5f :
		TR_134 = RG_rl_245 ;
	7'h60 :
		TR_134 = RG_rl_245 ;
	7'h61 :
		TR_134 = RG_rl_245 ;
	7'h62 :
		TR_134 = RG_rl_245 ;
	7'h63 :
		TR_134 = RG_rl_245 ;
	7'h64 :
		TR_134 = RG_rl_245 ;
	7'h65 :
		TR_134 = RG_rl_245 ;
	7'h66 :
		TR_134 = RG_rl_245 ;
	7'h67 :
		TR_134 = RG_rl_245 ;
	7'h68 :
		TR_134 = RG_rl_245 ;
	7'h69 :
		TR_134 = RG_rl_245 ;
	7'h6a :
		TR_134 = RG_rl_245 ;
	7'h6b :
		TR_134 = RG_rl_245 ;
	7'h6c :
		TR_134 = RG_rl_245 ;
	7'h6d :
		TR_134 = RG_rl_245 ;
	7'h6e :
		TR_134 = RG_rl_245 ;
	7'h6f :
		TR_134 = RG_rl_245 ;
	7'h70 :
		TR_134 = RG_rl_245 ;
	7'h71 :
		TR_134 = RG_rl_245 ;
	7'h72 :
		TR_134 = RG_rl_245 ;
	7'h73 :
		TR_134 = RG_rl_245 ;
	7'h74 :
		TR_134 = RG_rl_245 ;
	7'h75 :
		TR_134 = RG_rl_245 ;
	7'h76 :
		TR_134 = RG_rl_245 ;
	7'h77 :
		TR_134 = RG_rl_245 ;
	7'h78 :
		TR_134 = RG_rl_245 ;
	7'h79 :
		TR_134 = RG_rl_245 ;
	7'h7a :
		TR_134 = 9'h000 ;	// line#=../rle.cpp:68
	7'h7b :
		TR_134 = RG_rl_245 ;
	7'h7c :
		TR_134 = RG_rl_245 ;
	7'h7d :
		TR_134 = RG_rl_245 ;
	7'h7e :
		TR_134 = RG_rl_245 ;
	7'h7f :
		TR_134 = RG_rl_245 ;
	default :
		TR_134 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_60 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h01 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h02 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h03 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h04 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h05 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h06 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h07 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h08 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h09 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h0a :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h0b :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h0c :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h0d :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h0e :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h0f :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h10 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h11 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h12 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h13 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h14 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h15 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h16 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h17 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h18 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h19 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h1a :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h1b :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h1c :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h1d :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h1e :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h1f :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h20 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h21 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h22 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h23 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h24 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h25 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h26 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h27 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h28 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h29 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h2a :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h2b :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h2c :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h2d :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h2e :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h2f :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h30 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h31 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h32 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h33 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h34 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h35 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h36 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h37 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h38 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h39 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h3a :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h3b :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h3c :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h3d :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h3e :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h3f :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h40 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h41 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h42 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h43 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h44 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h45 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h46 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h47 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h48 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h49 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h4a :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h4b :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h4c :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h4d :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h4e :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h4f :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h50 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h51 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h52 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h53 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h54 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h55 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h56 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h57 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h58 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h59 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h5a :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h5b :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h5c :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h5d :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h5e :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h5f :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h60 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h61 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h62 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h63 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h64 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h65 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h66 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h67 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h68 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h69 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h6a :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h6b :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h6c :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h6d :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h6e :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h6f :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h70 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h71 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h72 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h73 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h74 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h75 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h76 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h77 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h78 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h79 :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h7a :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h7b :
		TR_135 = 9'h000 ;	// line#=../rle.cpp:68
	7'h7c :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h7d :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h7e :
		TR_135 = RG_quantized_block_rl_60 ;
	7'h7f :
		TR_135 = RG_quantized_block_rl_60 ;
	default :
		TR_135 = 9'hx ;
	endcase
always @ ( RG_rl_246 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_136 = RG_rl_246 ;
	7'h01 :
		TR_136 = RG_rl_246 ;
	7'h02 :
		TR_136 = RG_rl_246 ;
	7'h03 :
		TR_136 = RG_rl_246 ;
	7'h04 :
		TR_136 = RG_rl_246 ;
	7'h05 :
		TR_136 = RG_rl_246 ;
	7'h06 :
		TR_136 = RG_rl_246 ;
	7'h07 :
		TR_136 = RG_rl_246 ;
	7'h08 :
		TR_136 = RG_rl_246 ;
	7'h09 :
		TR_136 = RG_rl_246 ;
	7'h0a :
		TR_136 = RG_rl_246 ;
	7'h0b :
		TR_136 = RG_rl_246 ;
	7'h0c :
		TR_136 = RG_rl_246 ;
	7'h0d :
		TR_136 = RG_rl_246 ;
	7'h0e :
		TR_136 = RG_rl_246 ;
	7'h0f :
		TR_136 = RG_rl_246 ;
	7'h10 :
		TR_136 = RG_rl_246 ;
	7'h11 :
		TR_136 = RG_rl_246 ;
	7'h12 :
		TR_136 = RG_rl_246 ;
	7'h13 :
		TR_136 = RG_rl_246 ;
	7'h14 :
		TR_136 = RG_rl_246 ;
	7'h15 :
		TR_136 = RG_rl_246 ;
	7'h16 :
		TR_136 = RG_rl_246 ;
	7'h17 :
		TR_136 = RG_rl_246 ;
	7'h18 :
		TR_136 = RG_rl_246 ;
	7'h19 :
		TR_136 = RG_rl_246 ;
	7'h1a :
		TR_136 = RG_rl_246 ;
	7'h1b :
		TR_136 = RG_rl_246 ;
	7'h1c :
		TR_136 = RG_rl_246 ;
	7'h1d :
		TR_136 = RG_rl_246 ;
	7'h1e :
		TR_136 = RG_rl_246 ;
	7'h1f :
		TR_136 = RG_rl_246 ;
	7'h20 :
		TR_136 = RG_rl_246 ;
	7'h21 :
		TR_136 = RG_rl_246 ;
	7'h22 :
		TR_136 = RG_rl_246 ;
	7'h23 :
		TR_136 = RG_rl_246 ;
	7'h24 :
		TR_136 = RG_rl_246 ;
	7'h25 :
		TR_136 = RG_rl_246 ;
	7'h26 :
		TR_136 = RG_rl_246 ;
	7'h27 :
		TR_136 = RG_rl_246 ;
	7'h28 :
		TR_136 = RG_rl_246 ;
	7'h29 :
		TR_136 = RG_rl_246 ;
	7'h2a :
		TR_136 = RG_rl_246 ;
	7'h2b :
		TR_136 = RG_rl_246 ;
	7'h2c :
		TR_136 = RG_rl_246 ;
	7'h2d :
		TR_136 = RG_rl_246 ;
	7'h2e :
		TR_136 = RG_rl_246 ;
	7'h2f :
		TR_136 = RG_rl_246 ;
	7'h30 :
		TR_136 = RG_rl_246 ;
	7'h31 :
		TR_136 = RG_rl_246 ;
	7'h32 :
		TR_136 = RG_rl_246 ;
	7'h33 :
		TR_136 = RG_rl_246 ;
	7'h34 :
		TR_136 = RG_rl_246 ;
	7'h35 :
		TR_136 = RG_rl_246 ;
	7'h36 :
		TR_136 = RG_rl_246 ;
	7'h37 :
		TR_136 = RG_rl_246 ;
	7'h38 :
		TR_136 = RG_rl_246 ;
	7'h39 :
		TR_136 = RG_rl_246 ;
	7'h3a :
		TR_136 = RG_rl_246 ;
	7'h3b :
		TR_136 = RG_rl_246 ;
	7'h3c :
		TR_136 = RG_rl_246 ;
	7'h3d :
		TR_136 = RG_rl_246 ;
	7'h3e :
		TR_136 = RG_rl_246 ;
	7'h3f :
		TR_136 = RG_rl_246 ;
	7'h40 :
		TR_136 = RG_rl_246 ;
	7'h41 :
		TR_136 = RG_rl_246 ;
	7'h42 :
		TR_136 = RG_rl_246 ;
	7'h43 :
		TR_136 = RG_rl_246 ;
	7'h44 :
		TR_136 = RG_rl_246 ;
	7'h45 :
		TR_136 = RG_rl_246 ;
	7'h46 :
		TR_136 = RG_rl_246 ;
	7'h47 :
		TR_136 = RG_rl_246 ;
	7'h48 :
		TR_136 = RG_rl_246 ;
	7'h49 :
		TR_136 = RG_rl_246 ;
	7'h4a :
		TR_136 = RG_rl_246 ;
	7'h4b :
		TR_136 = RG_rl_246 ;
	7'h4c :
		TR_136 = RG_rl_246 ;
	7'h4d :
		TR_136 = RG_rl_246 ;
	7'h4e :
		TR_136 = RG_rl_246 ;
	7'h4f :
		TR_136 = RG_rl_246 ;
	7'h50 :
		TR_136 = RG_rl_246 ;
	7'h51 :
		TR_136 = RG_rl_246 ;
	7'h52 :
		TR_136 = RG_rl_246 ;
	7'h53 :
		TR_136 = RG_rl_246 ;
	7'h54 :
		TR_136 = RG_rl_246 ;
	7'h55 :
		TR_136 = RG_rl_246 ;
	7'h56 :
		TR_136 = RG_rl_246 ;
	7'h57 :
		TR_136 = RG_rl_246 ;
	7'h58 :
		TR_136 = RG_rl_246 ;
	7'h59 :
		TR_136 = RG_rl_246 ;
	7'h5a :
		TR_136 = RG_rl_246 ;
	7'h5b :
		TR_136 = RG_rl_246 ;
	7'h5c :
		TR_136 = RG_rl_246 ;
	7'h5d :
		TR_136 = RG_rl_246 ;
	7'h5e :
		TR_136 = RG_rl_246 ;
	7'h5f :
		TR_136 = RG_rl_246 ;
	7'h60 :
		TR_136 = RG_rl_246 ;
	7'h61 :
		TR_136 = RG_rl_246 ;
	7'h62 :
		TR_136 = RG_rl_246 ;
	7'h63 :
		TR_136 = RG_rl_246 ;
	7'h64 :
		TR_136 = RG_rl_246 ;
	7'h65 :
		TR_136 = RG_rl_246 ;
	7'h66 :
		TR_136 = RG_rl_246 ;
	7'h67 :
		TR_136 = RG_rl_246 ;
	7'h68 :
		TR_136 = RG_rl_246 ;
	7'h69 :
		TR_136 = RG_rl_246 ;
	7'h6a :
		TR_136 = RG_rl_246 ;
	7'h6b :
		TR_136 = RG_rl_246 ;
	7'h6c :
		TR_136 = RG_rl_246 ;
	7'h6d :
		TR_136 = RG_rl_246 ;
	7'h6e :
		TR_136 = RG_rl_246 ;
	7'h6f :
		TR_136 = RG_rl_246 ;
	7'h70 :
		TR_136 = RG_rl_246 ;
	7'h71 :
		TR_136 = RG_rl_246 ;
	7'h72 :
		TR_136 = RG_rl_246 ;
	7'h73 :
		TR_136 = RG_rl_246 ;
	7'h74 :
		TR_136 = RG_rl_246 ;
	7'h75 :
		TR_136 = RG_rl_246 ;
	7'h76 :
		TR_136 = RG_rl_246 ;
	7'h77 :
		TR_136 = RG_rl_246 ;
	7'h78 :
		TR_136 = RG_rl_246 ;
	7'h79 :
		TR_136 = RG_rl_246 ;
	7'h7a :
		TR_136 = RG_rl_246 ;
	7'h7b :
		TR_136 = RG_rl_246 ;
	7'h7c :
		TR_136 = 9'h000 ;	// line#=../rle.cpp:68
	7'h7d :
		TR_136 = RG_rl_246 ;
	7'h7e :
		TR_136 = RG_rl_246 ;
	7'h7f :
		TR_136 = RG_rl_246 ;
	default :
		TR_136 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_61 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h01 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h02 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h03 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h04 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h05 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h06 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h07 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h08 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h09 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h0a :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h0b :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h0c :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h0d :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h0e :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h0f :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h10 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h11 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h12 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h13 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h14 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h15 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h16 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h17 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h18 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h19 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h1a :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h1b :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h1c :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h1d :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h1e :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h1f :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h20 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h21 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h22 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h23 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h24 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h25 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h26 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h27 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h28 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h29 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h2a :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h2b :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h2c :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h2d :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h2e :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h2f :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h30 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h31 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h32 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h33 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h34 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h35 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h36 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h37 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h38 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h39 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h3a :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h3b :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h3c :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h3d :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h3e :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h3f :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h40 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h41 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h42 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h43 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h44 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h45 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h46 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h47 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h48 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h49 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h4a :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h4b :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h4c :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h4d :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h4e :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h4f :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h50 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h51 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h52 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h53 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h54 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h55 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h56 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h57 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h58 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h59 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h5a :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h5b :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h5c :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h5d :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h5e :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h5f :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h60 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h61 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h62 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h63 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h64 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h65 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h66 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h67 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h68 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h69 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h6a :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h6b :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h6c :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h6d :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h6e :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h6f :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h70 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h71 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h72 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h73 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h74 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h75 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h76 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h77 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h78 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h79 :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h7a :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h7b :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h7c :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h7d :
		TR_137 = 9'h000 ;	// line#=../rle.cpp:68
	7'h7e :
		TR_137 = RG_quantized_block_rl_61 ;
	7'h7f :
		TR_137 = RG_quantized_block_rl_61 ;
	default :
		TR_137 = 9'hx ;
	endcase
always @ ( RG_previous_dc_rl_1 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h01 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h02 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h03 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h04 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h05 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h06 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h07 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h08 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h09 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h0a :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h0b :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h0c :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h0d :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h0e :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h0f :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h10 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h11 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h12 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h13 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h14 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h15 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h16 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h17 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h18 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h19 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h1a :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h1b :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h1c :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h1d :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h1e :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h1f :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h20 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h21 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h22 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h23 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h24 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h25 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h26 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h27 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h28 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h29 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h2a :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h2b :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h2c :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h2d :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h2e :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h2f :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h30 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h31 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h32 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h33 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h34 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h35 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h36 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h37 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h38 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h39 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h3a :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h3b :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h3c :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h3d :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h3e :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h3f :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h40 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h41 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h42 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h43 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h44 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h45 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h46 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h47 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h48 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h49 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h4a :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h4b :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h4c :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h4d :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h4e :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h4f :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h50 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h51 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h52 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h53 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h54 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h55 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h56 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h57 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h58 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h59 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h5a :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h5b :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h5c :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h5d :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h5e :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h5f :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h60 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h61 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h62 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h63 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h64 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h65 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h66 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h67 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h68 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h69 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h6a :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h6b :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h6c :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h6d :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h6e :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h6f :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h70 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h71 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h72 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h73 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h74 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h75 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h76 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h77 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h78 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h79 :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h7a :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h7b :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h7c :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h7d :
		TR_138 = RG_previous_dc_rl_1 ;
	7'h7e :
		TR_138 = 9'h000 ;	// line#=../rle.cpp:68
	7'h7f :
		TR_138 = RG_previous_dc_rl_1 ;
	default :
		TR_138 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_62 or RG_len )	// line#=../rle.cpp:68
	case ( RG_len [6:0] )
	7'h00 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h01 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h02 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h03 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h04 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h05 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h06 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h07 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h08 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h09 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h0a :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h0b :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h0c :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h0d :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h0e :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h0f :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h10 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h11 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h12 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h13 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h14 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h15 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h16 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h17 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h18 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h19 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h1a :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h1b :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h1c :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h1d :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h1e :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h1f :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h20 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h21 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h22 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h23 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h24 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h25 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h26 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h27 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h28 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h29 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h2a :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h2b :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h2c :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h2d :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h2e :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h2f :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h30 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h31 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h32 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h33 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h34 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h35 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h36 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h37 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h38 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h39 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h3a :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h3b :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h3c :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h3d :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h3e :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h3f :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h40 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h41 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h42 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h43 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h44 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h45 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h46 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h47 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h48 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h49 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h4a :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h4b :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h4c :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h4d :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h4e :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h4f :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h50 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h51 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h52 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h53 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h54 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h55 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h56 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h57 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h58 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h59 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h5a :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h5b :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h5c :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h5d :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h5e :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h5f :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h60 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h61 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h62 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h63 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h64 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h65 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h66 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h67 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h68 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h69 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h6a :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h6b :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h6c :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h6d :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h6e :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h6f :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h70 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h71 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h72 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h73 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h74 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h75 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h76 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h77 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h78 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h79 :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h7a :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h7b :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h7c :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h7d :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h7e :
		TR_11 = RG_quantized_block_rl_62 ;
	7'h7f :
		TR_11 = 9'h000 ;	// line#=../rle.cpp:68
	default :
		TR_11 = 9'hx ;
	endcase
assign	CT_32 = ~|{ RG_i_j_01 [31:7] , ~RG_i_j_01 [6] , RG_i_j_01 [5:0] } ;	// line#=../rle.cpp:66,67
assign	CT_33 = ( M_01_t1 & ( RG_i_k_01 [31] | ( FF_len & ( ~&RG_i_k_01 [3:0] ) ) ) ) ;	// line#=../rle.cpp:61,62
assign	CT_33_port = CT_33 ;
always @ ( TR_12 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a00_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h1 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'h2 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'h3 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'h4 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'h5 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'h6 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'h7 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'h8 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'h9 :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'ha :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'hb :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'hc :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'hd :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'he :
		RG_rl_a00_d9_c0_t = TR_12 ;
	4'hf :
		RG_rl_a00_d9_c0_t = TR_12 ;
	default :
		RG_rl_a00_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a00_d9_c0 <= RG_rl_a00_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a00_d9_c1 <= TR_12 ;
always @ ( TR_13 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'h1 :
		RG_rl_a01_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h2 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'h3 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'h4 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'h5 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'h6 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'h7 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'h8 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'h9 :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'ha :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'hb :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'hc :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'hd :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'he :
		RG_rl_a01_d9_c0_t = TR_13 ;
	4'hf :
		RG_rl_a01_d9_c0_t = TR_13 ;
	default :
		RG_rl_a01_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a01_d9_c0 <= RG_rl_a01_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a01_d9_c1 <= TR_13 ;
always @ ( TR_14 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'h1 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'h2 :
		RG_rl_a02_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h3 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'h4 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'h5 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'h6 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'h7 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'h8 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'h9 :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'ha :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'hb :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'hc :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'hd :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'he :
		RG_rl_a02_d9_c0_t = TR_14 ;
	4'hf :
		RG_rl_a02_d9_c0_t = TR_14 ;
	default :
		RG_rl_a02_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a02_d9_c0 <= RG_rl_a02_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a02_d9_c1 <= TR_14 ;
always @ ( TR_15 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'h1 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'h2 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'h3 :
		RG_rl_a03_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h4 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'h5 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'h6 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'h7 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'h8 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'h9 :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'ha :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'hb :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'hc :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'hd :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'he :
		RG_rl_a03_d9_c0_t = TR_15 ;
	4'hf :
		RG_rl_a03_d9_c0_t = TR_15 ;
	default :
		RG_rl_a03_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a03_d9_c0 <= RG_rl_a03_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a03_d9_c1 <= TR_15 ;
always @ ( TR_16 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'h1 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'h2 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'h3 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'h4 :
		RG_rl_a04_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h5 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'h6 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'h7 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'h8 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'h9 :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'ha :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'hb :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'hc :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'hd :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'he :
		RG_rl_a04_d9_c0_t = TR_16 ;
	4'hf :
		RG_rl_a04_d9_c0_t = TR_16 ;
	default :
		RG_rl_a04_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a04_d9_c0 <= RG_rl_a04_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a04_d9_c1 <= TR_16 ;
always @ ( TR_17 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'h1 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'h2 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'h3 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'h4 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'h5 :
		RG_rl_a05_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h6 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'h7 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'h8 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'h9 :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'ha :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'hb :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'hc :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'hd :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'he :
		RG_rl_a05_d9_c0_t = TR_17 ;
	4'hf :
		RG_rl_a05_d9_c0_t = TR_17 ;
	default :
		RG_rl_a05_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a05_d9_c0 <= RG_rl_a05_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a05_d9_c1 <= TR_17 ;
always @ ( TR_18 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'h1 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'h2 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'h3 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'h4 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'h5 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'h6 :
		RG_rl_a06_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h7 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'h8 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'h9 :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'ha :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'hb :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'hc :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'hd :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'he :
		RG_rl_a06_d9_c0_t = TR_18 ;
	4'hf :
		RG_rl_a06_d9_c0_t = TR_18 ;
	default :
		RG_rl_a06_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a06_d9_c0 <= RG_rl_a06_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a06_d9_c1 <= TR_18 ;
always @ ( TR_19 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'h1 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'h2 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'h3 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'h4 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'h5 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'h6 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'h7 :
		RG_rl_a07_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h8 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'h9 :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'ha :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'hb :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'hc :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'hd :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'he :
		RG_rl_a07_d9_c0_t = TR_19 ;
	4'hf :
		RG_rl_a07_d9_c0_t = TR_19 ;
	default :
		RG_rl_a07_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a07_d9_c0 <= RG_rl_a07_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a07_d9_c1 <= TR_19 ;
always @ ( TR_20 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'h1 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'h2 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'h3 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'h4 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'h5 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'h6 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'h7 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'h8 :
		RG_rl_a08_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h9 :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'ha :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'hb :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'hc :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'hd :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'he :
		RG_rl_a08_d9_c0_t = TR_20 ;
	4'hf :
		RG_rl_a08_d9_c0_t = TR_20 ;
	default :
		RG_rl_a08_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a08_d9_c0 <= RG_rl_a08_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a08_d9_c1 <= TR_20 ;
always @ ( TR_21 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h1 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h2 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h3 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h4 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h5 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h6 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h7 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h8 :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'h9 :
		RG_rl_a09_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'ha :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'hb :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'hc :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'hd :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'he :
		RG_rl_a09_d9_c0_t = TR_21 ;
	4'hf :
		RG_rl_a09_d9_c0_t = TR_21 ;
	default :
		RG_rl_a09_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a09_d9_c0 <= RG_rl_a09_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a09_d9_c1 <= TR_21 ;
always @ ( TR_22 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h1 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h2 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h3 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h4 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h5 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h6 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h7 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h8 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'h9 :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'ha :
		RG_rl_a10_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hb :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'hc :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'hd :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'he :
		RG_rl_a10_d9_c0_t = TR_22 ;
	4'hf :
		RG_rl_a10_d9_c0_t = TR_22 ;
	default :
		RG_rl_a10_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a10_d9_c0 <= RG_rl_a10_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a10_d9_c1 <= TR_22 ;
always @ ( TR_23 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h1 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h2 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h3 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h4 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h5 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h6 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h7 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h8 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'h9 :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'ha :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'hb :
		RG_rl_a11_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hc :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'hd :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'he :
		RG_rl_a11_d9_c0_t = TR_23 ;
	4'hf :
		RG_rl_a11_d9_c0_t = TR_23 ;
	default :
		RG_rl_a11_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a11_d9_c0 <= RG_rl_a11_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a11_d9_c1 <= TR_23 ;
always @ ( TR_24 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h1 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h2 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h3 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h4 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h5 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h6 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h7 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h8 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'h9 :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'ha :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'hb :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'hc :
		RG_rl_a12_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hd :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'he :
		RG_rl_a12_d9_c0_t = TR_24 ;
	4'hf :
		RG_rl_a12_d9_c0_t = TR_24 ;
	default :
		RG_rl_a12_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a12_d9_c0 <= RG_rl_a12_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a12_d9_c1 <= TR_24 ;
always @ ( TR_25 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h1 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h2 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h3 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h4 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h5 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h6 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h7 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h8 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'h9 :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'ha :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'hb :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'hc :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'hd :
		RG_rl_a13_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'he :
		RG_rl_a13_d9_c0_t = TR_25 ;
	4'hf :
		RG_rl_a13_d9_c0_t = TR_25 ;
	default :
		RG_rl_a13_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a13_d9_c0 <= RG_rl_a13_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a13_d9_c1 <= TR_25 ;
always @ ( TR_26 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h1 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h2 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h3 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h4 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h5 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h6 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h7 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h8 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'h9 :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'ha :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'hb :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'hc :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'hd :
		RG_rl_a14_d9_c0_t = TR_26 ;
	4'he :
		RG_rl_a14_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hf :
		RG_rl_a14_d9_c0_t = TR_26 ;
	default :
		RG_rl_a14_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a14_d9_c0 <= RG_rl_a14_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a14_d9_c1 <= TR_26 ;
always @ ( TR_27 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h1 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h2 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h3 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h4 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h5 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h6 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h7 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h8 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'h9 :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'ha :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'hb :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'hc :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'hd :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'he :
		RG_rl_a15_d9_c0_t = TR_27 ;
	4'hf :
		RG_rl_a15_d9_c0_t = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_rl_a15_d9_c0_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a15_d9_c0 <= RG_rl_a15_d9_c0_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a15_d9_c1 <= TR_27 ;
always @ ( posedge clk )
	RG_rl_a16_d9_c0 <= TR_28 ;
always @ ( TR_28 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a16_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h1 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'h2 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'h3 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'h4 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'h5 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'h6 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'h7 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'h8 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'h9 :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'ha :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'hb :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'hc :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'hd :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'he :
		RG_rl_a16_d9_c1_t = TR_28 ;
	4'hf :
		RG_rl_a16_d9_c1_t = TR_28 ;
	default :
		RG_rl_a16_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a16_d9_c1 <= RG_rl_a16_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a17_d9_c0 <= TR_29 ;
always @ ( TR_29 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'h1 :
		RG_rl_a17_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h2 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'h3 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'h4 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'h5 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'h6 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'h7 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'h8 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'h9 :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'ha :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'hb :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'hc :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'hd :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'he :
		RG_rl_a17_d9_c1_t = TR_29 ;
	4'hf :
		RG_rl_a17_d9_c1_t = TR_29 ;
	default :
		RG_rl_a17_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a17_d9_c1 <= RG_rl_a17_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a18_d9_c0 <= TR_30 ;
always @ ( TR_30 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'h1 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'h2 :
		RG_rl_a18_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h3 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'h4 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'h5 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'h6 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'h7 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'h8 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'h9 :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'ha :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'hb :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'hc :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'hd :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'he :
		RG_rl_a18_d9_c1_t = TR_30 ;
	4'hf :
		RG_rl_a18_d9_c1_t = TR_30 ;
	default :
		RG_rl_a18_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a18_d9_c1 <= RG_rl_a18_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a19_d9_c0 <= TR_31 ;
always @ ( TR_31 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'h1 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'h2 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'h3 :
		RG_rl_a19_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h4 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'h5 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'h6 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'h7 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'h8 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'h9 :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'ha :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'hb :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'hc :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'hd :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'he :
		RG_rl_a19_d9_c1_t = TR_31 ;
	4'hf :
		RG_rl_a19_d9_c1_t = TR_31 ;
	default :
		RG_rl_a19_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a19_d9_c1 <= RG_rl_a19_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a20_d9_c0 <= TR_32 ;
always @ ( TR_32 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'h1 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'h2 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'h3 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'h4 :
		RG_rl_a20_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h5 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'h6 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'h7 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'h8 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'h9 :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'ha :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'hb :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'hc :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'hd :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'he :
		RG_rl_a20_d9_c1_t = TR_32 ;
	4'hf :
		RG_rl_a20_d9_c1_t = TR_32 ;
	default :
		RG_rl_a20_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a20_d9_c1 <= RG_rl_a20_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a21_d9_c0 <= TR_33 ;
always @ ( TR_33 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'h1 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'h2 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'h3 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'h4 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'h5 :
		RG_rl_a21_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h6 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'h7 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'h8 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'h9 :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'ha :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'hb :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'hc :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'hd :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'he :
		RG_rl_a21_d9_c1_t = TR_33 ;
	4'hf :
		RG_rl_a21_d9_c1_t = TR_33 ;
	default :
		RG_rl_a21_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a21_d9_c1 <= RG_rl_a21_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a22_d9_c0 <= TR_34 ;
always @ ( TR_34 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'h1 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'h2 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'h3 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'h4 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'h5 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'h6 :
		RG_rl_a22_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h7 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'h8 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'h9 :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'ha :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'hb :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'hc :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'hd :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'he :
		RG_rl_a22_d9_c1_t = TR_34 ;
	4'hf :
		RG_rl_a22_d9_c1_t = TR_34 ;
	default :
		RG_rl_a22_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a22_d9_c1 <= RG_rl_a22_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a23_d9_c0 <= TR_35 ;
always @ ( TR_35 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'h1 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'h2 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'h3 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'h4 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'h5 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'h6 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'h7 :
		RG_rl_a23_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h8 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'h9 :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'ha :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'hb :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'hc :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'hd :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'he :
		RG_rl_a23_d9_c1_t = TR_35 ;
	4'hf :
		RG_rl_a23_d9_c1_t = TR_35 ;
	default :
		RG_rl_a23_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a23_d9_c1 <= RG_rl_a23_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a24_d9_c0 <= TR_36 ;
always @ ( TR_36 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'h1 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'h2 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'h3 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'h4 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'h5 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'h6 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'h7 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'h8 :
		RG_rl_a24_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h9 :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'ha :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'hb :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'hc :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'hd :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'he :
		RG_rl_a24_d9_c1_t = TR_36 ;
	4'hf :
		RG_rl_a24_d9_c1_t = TR_36 ;
	default :
		RG_rl_a24_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a24_d9_c1 <= RG_rl_a24_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a25_d9_c0 <= TR_37 ;
always @ ( TR_37 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h1 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h2 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h3 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h4 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h5 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h6 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h7 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h8 :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'h9 :
		RG_rl_a25_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'ha :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'hb :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'hc :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'hd :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'he :
		RG_rl_a25_d9_c1_t = TR_37 ;
	4'hf :
		RG_rl_a25_d9_c1_t = TR_37 ;
	default :
		RG_rl_a25_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a25_d9_c1 <= RG_rl_a25_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a26_d9_c0 <= TR_38 ;
always @ ( TR_38 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h1 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h2 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h3 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h4 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h5 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h6 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h7 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h8 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'h9 :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'ha :
		RG_rl_a26_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hb :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'hc :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'hd :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'he :
		RG_rl_a26_d9_c1_t = TR_38 ;
	4'hf :
		RG_rl_a26_d9_c1_t = TR_38 ;
	default :
		RG_rl_a26_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a26_d9_c1 <= RG_rl_a26_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a27_d9_c0 <= TR_39 ;
always @ ( TR_39 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h1 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h2 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h3 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h4 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h5 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h6 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h7 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h8 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'h9 :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'ha :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'hb :
		RG_rl_a27_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hc :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'hd :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'he :
		RG_rl_a27_d9_c1_t = TR_39 ;
	4'hf :
		RG_rl_a27_d9_c1_t = TR_39 ;
	default :
		RG_rl_a27_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a27_d9_c1 <= RG_rl_a27_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a28_d9_c0 <= TR_40 ;
always @ ( TR_40 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h1 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h2 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h3 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h4 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h5 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h6 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h7 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h8 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'h9 :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'ha :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'hb :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'hc :
		RG_rl_a28_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hd :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'he :
		RG_rl_a28_d9_c1_t = TR_40 ;
	4'hf :
		RG_rl_a28_d9_c1_t = TR_40 ;
	default :
		RG_rl_a28_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a28_d9_c1 <= RG_rl_a28_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a29_d9_c0 <= TR_41 ;
always @ ( TR_41 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h1 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h2 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h3 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h4 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h5 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h6 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h7 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h8 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'h9 :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'ha :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'hb :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'hc :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'hd :
		RG_rl_a29_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'he :
		RG_rl_a29_d9_c1_t = TR_41 ;
	4'hf :
		RG_rl_a29_d9_c1_t = TR_41 ;
	default :
		RG_rl_a29_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a29_d9_c1 <= RG_rl_a29_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a30_d9_c0 <= TR_42 ;
always @ ( TR_42 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h1 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h2 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h3 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h4 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h5 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h6 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h7 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h8 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'h9 :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'ha :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'hb :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'hc :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'hd :
		RG_rl_a30_d9_c1_t = TR_42 ;
	4'he :
		RG_rl_a30_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hf :
		RG_rl_a30_d9_c1_t = TR_42 ;
	default :
		RG_rl_a30_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a30_d9_c1 <= RG_rl_a30_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a31_d9_c0 <= TR_43 ;
always @ ( TR_43 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h1 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h2 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h3 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h4 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h5 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h6 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h7 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h8 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'h9 :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'ha :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'hb :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'hc :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'hd :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'he :
		RG_rl_a31_d9_c1_t = TR_43 ;
	4'hf :
		RG_rl_a31_d9_c1_t = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_rl_a31_d9_c1_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a31_d9_c1 <= RG_rl_a31_d9_c1_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a32_d9_c0 <= TR_44 ;
always @ ( TR_44 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a32_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h1 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'h2 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'h3 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'h4 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'h5 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'h6 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'h7 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'h8 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'h9 :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'ha :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'hb :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'hc :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'hd :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'he :
		RG_rl_a32_d9_c2_t = TR_44 ;
	4'hf :
		RG_rl_a32_d9_c2_t = TR_44 ;
	default :
		RG_rl_a32_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a32_d9_c2 <= RG_rl_a32_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a33_d9_c0 <= TR_45 ;
always @ ( TR_45 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'h1 :
		RG_rl_a33_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h2 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'h3 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'h4 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'h5 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'h6 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'h7 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'h8 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'h9 :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'ha :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'hb :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'hc :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'hd :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'he :
		RG_rl_a33_d9_c2_t = TR_45 ;
	4'hf :
		RG_rl_a33_d9_c2_t = TR_45 ;
	default :
		RG_rl_a33_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a33_d9_c2 <= RG_rl_a33_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a34_d9_c0 <= TR_46 ;
always @ ( TR_46 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'h1 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'h2 :
		RG_rl_a34_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h3 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'h4 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'h5 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'h6 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'h7 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'h8 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'h9 :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'ha :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'hb :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'hc :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'hd :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'he :
		RG_rl_a34_d9_c2_t = TR_46 ;
	4'hf :
		RG_rl_a34_d9_c2_t = TR_46 ;
	default :
		RG_rl_a34_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a34_d9_c2 <= RG_rl_a34_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a35_d9_c0 <= TR_47 ;
always @ ( TR_47 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'h1 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'h2 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'h3 :
		RG_rl_a35_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h4 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'h5 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'h6 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'h7 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'h8 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'h9 :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'ha :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'hb :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'hc :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'hd :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'he :
		RG_rl_a35_d9_c2_t = TR_47 ;
	4'hf :
		RG_rl_a35_d9_c2_t = TR_47 ;
	default :
		RG_rl_a35_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a35_d9_c2 <= RG_rl_a35_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a36_d9_c0 <= TR_48 ;
always @ ( TR_48 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'h1 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'h2 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'h3 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'h4 :
		RG_rl_a36_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h5 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'h6 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'h7 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'h8 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'h9 :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'ha :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'hb :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'hc :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'hd :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'he :
		RG_rl_a36_d9_c2_t = TR_48 ;
	4'hf :
		RG_rl_a36_d9_c2_t = TR_48 ;
	default :
		RG_rl_a36_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a36_d9_c2 <= RG_rl_a36_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a37_d9_c0 <= TR_49 ;
always @ ( TR_49 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'h1 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'h2 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'h3 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'h4 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'h5 :
		RG_rl_a37_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h6 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'h7 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'h8 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'h9 :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'ha :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'hb :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'hc :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'hd :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'he :
		RG_rl_a37_d9_c2_t = TR_49 ;
	4'hf :
		RG_rl_a37_d9_c2_t = TR_49 ;
	default :
		RG_rl_a37_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a37_d9_c2 <= RG_rl_a37_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a38_d9_c0 <= TR_50 ;
always @ ( TR_50 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'h1 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'h2 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'h3 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'h4 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'h5 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'h6 :
		RG_rl_a38_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h7 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'h8 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'h9 :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'ha :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'hb :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'hc :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'hd :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'he :
		RG_rl_a38_d9_c2_t = TR_50 ;
	4'hf :
		RG_rl_a38_d9_c2_t = TR_50 ;
	default :
		RG_rl_a38_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a38_d9_c2 <= RG_rl_a38_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a39_d9_c0 <= TR_51 ;
always @ ( TR_51 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'h1 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'h2 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'h3 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'h4 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'h5 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'h6 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'h7 :
		RG_rl_a39_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h8 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'h9 :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'ha :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'hb :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'hc :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'hd :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'he :
		RG_rl_a39_d9_c2_t = TR_51 ;
	4'hf :
		RG_rl_a39_d9_c2_t = TR_51 ;
	default :
		RG_rl_a39_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a39_d9_c2 <= RG_rl_a39_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a40_d9_c0 <= TR_52 ;
always @ ( TR_52 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'h1 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'h2 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'h3 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'h4 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'h5 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'h6 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'h7 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'h8 :
		RG_rl_a40_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h9 :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'ha :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'hb :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'hc :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'hd :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'he :
		RG_rl_a40_d9_c2_t = TR_52 ;
	4'hf :
		RG_rl_a40_d9_c2_t = TR_52 ;
	default :
		RG_rl_a40_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a40_d9_c2 <= RG_rl_a40_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a41_d9_c0 <= TR_53 ;
always @ ( TR_53 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h1 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h2 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h3 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h4 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h5 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h6 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h7 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h8 :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'h9 :
		RG_rl_a41_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'ha :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'hb :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'hc :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'hd :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'he :
		RG_rl_a41_d9_c2_t = TR_53 ;
	4'hf :
		RG_rl_a41_d9_c2_t = TR_53 ;
	default :
		RG_rl_a41_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a41_d9_c2 <= RG_rl_a41_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a42_d9_c0 <= TR_54 ;
always @ ( TR_54 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h1 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h2 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h3 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h4 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h5 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h6 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h7 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h8 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'h9 :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'ha :
		RG_rl_a42_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hb :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'hc :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'hd :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'he :
		RG_rl_a42_d9_c2_t = TR_54 ;
	4'hf :
		RG_rl_a42_d9_c2_t = TR_54 ;
	default :
		RG_rl_a42_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a42_d9_c2 <= RG_rl_a42_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a43_d9_c0 <= TR_55 ;
always @ ( TR_55 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h1 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h2 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h3 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h4 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h5 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h6 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h7 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h8 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'h9 :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'ha :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'hb :
		RG_rl_a43_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hc :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'hd :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'he :
		RG_rl_a43_d9_c2_t = TR_55 ;
	4'hf :
		RG_rl_a43_d9_c2_t = TR_55 ;
	default :
		RG_rl_a43_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a43_d9_c2 <= RG_rl_a43_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a44_d9_c0 <= TR_56 ;
always @ ( TR_56 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h1 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h2 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h3 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h4 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h5 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h6 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h7 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h8 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'h9 :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'ha :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'hb :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'hc :
		RG_rl_a44_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hd :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'he :
		RG_rl_a44_d9_c2_t = TR_56 ;
	4'hf :
		RG_rl_a44_d9_c2_t = TR_56 ;
	default :
		RG_rl_a44_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a44_d9_c2 <= RG_rl_a44_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a45_d9_c0 <= TR_57 ;
always @ ( TR_57 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h1 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h2 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h3 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h4 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h5 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h6 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h7 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h8 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'h9 :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'ha :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'hb :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'hc :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'hd :
		RG_rl_a45_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'he :
		RG_rl_a45_d9_c2_t = TR_57 ;
	4'hf :
		RG_rl_a45_d9_c2_t = TR_57 ;
	default :
		RG_rl_a45_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a45_d9_c2 <= RG_rl_a45_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a46_d9_c0 <= TR_58 ;
always @ ( TR_58 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h1 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h2 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h3 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h4 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h5 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h6 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h7 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h8 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'h9 :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'ha :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'hb :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'hc :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'hd :
		RG_rl_a46_d9_c2_t = TR_58 ;
	4'he :
		RG_rl_a46_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hf :
		RG_rl_a46_d9_c2_t = TR_58 ;
	default :
		RG_rl_a46_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a46_d9_c2 <= RG_rl_a46_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a47_d9_c0 <= TR_59 ;
always @ ( TR_59 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h1 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h2 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h3 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h4 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h5 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h6 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h7 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h8 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'h9 :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'ha :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'hb :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'hc :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'hd :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'he :
		RG_rl_a47_d9_c2_t = TR_59 ;
	4'hf :
		RG_rl_a47_d9_c2_t = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_rl_a47_d9_c2_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a47_d9_c2 <= RG_rl_a47_d9_c2_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a48_d9_c0 <= TR_60 ;
always @ ( TR_60 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a48_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h1 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'h2 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'h3 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'h4 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'h5 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'h6 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'h7 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'h8 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'h9 :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'ha :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'hb :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'hc :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'hd :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'he :
		RG_rl_a48_d9_c3_t = TR_60 ;
	4'hf :
		RG_rl_a48_d9_c3_t = TR_60 ;
	default :
		RG_rl_a48_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a48_d9_c3 <= RG_rl_a48_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a49_d9_c0 <= TR_61 ;
always @ ( TR_61 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'h1 :
		RG_rl_a49_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h2 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'h3 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'h4 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'h5 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'h6 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'h7 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'h8 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'h9 :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'ha :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'hb :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'hc :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'hd :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'he :
		RG_rl_a49_d9_c3_t = TR_61 ;
	4'hf :
		RG_rl_a49_d9_c3_t = TR_61 ;
	default :
		RG_rl_a49_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a49_d9_c3 <= RG_rl_a49_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a50_d9_c0 <= TR_62 ;
always @ ( TR_62 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'h1 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'h2 :
		RG_rl_a50_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h3 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'h4 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'h5 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'h6 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'h7 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'h8 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'h9 :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'ha :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'hb :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'hc :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'hd :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'he :
		RG_rl_a50_d9_c3_t = TR_62 ;
	4'hf :
		RG_rl_a50_d9_c3_t = TR_62 ;
	default :
		RG_rl_a50_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a50_d9_c3 <= RG_rl_a50_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a51_d9_c0 <= TR_63 ;
always @ ( TR_63 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'h1 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'h2 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'h3 :
		RG_rl_a51_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h4 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'h5 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'h6 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'h7 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'h8 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'h9 :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'ha :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'hb :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'hc :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'hd :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'he :
		RG_rl_a51_d9_c3_t = TR_63 ;
	4'hf :
		RG_rl_a51_d9_c3_t = TR_63 ;
	default :
		RG_rl_a51_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a51_d9_c3 <= RG_rl_a51_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a52_d9_c0 <= TR_64 ;
always @ ( TR_64 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'h1 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'h2 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'h3 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'h4 :
		RG_rl_a52_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h5 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'h6 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'h7 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'h8 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'h9 :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'ha :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'hb :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'hc :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'hd :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'he :
		RG_rl_a52_d9_c3_t = TR_64 ;
	4'hf :
		RG_rl_a52_d9_c3_t = TR_64 ;
	default :
		RG_rl_a52_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a52_d9_c3 <= RG_rl_a52_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a53_d9_c0 <= TR_65 ;
always @ ( TR_65 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'h1 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'h2 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'h3 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'h4 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'h5 :
		RG_rl_a53_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h6 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'h7 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'h8 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'h9 :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'ha :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'hb :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'hc :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'hd :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'he :
		RG_rl_a53_d9_c3_t = TR_65 ;
	4'hf :
		RG_rl_a53_d9_c3_t = TR_65 ;
	default :
		RG_rl_a53_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a53_d9_c3 <= RG_rl_a53_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a54_d9_c0 <= TR_66 ;
always @ ( TR_66 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'h1 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'h2 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'h3 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'h4 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'h5 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'h6 :
		RG_rl_a54_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h7 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'h8 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'h9 :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'ha :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'hb :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'hc :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'hd :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'he :
		RG_rl_a54_d9_c3_t = TR_66 ;
	4'hf :
		RG_rl_a54_d9_c3_t = TR_66 ;
	default :
		RG_rl_a54_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a54_d9_c3 <= RG_rl_a54_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a55_d9_c0 <= TR_67 ;
always @ ( TR_67 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'h1 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'h2 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'h3 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'h4 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'h5 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'h6 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'h7 :
		RG_rl_a55_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h8 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'h9 :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'ha :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'hb :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'hc :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'hd :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'he :
		RG_rl_a55_d9_c3_t = TR_67 ;
	4'hf :
		RG_rl_a55_d9_c3_t = TR_67 ;
	default :
		RG_rl_a55_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a55_d9_c3 <= RG_rl_a55_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a56_d9_c0 <= TR_68 ;
always @ ( TR_68 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'h1 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'h2 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'h3 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'h4 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'h5 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'h6 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'h7 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'h8 :
		RG_rl_a56_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h9 :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'ha :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'hb :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'hc :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'hd :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'he :
		RG_rl_a56_d9_c3_t = TR_68 ;
	4'hf :
		RG_rl_a56_d9_c3_t = TR_68 ;
	default :
		RG_rl_a56_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a56_d9_c3 <= RG_rl_a56_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a57_d9_c0 <= TR_69 ;
always @ ( TR_69 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h1 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h2 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h3 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h4 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h5 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h6 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h7 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h8 :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'h9 :
		RG_rl_a57_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'ha :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'hb :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'hc :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'hd :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'he :
		RG_rl_a57_d9_c3_t = TR_69 ;
	4'hf :
		RG_rl_a57_d9_c3_t = TR_69 ;
	default :
		RG_rl_a57_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a57_d9_c3 <= RG_rl_a57_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a58_d9_c0 <= TR_70 ;
always @ ( TR_70 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h1 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h2 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h3 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h4 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h5 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h6 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h7 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h8 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'h9 :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'ha :
		RG_rl_a58_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hb :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'hc :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'hd :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'he :
		RG_rl_a58_d9_c3_t = TR_70 ;
	4'hf :
		RG_rl_a58_d9_c3_t = TR_70 ;
	default :
		RG_rl_a58_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a58_d9_c3 <= RG_rl_a58_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a59_d9_c0 <= TR_71 ;
always @ ( TR_71 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h1 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h2 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h3 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h4 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h5 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h6 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h7 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h8 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'h9 :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'ha :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'hb :
		RG_rl_a59_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hc :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'hd :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'he :
		RG_rl_a59_d9_c3_t = TR_71 ;
	4'hf :
		RG_rl_a59_d9_c3_t = TR_71 ;
	default :
		RG_rl_a59_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a59_d9_c3 <= RG_rl_a59_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a60_d9_c0 <= TR_72 ;
always @ ( TR_72 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h1 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h2 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h3 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h4 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h5 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h6 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h7 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h8 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'h9 :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'ha :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'hb :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'hc :
		RG_rl_a60_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hd :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'he :
		RG_rl_a60_d9_c3_t = TR_72 ;
	4'hf :
		RG_rl_a60_d9_c3_t = TR_72 ;
	default :
		RG_rl_a60_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a60_d9_c3 <= RG_rl_a60_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a61_d9_c0 <= TR_73 ;
always @ ( TR_73 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h1 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h2 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h3 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h4 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h5 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h6 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h7 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h8 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'h9 :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'ha :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'hb :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'hc :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'hd :
		RG_rl_a61_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'he :
		RG_rl_a61_d9_c3_t = TR_73 ;
	4'hf :
		RG_rl_a61_d9_c3_t = TR_73 ;
	default :
		RG_rl_a61_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a61_d9_c3 <= RG_rl_a61_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a62_d9_c0 <= TR_74 ;
always @ ( TR_74 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h1 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h2 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h3 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h4 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h5 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h6 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h7 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h8 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'h9 :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'ha :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'hb :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'hc :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'hd :
		RG_rl_a62_d9_c3_t = TR_74 ;
	4'he :
		RG_rl_a62_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hf :
		RG_rl_a62_d9_c3_t = TR_74 ;
	default :
		RG_rl_a62_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a62_d9_c3 <= RG_rl_a62_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a63_d9_c0 <= TR_75 ;
always @ ( TR_75 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h1 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h2 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h3 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h4 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h5 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h6 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h7 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h8 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'h9 :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'ha :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'hb :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'hc :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'hd :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'he :
		RG_rl_a63_d9_c3_t = TR_75 ;
	4'hf :
		RG_rl_a63_d9_c3_t = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_rl_a63_d9_c3_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a63_d9_c3 <= RG_rl_a63_d9_c3_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a64_d9_c0 <= TR_76 ;
always @ ( TR_76 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a64_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h1 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'h2 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'h3 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'h4 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'h5 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'h6 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'h7 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'h8 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'h9 :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'ha :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'hb :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'hc :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'hd :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'he :
		RG_rl_a64_d9_c4_t = TR_76 ;
	4'hf :
		RG_rl_a64_d9_c4_t = TR_76 ;
	default :
		RG_rl_a64_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a64_d9_c4 <= RG_rl_a64_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a65_d9_c0 <= TR_77 ;
always @ ( TR_77 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'h1 :
		RG_rl_a65_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h2 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'h3 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'h4 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'h5 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'h6 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'h7 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'h8 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'h9 :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'ha :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'hb :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'hc :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'hd :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'he :
		RG_rl_a65_d9_c4_t = TR_77 ;
	4'hf :
		RG_rl_a65_d9_c4_t = TR_77 ;
	default :
		RG_rl_a65_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a65_d9_c4 <= RG_rl_a65_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a66_d9_c0 <= TR_78 ;
always @ ( TR_78 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'h1 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'h2 :
		RG_rl_a66_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h3 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'h4 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'h5 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'h6 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'h7 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'h8 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'h9 :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'ha :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'hb :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'hc :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'hd :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'he :
		RG_rl_a66_d9_c4_t = TR_78 ;
	4'hf :
		RG_rl_a66_d9_c4_t = TR_78 ;
	default :
		RG_rl_a66_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a66_d9_c4 <= RG_rl_a66_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a67_d9_c0 <= TR_79 ;
always @ ( TR_79 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'h1 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'h2 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'h3 :
		RG_rl_a67_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h4 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'h5 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'h6 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'h7 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'h8 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'h9 :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'ha :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'hb :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'hc :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'hd :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'he :
		RG_rl_a67_d9_c4_t = TR_79 ;
	4'hf :
		RG_rl_a67_d9_c4_t = TR_79 ;
	default :
		RG_rl_a67_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a67_d9_c4 <= RG_rl_a67_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a68_d9_c0 <= TR_80 ;
always @ ( TR_80 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'h1 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'h2 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'h3 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'h4 :
		RG_rl_a68_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h5 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'h6 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'h7 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'h8 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'h9 :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'ha :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'hb :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'hc :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'hd :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'he :
		RG_rl_a68_d9_c4_t = TR_80 ;
	4'hf :
		RG_rl_a68_d9_c4_t = TR_80 ;
	default :
		RG_rl_a68_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a68_d9_c4 <= RG_rl_a68_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a69_d9_c0 <= TR_81 ;
always @ ( TR_81 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'h1 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'h2 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'h3 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'h4 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'h5 :
		RG_rl_a69_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h6 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'h7 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'h8 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'h9 :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'ha :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'hb :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'hc :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'hd :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'he :
		RG_rl_a69_d9_c4_t = TR_81 ;
	4'hf :
		RG_rl_a69_d9_c4_t = TR_81 ;
	default :
		RG_rl_a69_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a69_d9_c4 <= RG_rl_a69_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a70_d9_c0 <= TR_82 ;
always @ ( TR_82 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'h1 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'h2 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'h3 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'h4 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'h5 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'h6 :
		RG_rl_a70_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h7 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'h8 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'h9 :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'ha :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'hb :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'hc :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'hd :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'he :
		RG_rl_a70_d9_c4_t = TR_82 ;
	4'hf :
		RG_rl_a70_d9_c4_t = TR_82 ;
	default :
		RG_rl_a70_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a70_d9_c4 <= RG_rl_a70_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a71_d9_c0 <= TR_83 ;
always @ ( TR_83 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'h1 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'h2 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'h3 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'h4 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'h5 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'h6 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'h7 :
		RG_rl_a71_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h8 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'h9 :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'ha :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'hb :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'hc :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'hd :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'he :
		RG_rl_a71_d9_c4_t = TR_83 ;
	4'hf :
		RG_rl_a71_d9_c4_t = TR_83 ;
	default :
		RG_rl_a71_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a71_d9_c4 <= RG_rl_a71_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a72_d9_c0 <= TR_84 ;
always @ ( TR_84 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'h1 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'h2 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'h3 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'h4 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'h5 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'h6 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'h7 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'h8 :
		RG_rl_a72_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h9 :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'ha :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'hb :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'hc :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'hd :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'he :
		RG_rl_a72_d9_c4_t = TR_84 ;
	4'hf :
		RG_rl_a72_d9_c4_t = TR_84 ;
	default :
		RG_rl_a72_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a72_d9_c4 <= RG_rl_a72_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a73_d9_c0 <= TR_85 ;
always @ ( TR_85 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h1 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h2 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h3 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h4 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h5 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h6 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h7 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h8 :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'h9 :
		RG_rl_a73_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'ha :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'hb :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'hc :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'hd :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'he :
		RG_rl_a73_d9_c4_t = TR_85 ;
	4'hf :
		RG_rl_a73_d9_c4_t = TR_85 ;
	default :
		RG_rl_a73_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a73_d9_c4 <= RG_rl_a73_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a74_d9_c0 <= TR_86 ;
always @ ( TR_86 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h1 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h2 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h3 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h4 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h5 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h6 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h7 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h8 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'h9 :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'ha :
		RG_rl_a74_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hb :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'hc :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'hd :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'he :
		RG_rl_a74_d9_c4_t = TR_86 ;
	4'hf :
		RG_rl_a74_d9_c4_t = TR_86 ;
	default :
		RG_rl_a74_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a74_d9_c4 <= RG_rl_a74_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a75_d9_c0 <= TR_87 ;
always @ ( TR_87 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h1 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h2 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h3 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h4 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h5 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h6 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h7 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h8 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'h9 :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'ha :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'hb :
		RG_rl_a75_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hc :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'hd :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'he :
		RG_rl_a75_d9_c4_t = TR_87 ;
	4'hf :
		RG_rl_a75_d9_c4_t = TR_87 ;
	default :
		RG_rl_a75_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a75_d9_c4 <= RG_rl_a75_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a76_d9_c0 <= TR_88 ;
always @ ( TR_88 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h1 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h2 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h3 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h4 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h5 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h6 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h7 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h8 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'h9 :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'ha :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'hb :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'hc :
		RG_rl_a76_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hd :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'he :
		RG_rl_a76_d9_c4_t = TR_88 ;
	4'hf :
		RG_rl_a76_d9_c4_t = TR_88 ;
	default :
		RG_rl_a76_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a76_d9_c4 <= RG_rl_a76_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a77_d9_c0 <= TR_89 ;
always @ ( TR_89 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h1 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h2 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h3 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h4 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h5 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h6 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h7 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h8 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'h9 :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'ha :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'hb :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'hc :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'hd :
		RG_rl_a77_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'he :
		RG_rl_a77_d9_c4_t = TR_89 ;
	4'hf :
		RG_rl_a77_d9_c4_t = TR_89 ;
	default :
		RG_rl_a77_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a77_d9_c4 <= RG_rl_a77_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a78_d9_c0 <= TR_90 ;
always @ ( TR_90 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h1 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h2 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h3 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h4 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h5 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h6 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h7 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h8 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'h9 :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'ha :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'hb :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'hc :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'hd :
		RG_rl_a78_d9_c4_t = TR_90 ;
	4'he :
		RG_rl_a78_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hf :
		RG_rl_a78_d9_c4_t = TR_90 ;
	default :
		RG_rl_a78_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a78_d9_c4 <= RG_rl_a78_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a79_d9_c0 <= TR_91 ;
always @ ( TR_91 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h1 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h2 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h3 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h4 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h5 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h6 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h7 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h8 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'h9 :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'ha :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'hb :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'hc :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'hd :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'he :
		RG_rl_a79_d9_c4_t = TR_91 ;
	4'hf :
		RG_rl_a79_d9_c4_t = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_rl_a79_d9_c4_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a79_d9_c4 <= RG_rl_a79_d9_c4_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a80_d9_c0 <= TR_92 ;
always @ ( TR_92 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a80_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h1 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'h2 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'h3 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'h4 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'h5 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'h6 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'h7 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'h8 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'h9 :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'ha :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'hb :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'hc :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'hd :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'he :
		RG_rl_a80_d9_c5_t = TR_92 ;
	4'hf :
		RG_rl_a80_d9_c5_t = TR_92 ;
	default :
		RG_rl_a80_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a80_d9_c5 <= RG_rl_a80_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a81_d9_c0 <= TR_93 ;
always @ ( TR_93 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'h1 :
		RG_rl_a81_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h2 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'h3 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'h4 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'h5 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'h6 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'h7 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'h8 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'h9 :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'ha :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'hb :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'hc :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'hd :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'he :
		RG_rl_a81_d9_c5_t = TR_93 ;
	4'hf :
		RG_rl_a81_d9_c5_t = TR_93 ;
	default :
		RG_rl_a81_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a81_d9_c5 <= RG_rl_a81_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a82_d9_c0 <= TR_94 ;
always @ ( TR_94 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'h1 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'h2 :
		RG_rl_a82_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h3 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'h4 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'h5 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'h6 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'h7 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'h8 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'h9 :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'ha :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'hb :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'hc :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'hd :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'he :
		RG_rl_a82_d9_c5_t = TR_94 ;
	4'hf :
		RG_rl_a82_d9_c5_t = TR_94 ;
	default :
		RG_rl_a82_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a82_d9_c5 <= RG_rl_a82_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a83_d9_c0 <= TR_95 ;
always @ ( TR_95 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'h1 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'h2 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'h3 :
		RG_rl_a83_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h4 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'h5 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'h6 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'h7 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'h8 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'h9 :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'ha :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'hb :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'hc :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'hd :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'he :
		RG_rl_a83_d9_c5_t = TR_95 ;
	4'hf :
		RG_rl_a83_d9_c5_t = TR_95 ;
	default :
		RG_rl_a83_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a83_d9_c5 <= RG_rl_a83_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a84_d9_c0 <= TR_96 ;
always @ ( TR_96 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'h1 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'h2 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'h3 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'h4 :
		RG_rl_a84_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h5 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'h6 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'h7 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'h8 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'h9 :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'ha :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'hb :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'hc :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'hd :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'he :
		RG_rl_a84_d9_c5_t = TR_96 ;
	4'hf :
		RG_rl_a84_d9_c5_t = TR_96 ;
	default :
		RG_rl_a84_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a84_d9_c5 <= RG_rl_a84_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a85_d9_c0 <= TR_97 ;
always @ ( TR_97 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'h1 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'h2 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'h3 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'h4 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'h5 :
		RG_rl_a85_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h6 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'h7 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'h8 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'h9 :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'ha :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'hb :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'hc :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'hd :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'he :
		RG_rl_a85_d9_c5_t = TR_97 ;
	4'hf :
		RG_rl_a85_d9_c5_t = TR_97 ;
	default :
		RG_rl_a85_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a85_d9_c5 <= RG_rl_a85_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a86_d9_c0 <= TR_98 ;
always @ ( TR_98 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'h1 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'h2 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'h3 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'h4 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'h5 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'h6 :
		RG_rl_a86_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h7 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'h8 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'h9 :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'ha :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'hb :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'hc :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'hd :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'he :
		RG_rl_a86_d9_c5_t = TR_98 ;
	4'hf :
		RG_rl_a86_d9_c5_t = TR_98 ;
	default :
		RG_rl_a86_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a86_d9_c5 <= RG_rl_a86_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a87_d9_c0 <= TR_99 ;
always @ ( TR_99 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'h1 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'h2 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'h3 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'h4 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'h5 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'h6 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'h7 :
		RG_rl_a87_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h8 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'h9 :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'ha :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'hb :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'hc :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'hd :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'he :
		RG_rl_a87_d9_c5_t = TR_99 ;
	4'hf :
		RG_rl_a87_d9_c5_t = TR_99 ;
	default :
		RG_rl_a87_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a87_d9_c5 <= RG_rl_a87_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a88_d9_c0 <= TR_100 ;
always @ ( TR_100 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'h1 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'h2 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'h3 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'h4 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'h5 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'h6 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'h7 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'h8 :
		RG_rl_a88_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h9 :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'ha :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'hb :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'hc :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'hd :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'he :
		RG_rl_a88_d9_c5_t = TR_100 ;
	4'hf :
		RG_rl_a88_d9_c5_t = TR_100 ;
	default :
		RG_rl_a88_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a88_d9_c5 <= RG_rl_a88_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a89_d9_c0 <= TR_101 ;
always @ ( TR_101 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h1 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h2 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h3 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h4 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h5 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h6 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h7 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h8 :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'h9 :
		RG_rl_a89_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'ha :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'hb :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'hc :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'hd :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'he :
		RG_rl_a89_d9_c5_t = TR_101 ;
	4'hf :
		RG_rl_a89_d9_c5_t = TR_101 ;
	default :
		RG_rl_a89_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a89_d9_c5 <= RG_rl_a89_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a90_d9_c0 <= TR_102 ;
always @ ( TR_102 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h1 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h2 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h3 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h4 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h5 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h6 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h7 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h8 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'h9 :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'ha :
		RG_rl_a90_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hb :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'hc :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'hd :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'he :
		RG_rl_a90_d9_c5_t = TR_102 ;
	4'hf :
		RG_rl_a90_d9_c5_t = TR_102 ;
	default :
		RG_rl_a90_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a90_d9_c5 <= RG_rl_a90_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a91_d9_c0 <= TR_103 ;
always @ ( TR_103 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h1 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h2 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h3 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h4 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h5 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h6 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h7 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h8 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'h9 :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'ha :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'hb :
		RG_rl_a91_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hc :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'hd :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'he :
		RG_rl_a91_d9_c5_t = TR_103 ;
	4'hf :
		RG_rl_a91_d9_c5_t = TR_103 ;
	default :
		RG_rl_a91_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a91_d9_c5 <= RG_rl_a91_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a92_d9_c0 <= TR_104 ;
always @ ( TR_104 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h1 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h2 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h3 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h4 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h5 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h6 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h7 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h8 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'h9 :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'ha :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'hb :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'hc :
		RG_rl_a92_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hd :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'he :
		RG_rl_a92_d9_c5_t = TR_104 ;
	4'hf :
		RG_rl_a92_d9_c5_t = TR_104 ;
	default :
		RG_rl_a92_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a92_d9_c5 <= RG_rl_a92_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a93_d9_c0 <= TR_105 ;
always @ ( TR_105 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h1 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h2 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h3 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h4 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h5 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h6 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h7 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h8 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'h9 :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'ha :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'hb :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'hc :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'hd :
		RG_rl_a93_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'he :
		RG_rl_a93_d9_c5_t = TR_105 ;
	4'hf :
		RG_rl_a93_d9_c5_t = TR_105 ;
	default :
		RG_rl_a93_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a93_d9_c5 <= RG_rl_a93_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a94_d9_c0 <= TR_106 ;
always @ ( TR_106 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h1 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h2 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h3 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h4 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h5 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h6 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h7 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h8 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'h9 :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'ha :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'hb :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'hc :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'hd :
		RG_rl_a94_d9_c5_t = TR_106 ;
	4'he :
		RG_rl_a94_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hf :
		RG_rl_a94_d9_c5_t = TR_106 ;
	default :
		RG_rl_a94_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a94_d9_c5 <= RG_rl_a94_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a95_d9_c0 <= TR_107 ;
always @ ( TR_107 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h1 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h2 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h3 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h4 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h5 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h6 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h7 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h8 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'h9 :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'ha :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'hb :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'hc :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'hd :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'he :
		RG_rl_a95_d9_c5_t = TR_107 ;
	4'hf :
		RG_rl_a95_d9_c5_t = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_rl_a95_d9_c5_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a95_d9_c5 <= RG_rl_a95_d9_c5_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a96_d9_c0 <= TR_108 ;
always @ ( TR_108 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a96_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h1 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'h2 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'h3 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'h4 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'h5 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'h6 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'h7 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'h8 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'h9 :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'ha :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'hb :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'hc :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'hd :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'he :
		RG_rl_a96_d9_c6_t = TR_108 ;
	4'hf :
		RG_rl_a96_d9_c6_t = TR_108 ;
	default :
		RG_rl_a96_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a96_d9_c6 <= RG_rl_a96_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a97_d9_c0 <= TR_109 ;
always @ ( TR_109 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'h1 :
		RG_rl_a97_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h2 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'h3 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'h4 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'h5 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'h6 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'h7 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'h8 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'h9 :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'ha :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'hb :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'hc :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'hd :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'he :
		RG_rl_a97_d9_c6_t = TR_109 ;
	4'hf :
		RG_rl_a97_d9_c6_t = TR_109 ;
	default :
		RG_rl_a97_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a97_d9_c6 <= RG_rl_a97_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a98_d9_c0 <= TR_110 ;
always @ ( TR_110 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'h1 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'h2 :
		RG_rl_a98_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h3 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'h4 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'h5 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'h6 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'h7 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'h8 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'h9 :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'ha :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'hb :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'hc :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'hd :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'he :
		RG_rl_a98_d9_c6_t = TR_110 ;
	4'hf :
		RG_rl_a98_d9_c6_t = TR_110 ;
	default :
		RG_rl_a98_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a98_d9_c6 <= RG_rl_a98_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a99_d9_c0 <= TR_111 ;
always @ ( TR_111 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'h1 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'h2 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'h3 :
		RG_rl_a99_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h4 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'h5 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'h6 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'h7 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'h8 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'h9 :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'ha :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'hb :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'hc :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'hd :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'he :
		RG_rl_a99_d9_c6_t = TR_111 ;
	4'hf :
		RG_rl_a99_d9_c6_t = TR_111 ;
	default :
		RG_rl_a99_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a99_d9_c6 <= RG_rl_a99_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a100_d9_c0 <= TR_112 ;
always @ ( TR_112 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'h1 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'h2 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'h3 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'h4 :
		RG_rl_a100_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h5 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'h6 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'h7 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'h8 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'h9 :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'ha :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'hb :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'hc :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'hd :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'he :
		RG_rl_a100_d9_c6_t = TR_112 ;
	4'hf :
		RG_rl_a100_d9_c6_t = TR_112 ;
	default :
		RG_rl_a100_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a100_d9_c6 <= RG_rl_a100_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a101_d9_c0 <= TR_113 ;
always @ ( TR_113 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'h1 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'h2 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'h3 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'h4 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'h5 :
		RG_rl_a101_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h6 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'h7 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'h8 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'h9 :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'ha :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'hb :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'hc :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'hd :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'he :
		RG_rl_a101_d9_c6_t = TR_113 ;
	4'hf :
		RG_rl_a101_d9_c6_t = TR_113 ;
	default :
		RG_rl_a101_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a101_d9_c6 <= RG_rl_a101_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a102_d9_c0 <= TR_114 ;
always @ ( TR_114 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'h1 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'h2 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'h3 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'h4 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'h5 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'h6 :
		RG_rl_a102_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h7 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'h8 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'h9 :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'ha :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'hb :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'hc :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'hd :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'he :
		RG_rl_a102_d9_c6_t = TR_114 ;
	4'hf :
		RG_rl_a102_d9_c6_t = TR_114 ;
	default :
		RG_rl_a102_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a102_d9_c6 <= RG_rl_a102_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a103_d9_c0 <= TR_115 ;
always @ ( TR_115 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'h1 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'h2 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'h3 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'h4 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'h5 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'h6 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'h7 :
		RG_rl_a103_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h8 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'h9 :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'ha :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'hb :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'hc :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'hd :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'he :
		RG_rl_a103_d9_c6_t = TR_115 ;
	4'hf :
		RG_rl_a103_d9_c6_t = TR_115 ;
	default :
		RG_rl_a103_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a103_d9_c6 <= RG_rl_a103_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a104_d9_c0 <= TR_116 ;
always @ ( TR_116 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'h1 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'h2 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'h3 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'h4 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'h5 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'h6 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'h7 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'h8 :
		RG_rl_a104_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h9 :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'ha :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'hb :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'hc :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'hd :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'he :
		RG_rl_a104_d9_c6_t = TR_116 ;
	4'hf :
		RG_rl_a104_d9_c6_t = TR_116 ;
	default :
		RG_rl_a104_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a104_d9_c6 <= RG_rl_a104_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a105_d9_c0 <= TR_117 ;
always @ ( TR_117 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h1 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h2 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h3 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h4 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h5 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h6 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h7 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h8 :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'h9 :
		RG_rl_a105_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'ha :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'hb :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'hc :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'hd :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'he :
		RG_rl_a105_d9_c6_t = TR_117 ;
	4'hf :
		RG_rl_a105_d9_c6_t = TR_117 ;
	default :
		RG_rl_a105_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a105_d9_c6 <= RG_rl_a105_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a106_d9_c0 <= TR_118 ;
always @ ( TR_118 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h1 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h2 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h3 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h4 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h5 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h6 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h7 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h8 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'h9 :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'ha :
		RG_rl_a106_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hb :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'hc :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'hd :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'he :
		RG_rl_a106_d9_c6_t = TR_118 ;
	4'hf :
		RG_rl_a106_d9_c6_t = TR_118 ;
	default :
		RG_rl_a106_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a106_d9_c6 <= RG_rl_a106_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a107_d9_c0 <= TR_119 ;
always @ ( TR_119 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h1 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h2 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h3 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h4 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h5 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h6 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h7 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h8 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'h9 :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'ha :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'hb :
		RG_rl_a107_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hc :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'hd :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'he :
		RG_rl_a107_d9_c6_t = TR_119 ;
	4'hf :
		RG_rl_a107_d9_c6_t = TR_119 ;
	default :
		RG_rl_a107_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a107_d9_c6 <= RG_rl_a107_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a108_d9_c0 <= TR_120 ;
always @ ( TR_120 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h1 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h2 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h3 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h4 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h5 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h6 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h7 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h8 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'h9 :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'ha :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'hb :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'hc :
		RG_rl_a108_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hd :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'he :
		RG_rl_a108_d9_c6_t = TR_120 ;
	4'hf :
		RG_rl_a108_d9_c6_t = TR_120 ;
	default :
		RG_rl_a108_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a108_d9_c6 <= RG_rl_a108_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a109_d9_c0 <= TR_121 ;
always @ ( TR_121 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h1 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h2 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h3 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h4 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h5 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h6 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h7 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h8 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'h9 :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'ha :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'hb :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'hc :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'hd :
		RG_rl_a109_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'he :
		RG_rl_a109_d9_c6_t = TR_121 ;
	4'hf :
		RG_rl_a109_d9_c6_t = TR_121 ;
	default :
		RG_rl_a109_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a109_d9_c6 <= RG_rl_a109_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a110_d9_c0 <= TR_122 ;
always @ ( TR_122 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h1 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h2 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h3 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h4 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h5 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h6 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h7 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h8 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'h9 :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'ha :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'hb :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'hc :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'hd :
		RG_rl_a110_d9_c6_t = TR_122 ;
	4'he :
		RG_rl_a110_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hf :
		RG_rl_a110_d9_c6_t = TR_122 ;
	default :
		RG_rl_a110_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a110_d9_c6 <= RG_rl_a110_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a111_d9_c0 <= TR_123 ;
always @ ( TR_123 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h1 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h2 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h3 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h4 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h5 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h6 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h7 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h8 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'h9 :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'ha :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'hb :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'hc :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'hd :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'he :
		RG_rl_a111_d9_c6_t = TR_123 ;
	4'hf :
		RG_rl_a111_d9_c6_t = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_rl_a111_d9_c6_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a111_d9_c6 <= RG_rl_a111_d9_c6_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a112_d9_c0 <= TR_124 ;
always @ ( TR_124 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a112_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h1 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'h2 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'h3 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'h4 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'h5 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'h6 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'h7 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'h8 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'h9 :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'ha :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'hb :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'hc :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'hd :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'he :
		RG_rl_a112_d9_c7_t = TR_124 ;
	4'hf :
		RG_rl_a112_d9_c7_t = TR_124 ;
	default :
		RG_rl_a112_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a112_d9_c7 <= RG_rl_a112_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a113_d9_c0 <= TR_125 ;
always @ ( TR_125 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'h1 :
		RG_rl_a113_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h2 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'h3 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'h4 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'h5 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'h6 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'h7 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'h8 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'h9 :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'ha :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'hb :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'hc :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'hd :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'he :
		RG_rl_a113_d9_c7_t = TR_125 ;
	4'hf :
		RG_rl_a113_d9_c7_t = TR_125 ;
	default :
		RG_rl_a113_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a113_d9_c7 <= RG_rl_a113_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a114_d9_c0 <= TR_126 ;
always @ ( TR_126 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'h1 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'h2 :
		RG_rl_a114_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h3 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'h4 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'h5 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'h6 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'h7 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'h8 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'h9 :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'ha :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'hb :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'hc :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'hd :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'he :
		RG_rl_a114_d9_c7_t = TR_126 ;
	4'hf :
		RG_rl_a114_d9_c7_t = TR_126 ;
	default :
		RG_rl_a114_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a114_d9_c7 <= RG_rl_a114_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a115_d9_c0 <= TR_127 ;
always @ ( TR_127 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'h1 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'h2 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'h3 :
		RG_rl_a115_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h4 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'h5 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'h6 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'h7 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'h8 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'h9 :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'ha :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'hb :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'hc :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'hd :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'he :
		RG_rl_a115_d9_c7_t = TR_127 ;
	4'hf :
		RG_rl_a115_d9_c7_t = TR_127 ;
	default :
		RG_rl_a115_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a115_d9_c7 <= RG_rl_a115_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a116_d9_c0 <= TR_128 ;
always @ ( TR_128 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'h1 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'h2 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'h3 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'h4 :
		RG_rl_a116_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h5 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'h6 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'h7 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'h8 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'h9 :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'ha :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'hb :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'hc :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'hd :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'he :
		RG_rl_a116_d9_c7_t = TR_128 ;
	4'hf :
		RG_rl_a116_d9_c7_t = TR_128 ;
	default :
		RG_rl_a116_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a116_d9_c7 <= RG_rl_a116_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a117_d9_c0 <= TR_129 ;
always @ ( TR_129 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'h1 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'h2 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'h3 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'h4 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'h5 :
		RG_rl_a117_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h6 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'h7 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'h8 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'h9 :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'ha :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'hb :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'hc :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'hd :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'he :
		RG_rl_a117_d9_c7_t = TR_129 ;
	4'hf :
		RG_rl_a117_d9_c7_t = TR_129 ;
	default :
		RG_rl_a117_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a117_d9_c7 <= RG_rl_a117_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a118_d9_c0 <= TR_130 ;
always @ ( TR_130 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'h1 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'h2 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'h3 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'h4 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'h5 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'h6 :
		RG_rl_a118_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h7 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'h8 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'h9 :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'ha :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'hb :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'hc :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'hd :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'he :
		RG_rl_a118_d9_c7_t = TR_130 ;
	4'hf :
		RG_rl_a118_d9_c7_t = TR_130 ;
	default :
		RG_rl_a118_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a118_d9_c7 <= RG_rl_a118_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a119_d9_c0 <= TR_131 ;
always @ ( TR_131 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'h1 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'h2 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'h3 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'h4 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'h5 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'h6 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'h7 :
		RG_rl_a119_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h8 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'h9 :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'ha :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'hb :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'hc :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'hd :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'he :
		RG_rl_a119_d9_c7_t = TR_131 ;
	4'hf :
		RG_rl_a119_d9_c7_t = TR_131 ;
	default :
		RG_rl_a119_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a119_d9_c7 <= RG_rl_a119_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a120_d9_c0 <= TR_132 ;
always @ ( TR_132 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'h1 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'h2 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'h3 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'h4 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'h5 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'h6 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'h7 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'h8 :
		RG_rl_a120_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'h9 :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'ha :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'hb :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'hc :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'hd :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'he :
		RG_rl_a120_d9_c7_t = TR_132 ;
	4'hf :
		RG_rl_a120_d9_c7_t = TR_132 ;
	default :
		RG_rl_a120_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a120_d9_c7 <= RG_rl_a120_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a121_d9_c0 <= TR_133 ;
always @ ( TR_133 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h1 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h2 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h3 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h4 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h5 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h6 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h7 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h8 :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'h9 :
		RG_rl_a121_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'ha :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'hb :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'hc :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'hd :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'he :
		RG_rl_a121_d9_c7_t = TR_133 ;
	4'hf :
		RG_rl_a121_d9_c7_t = TR_133 ;
	default :
		RG_rl_a121_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a121_d9_c7 <= RG_rl_a121_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a122_d9_c0 <= TR_134 ;
always @ ( TR_134 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h1 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h2 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h3 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h4 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h5 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h6 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h7 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h8 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'h9 :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'ha :
		RG_rl_a122_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hb :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'hc :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'hd :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'he :
		RG_rl_a122_d9_c7_t = TR_134 ;
	4'hf :
		RG_rl_a122_d9_c7_t = TR_134 ;
	default :
		RG_rl_a122_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a122_d9_c7 <= RG_rl_a122_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a123_d9_c0 <= TR_135 ;
always @ ( TR_135 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h1 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h2 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h3 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h4 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h5 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h6 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h7 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h8 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'h9 :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'ha :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'hb :
		RG_rl_a123_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hc :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'hd :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'he :
		RG_rl_a123_d9_c7_t = TR_135 ;
	4'hf :
		RG_rl_a123_d9_c7_t = TR_135 ;
	default :
		RG_rl_a123_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a123_d9_c7 <= RG_rl_a123_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a124_d9_c0 <= TR_136 ;
always @ ( TR_136 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h1 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h2 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h3 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h4 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h5 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h6 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h7 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h8 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'h9 :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'ha :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'hb :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'hc :
		RG_rl_a124_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hd :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'he :
		RG_rl_a124_d9_c7_t = TR_136 ;
	4'hf :
		RG_rl_a124_d9_c7_t = TR_136 ;
	default :
		RG_rl_a124_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a124_d9_c7 <= RG_rl_a124_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a125_d9_c0 <= TR_137 ;
always @ ( TR_137 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h1 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h2 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h3 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h4 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h5 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h6 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h7 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h8 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'h9 :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'ha :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'hb :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'hc :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'hd :
		RG_rl_a125_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'he :
		RG_rl_a125_d9_c7_t = TR_137 ;
	4'hf :
		RG_rl_a125_d9_c7_t = TR_137 ;
	default :
		RG_rl_a125_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a125_d9_c7 <= RG_rl_a125_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a126_d9_c0 <= TR_138 ;
always @ ( TR_138 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h1 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h2 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h3 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h4 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h5 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h6 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h7 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h8 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'h9 :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'ha :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'hb :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'hc :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'hd :
		RG_rl_a126_d9_c7_t = TR_138 ;
	4'he :
		RG_rl_a126_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	4'hf :
		RG_rl_a126_d9_c7_t = TR_138 ;
	default :
		RG_rl_a126_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a126_d9_c7 <= RG_rl_a126_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( posedge clk )
	RG_rl_a127_d9_c0 <= TR_11 ;
always @ ( TR_11 or incr8u1ot )	// line#=../rle.cpp:68,69
	case ( incr8u1ot [3:0] )
	4'h0 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h1 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h2 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h3 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h4 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h5 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h6 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h7 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h8 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'h9 :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'ha :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'hb :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'hc :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'hd :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'he :
		RG_rl_a127_d9_c7_t = TR_11 ;
	4'hf :
		RG_rl_a127_d9_c7_t = 9'h000 ;	// line#=../rle.cpp:69
	default :
		RG_rl_a127_d9_c7_t = 9'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:68,69
	RG_rl_a127_d9_c7 <= RG_rl_a127_d9_c7_t ;	// line#=../rle.cpp:69
always @ ( RG_rl_a00_d9_c1 or RG_rl_a00_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a00_t5 = RG_rl_a00_d9_c0 ;
	3'h1 :
		rl_a00_t5 = RG_rl_a00_d9_c1 ;
	3'h2 :
		rl_a00_t5 = RG_rl_a00_d9_c1 ;
	3'h3 :
		rl_a00_t5 = RG_rl_a00_d9_c1 ;
	3'h4 :
		rl_a00_t5 = RG_rl_a00_d9_c1 ;
	3'h5 :
		rl_a00_t5 = RG_rl_a00_d9_c1 ;
	3'h6 :
		rl_a00_t5 = RG_rl_a00_d9_c1 ;
	3'h7 :
		rl_a00_t5 = RG_rl_a00_d9_c1 ;
	default :
		rl_a00_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a01_d9_c1 or RG_rl_a01_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a01_t5 = RG_rl_a01_d9_c0 ;
	3'h1 :
		rl_a01_t5 = RG_rl_a01_d9_c1 ;
	3'h2 :
		rl_a01_t5 = RG_rl_a01_d9_c1 ;
	3'h3 :
		rl_a01_t5 = RG_rl_a01_d9_c1 ;
	3'h4 :
		rl_a01_t5 = RG_rl_a01_d9_c1 ;
	3'h5 :
		rl_a01_t5 = RG_rl_a01_d9_c1 ;
	3'h6 :
		rl_a01_t5 = RG_rl_a01_d9_c1 ;
	3'h7 :
		rl_a01_t5 = RG_rl_a01_d9_c1 ;
	default :
		rl_a01_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a02_d9_c1 or RG_rl_a02_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a02_t5 = RG_rl_a02_d9_c0 ;
	3'h1 :
		rl_a02_t5 = RG_rl_a02_d9_c1 ;
	3'h2 :
		rl_a02_t5 = RG_rl_a02_d9_c1 ;
	3'h3 :
		rl_a02_t5 = RG_rl_a02_d9_c1 ;
	3'h4 :
		rl_a02_t5 = RG_rl_a02_d9_c1 ;
	3'h5 :
		rl_a02_t5 = RG_rl_a02_d9_c1 ;
	3'h6 :
		rl_a02_t5 = RG_rl_a02_d9_c1 ;
	3'h7 :
		rl_a02_t5 = RG_rl_a02_d9_c1 ;
	default :
		rl_a02_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a03_d9_c1 or RG_rl_a03_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a03_t5 = RG_rl_a03_d9_c0 ;
	3'h1 :
		rl_a03_t5 = RG_rl_a03_d9_c1 ;
	3'h2 :
		rl_a03_t5 = RG_rl_a03_d9_c1 ;
	3'h3 :
		rl_a03_t5 = RG_rl_a03_d9_c1 ;
	3'h4 :
		rl_a03_t5 = RG_rl_a03_d9_c1 ;
	3'h5 :
		rl_a03_t5 = RG_rl_a03_d9_c1 ;
	3'h6 :
		rl_a03_t5 = RG_rl_a03_d9_c1 ;
	3'h7 :
		rl_a03_t5 = RG_rl_a03_d9_c1 ;
	default :
		rl_a03_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a04_d9_c1 or RG_rl_a04_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a04_t5 = RG_rl_a04_d9_c0 ;
	3'h1 :
		rl_a04_t5 = RG_rl_a04_d9_c1 ;
	3'h2 :
		rl_a04_t5 = RG_rl_a04_d9_c1 ;
	3'h3 :
		rl_a04_t5 = RG_rl_a04_d9_c1 ;
	3'h4 :
		rl_a04_t5 = RG_rl_a04_d9_c1 ;
	3'h5 :
		rl_a04_t5 = RG_rl_a04_d9_c1 ;
	3'h6 :
		rl_a04_t5 = RG_rl_a04_d9_c1 ;
	3'h7 :
		rl_a04_t5 = RG_rl_a04_d9_c1 ;
	default :
		rl_a04_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a05_d9_c1 or RG_rl_a05_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a05_t5 = RG_rl_a05_d9_c0 ;
	3'h1 :
		rl_a05_t5 = RG_rl_a05_d9_c1 ;
	3'h2 :
		rl_a05_t5 = RG_rl_a05_d9_c1 ;
	3'h3 :
		rl_a05_t5 = RG_rl_a05_d9_c1 ;
	3'h4 :
		rl_a05_t5 = RG_rl_a05_d9_c1 ;
	3'h5 :
		rl_a05_t5 = RG_rl_a05_d9_c1 ;
	3'h6 :
		rl_a05_t5 = RG_rl_a05_d9_c1 ;
	3'h7 :
		rl_a05_t5 = RG_rl_a05_d9_c1 ;
	default :
		rl_a05_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a06_d9_c1 or RG_rl_a06_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a06_t5 = RG_rl_a06_d9_c0 ;
	3'h1 :
		rl_a06_t5 = RG_rl_a06_d9_c1 ;
	3'h2 :
		rl_a06_t5 = RG_rl_a06_d9_c1 ;
	3'h3 :
		rl_a06_t5 = RG_rl_a06_d9_c1 ;
	3'h4 :
		rl_a06_t5 = RG_rl_a06_d9_c1 ;
	3'h5 :
		rl_a06_t5 = RG_rl_a06_d9_c1 ;
	3'h6 :
		rl_a06_t5 = RG_rl_a06_d9_c1 ;
	3'h7 :
		rl_a06_t5 = RG_rl_a06_d9_c1 ;
	default :
		rl_a06_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a07_d9_c1 or RG_rl_a07_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a07_t5 = RG_rl_a07_d9_c0 ;
	3'h1 :
		rl_a07_t5 = RG_rl_a07_d9_c1 ;
	3'h2 :
		rl_a07_t5 = RG_rl_a07_d9_c1 ;
	3'h3 :
		rl_a07_t5 = RG_rl_a07_d9_c1 ;
	3'h4 :
		rl_a07_t5 = RG_rl_a07_d9_c1 ;
	3'h5 :
		rl_a07_t5 = RG_rl_a07_d9_c1 ;
	3'h6 :
		rl_a07_t5 = RG_rl_a07_d9_c1 ;
	3'h7 :
		rl_a07_t5 = RG_rl_a07_d9_c1 ;
	default :
		rl_a07_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a08_d9_c1 or RG_rl_a08_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a08_t5 = RG_rl_a08_d9_c0 ;
	3'h1 :
		rl_a08_t5 = RG_rl_a08_d9_c1 ;
	3'h2 :
		rl_a08_t5 = RG_rl_a08_d9_c1 ;
	3'h3 :
		rl_a08_t5 = RG_rl_a08_d9_c1 ;
	3'h4 :
		rl_a08_t5 = RG_rl_a08_d9_c1 ;
	3'h5 :
		rl_a08_t5 = RG_rl_a08_d9_c1 ;
	3'h6 :
		rl_a08_t5 = RG_rl_a08_d9_c1 ;
	3'h7 :
		rl_a08_t5 = RG_rl_a08_d9_c1 ;
	default :
		rl_a08_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a09_d9_c1 or RG_rl_a09_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a09_t5 = RG_rl_a09_d9_c0 ;
	3'h1 :
		rl_a09_t5 = RG_rl_a09_d9_c1 ;
	3'h2 :
		rl_a09_t5 = RG_rl_a09_d9_c1 ;
	3'h3 :
		rl_a09_t5 = RG_rl_a09_d9_c1 ;
	3'h4 :
		rl_a09_t5 = RG_rl_a09_d9_c1 ;
	3'h5 :
		rl_a09_t5 = RG_rl_a09_d9_c1 ;
	3'h6 :
		rl_a09_t5 = RG_rl_a09_d9_c1 ;
	3'h7 :
		rl_a09_t5 = RG_rl_a09_d9_c1 ;
	default :
		rl_a09_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a10_d9_c1 or RG_rl_a10_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a10_t5 = RG_rl_a10_d9_c0 ;
	3'h1 :
		rl_a10_t5 = RG_rl_a10_d9_c1 ;
	3'h2 :
		rl_a10_t5 = RG_rl_a10_d9_c1 ;
	3'h3 :
		rl_a10_t5 = RG_rl_a10_d9_c1 ;
	3'h4 :
		rl_a10_t5 = RG_rl_a10_d9_c1 ;
	3'h5 :
		rl_a10_t5 = RG_rl_a10_d9_c1 ;
	3'h6 :
		rl_a10_t5 = RG_rl_a10_d9_c1 ;
	3'h7 :
		rl_a10_t5 = RG_rl_a10_d9_c1 ;
	default :
		rl_a10_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a11_d9_c1 or RG_rl_a11_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a11_t5 = RG_rl_a11_d9_c0 ;
	3'h1 :
		rl_a11_t5 = RG_rl_a11_d9_c1 ;
	3'h2 :
		rl_a11_t5 = RG_rl_a11_d9_c1 ;
	3'h3 :
		rl_a11_t5 = RG_rl_a11_d9_c1 ;
	3'h4 :
		rl_a11_t5 = RG_rl_a11_d9_c1 ;
	3'h5 :
		rl_a11_t5 = RG_rl_a11_d9_c1 ;
	3'h6 :
		rl_a11_t5 = RG_rl_a11_d9_c1 ;
	3'h7 :
		rl_a11_t5 = RG_rl_a11_d9_c1 ;
	default :
		rl_a11_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a12_d9_c1 or RG_rl_a12_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a12_t5 = RG_rl_a12_d9_c0 ;
	3'h1 :
		rl_a12_t5 = RG_rl_a12_d9_c1 ;
	3'h2 :
		rl_a12_t5 = RG_rl_a12_d9_c1 ;
	3'h3 :
		rl_a12_t5 = RG_rl_a12_d9_c1 ;
	3'h4 :
		rl_a12_t5 = RG_rl_a12_d9_c1 ;
	3'h5 :
		rl_a12_t5 = RG_rl_a12_d9_c1 ;
	3'h6 :
		rl_a12_t5 = RG_rl_a12_d9_c1 ;
	3'h7 :
		rl_a12_t5 = RG_rl_a12_d9_c1 ;
	default :
		rl_a12_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a13_d9_c1 or RG_rl_a13_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a13_t5 = RG_rl_a13_d9_c0 ;
	3'h1 :
		rl_a13_t5 = RG_rl_a13_d9_c1 ;
	3'h2 :
		rl_a13_t5 = RG_rl_a13_d9_c1 ;
	3'h3 :
		rl_a13_t5 = RG_rl_a13_d9_c1 ;
	3'h4 :
		rl_a13_t5 = RG_rl_a13_d9_c1 ;
	3'h5 :
		rl_a13_t5 = RG_rl_a13_d9_c1 ;
	3'h6 :
		rl_a13_t5 = RG_rl_a13_d9_c1 ;
	3'h7 :
		rl_a13_t5 = RG_rl_a13_d9_c1 ;
	default :
		rl_a13_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a14_d9_c1 or RG_rl_a14_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a14_t5 = RG_rl_a14_d9_c0 ;
	3'h1 :
		rl_a14_t5 = RG_rl_a14_d9_c1 ;
	3'h2 :
		rl_a14_t5 = RG_rl_a14_d9_c1 ;
	3'h3 :
		rl_a14_t5 = RG_rl_a14_d9_c1 ;
	3'h4 :
		rl_a14_t5 = RG_rl_a14_d9_c1 ;
	3'h5 :
		rl_a14_t5 = RG_rl_a14_d9_c1 ;
	3'h6 :
		rl_a14_t5 = RG_rl_a14_d9_c1 ;
	3'h7 :
		rl_a14_t5 = RG_rl_a14_d9_c1 ;
	default :
		rl_a14_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a15_d9_c1 or RG_rl_a15_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a15_t5 = RG_rl_a15_d9_c0 ;
	3'h1 :
		rl_a15_t5 = RG_rl_a15_d9_c1 ;
	3'h2 :
		rl_a15_t5 = RG_rl_a15_d9_c1 ;
	3'h3 :
		rl_a15_t5 = RG_rl_a15_d9_c1 ;
	3'h4 :
		rl_a15_t5 = RG_rl_a15_d9_c1 ;
	3'h5 :
		rl_a15_t5 = RG_rl_a15_d9_c1 ;
	3'h6 :
		rl_a15_t5 = RG_rl_a15_d9_c1 ;
	3'h7 :
		rl_a15_t5 = RG_rl_a15_d9_c1 ;
	default :
		rl_a15_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a16_d9_c1 or RG_rl_a16_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a16_t5 = RG_rl_a16_d9_c0 ;
	3'h1 :
		rl_a16_t5 = RG_rl_a16_d9_c1 ;
	3'h2 :
		rl_a16_t5 = RG_rl_a16_d9_c0 ;
	3'h3 :
		rl_a16_t5 = RG_rl_a16_d9_c0 ;
	3'h4 :
		rl_a16_t5 = RG_rl_a16_d9_c0 ;
	3'h5 :
		rl_a16_t5 = RG_rl_a16_d9_c0 ;
	3'h6 :
		rl_a16_t5 = RG_rl_a16_d9_c0 ;
	3'h7 :
		rl_a16_t5 = RG_rl_a16_d9_c0 ;
	default :
		rl_a16_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a17_d9_c1 or RG_rl_a17_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a17_t5 = RG_rl_a17_d9_c0 ;
	3'h1 :
		rl_a17_t5 = RG_rl_a17_d9_c1 ;
	3'h2 :
		rl_a17_t5 = RG_rl_a17_d9_c0 ;
	3'h3 :
		rl_a17_t5 = RG_rl_a17_d9_c0 ;
	3'h4 :
		rl_a17_t5 = RG_rl_a17_d9_c0 ;
	3'h5 :
		rl_a17_t5 = RG_rl_a17_d9_c0 ;
	3'h6 :
		rl_a17_t5 = RG_rl_a17_d9_c0 ;
	3'h7 :
		rl_a17_t5 = RG_rl_a17_d9_c0 ;
	default :
		rl_a17_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a18_d9_c1 or RG_rl_a18_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a18_t5 = RG_rl_a18_d9_c0 ;
	3'h1 :
		rl_a18_t5 = RG_rl_a18_d9_c1 ;
	3'h2 :
		rl_a18_t5 = RG_rl_a18_d9_c0 ;
	3'h3 :
		rl_a18_t5 = RG_rl_a18_d9_c0 ;
	3'h4 :
		rl_a18_t5 = RG_rl_a18_d9_c0 ;
	3'h5 :
		rl_a18_t5 = RG_rl_a18_d9_c0 ;
	3'h6 :
		rl_a18_t5 = RG_rl_a18_d9_c0 ;
	3'h7 :
		rl_a18_t5 = RG_rl_a18_d9_c0 ;
	default :
		rl_a18_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a19_d9_c1 or RG_rl_a19_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a19_t5 = RG_rl_a19_d9_c0 ;
	3'h1 :
		rl_a19_t5 = RG_rl_a19_d9_c1 ;
	3'h2 :
		rl_a19_t5 = RG_rl_a19_d9_c0 ;
	3'h3 :
		rl_a19_t5 = RG_rl_a19_d9_c0 ;
	3'h4 :
		rl_a19_t5 = RG_rl_a19_d9_c0 ;
	3'h5 :
		rl_a19_t5 = RG_rl_a19_d9_c0 ;
	3'h6 :
		rl_a19_t5 = RG_rl_a19_d9_c0 ;
	3'h7 :
		rl_a19_t5 = RG_rl_a19_d9_c0 ;
	default :
		rl_a19_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a20_d9_c1 or RG_rl_a20_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a20_t5 = RG_rl_a20_d9_c0 ;
	3'h1 :
		rl_a20_t5 = RG_rl_a20_d9_c1 ;
	3'h2 :
		rl_a20_t5 = RG_rl_a20_d9_c0 ;
	3'h3 :
		rl_a20_t5 = RG_rl_a20_d9_c0 ;
	3'h4 :
		rl_a20_t5 = RG_rl_a20_d9_c0 ;
	3'h5 :
		rl_a20_t5 = RG_rl_a20_d9_c0 ;
	3'h6 :
		rl_a20_t5 = RG_rl_a20_d9_c0 ;
	3'h7 :
		rl_a20_t5 = RG_rl_a20_d9_c0 ;
	default :
		rl_a20_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a21_d9_c1 or RG_rl_a21_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a21_t5 = RG_rl_a21_d9_c0 ;
	3'h1 :
		rl_a21_t5 = RG_rl_a21_d9_c1 ;
	3'h2 :
		rl_a21_t5 = RG_rl_a21_d9_c0 ;
	3'h3 :
		rl_a21_t5 = RG_rl_a21_d9_c0 ;
	3'h4 :
		rl_a21_t5 = RG_rl_a21_d9_c0 ;
	3'h5 :
		rl_a21_t5 = RG_rl_a21_d9_c0 ;
	3'h6 :
		rl_a21_t5 = RG_rl_a21_d9_c0 ;
	3'h7 :
		rl_a21_t5 = RG_rl_a21_d9_c0 ;
	default :
		rl_a21_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a22_d9_c1 or RG_rl_a22_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a22_t5 = RG_rl_a22_d9_c0 ;
	3'h1 :
		rl_a22_t5 = RG_rl_a22_d9_c1 ;
	3'h2 :
		rl_a22_t5 = RG_rl_a22_d9_c0 ;
	3'h3 :
		rl_a22_t5 = RG_rl_a22_d9_c0 ;
	3'h4 :
		rl_a22_t5 = RG_rl_a22_d9_c0 ;
	3'h5 :
		rl_a22_t5 = RG_rl_a22_d9_c0 ;
	3'h6 :
		rl_a22_t5 = RG_rl_a22_d9_c0 ;
	3'h7 :
		rl_a22_t5 = RG_rl_a22_d9_c0 ;
	default :
		rl_a22_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a23_d9_c1 or RG_rl_a23_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a23_t5 = RG_rl_a23_d9_c0 ;
	3'h1 :
		rl_a23_t5 = RG_rl_a23_d9_c1 ;
	3'h2 :
		rl_a23_t5 = RG_rl_a23_d9_c0 ;
	3'h3 :
		rl_a23_t5 = RG_rl_a23_d9_c0 ;
	3'h4 :
		rl_a23_t5 = RG_rl_a23_d9_c0 ;
	3'h5 :
		rl_a23_t5 = RG_rl_a23_d9_c0 ;
	3'h6 :
		rl_a23_t5 = RG_rl_a23_d9_c0 ;
	3'h7 :
		rl_a23_t5 = RG_rl_a23_d9_c0 ;
	default :
		rl_a23_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a24_d9_c1 or RG_rl_a24_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a24_t5 = RG_rl_a24_d9_c0 ;
	3'h1 :
		rl_a24_t5 = RG_rl_a24_d9_c1 ;
	3'h2 :
		rl_a24_t5 = RG_rl_a24_d9_c0 ;
	3'h3 :
		rl_a24_t5 = RG_rl_a24_d9_c0 ;
	3'h4 :
		rl_a24_t5 = RG_rl_a24_d9_c0 ;
	3'h5 :
		rl_a24_t5 = RG_rl_a24_d9_c0 ;
	3'h6 :
		rl_a24_t5 = RG_rl_a24_d9_c0 ;
	3'h7 :
		rl_a24_t5 = RG_rl_a24_d9_c0 ;
	default :
		rl_a24_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a25_d9_c1 or RG_rl_a25_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a25_t5 = RG_rl_a25_d9_c0 ;
	3'h1 :
		rl_a25_t5 = RG_rl_a25_d9_c1 ;
	3'h2 :
		rl_a25_t5 = RG_rl_a25_d9_c0 ;
	3'h3 :
		rl_a25_t5 = RG_rl_a25_d9_c0 ;
	3'h4 :
		rl_a25_t5 = RG_rl_a25_d9_c0 ;
	3'h5 :
		rl_a25_t5 = RG_rl_a25_d9_c0 ;
	3'h6 :
		rl_a25_t5 = RG_rl_a25_d9_c0 ;
	3'h7 :
		rl_a25_t5 = RG_rl_a25_d9_c0 ;
	default :
		rl_a25_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a26_d9_c1 or RG_rl_a26_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a26_t5 = RG_rl_a26_d9_c0 ;
	3'h1 :
		rl_a26_t5 = RG_rl_a26_d9_c1 ;
	3'h2 :
		rl_a26_t5 = RG_rl_a26_d9_c0 ;
	3'h3 :
		rl_a26_t5 = RG_rl_a26_d9_c0 ;
	3'h4 :
		rl_a26_t5 = RG_rl_a26_d9_c0 ;
	3'h5 :
		rl_a26_t5 = RG_rl_a26_d9_c0 ;
	3'h6 :
		rl_a26_t5 = RG_rl_a26_d9_c0 ;
	3'h7 :
		rl_a26_t5 = RG_rl_a26_d9_c0 ;
	default :
		rl_a26_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a27_d9_c1 or RG_rl_a27_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a27_t5 = RG_rl_a27_d9_c0 ;
	3'h1 :
		rl_a27_t5 = RG_rl_a27_d9_c1 ;
	3'h2 :
		rl_a27_t5 = RG_rl_a27_d9_c0 ;
	3'h3 :
		rl_a27_t5 = RG_rl_a27_d9_c0 ;
	3'h4 :
		rl_a27_t5 = RG_rl_a27_d9_c0 ;
	3'h5 :
		rl_a27_t5 = RG_rl_a27_d9_c0 ;
	3'h6 :
		rl_a27_t5 = RG_rl_a27_d9_c0 ;
	3'h7 :
		rl_a27_t5 = RG_rl_a27_d9_c0 ;
	default :
		rl_a27_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a28_d9_c1 or RG_rl_a28_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a28_t5 = RG_rl_a28_d9_c0 ;
	3'h1 :
		rl_a28_t5 = RG_rl_a28_d9_c1 ;
	3'h2 :
		rl_a28_t5 = RG_rl_a28_d9_c0 ;
	3'h3 :
		rl_a28_t5 = RG_rl_a28_d9_c0 ;
	3'h4 :
		rl_a28_t5 = RG_rl_a28_d9_c0 ;
	3'h5 :
		rl_a28_t5 = RG_rl_a28_d9_c0 ;
	3'h6 :
		rl_a28_t5 = RG_rl_a28_d9_c0 ;
	3'h7 :
		rl_a28_t5 = RG_rl_a28_d9_c0 ;
	default :
		rl_a28_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a29_d9_c1 or RG_rl_a29_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a29_t5 = RG_rl_a29_d9_c0 ;
	3'h1 :
		rl_a29_t5 = RG_rl_a29_d9_c1 ;
	3'h2 :
		rl_a29_t5 = RG_rl_a29_d9_c0 ;
	3'h3 :
		rl_a29_t5 = RG_rl_a29_d9_c0 ;
	3'h4 :
		rl_a29_t5 = RG_rl_a29_d9_c0 ;
	3'h5 :
		rl_a29_t5 = RG_rl_a29_d9_c0 ;
	3'h6 :
		rl_a29_t5 = RG_rl_a29_d9_c0 ;
	3'h7 :
		rl_a29_t5 = RG_rl_a29_d9_c0 ;
	default :
		rl_a29_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a30_d9_c1 or RG_rl_a30_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a30_t5 = RG_rl_a30_d9_c0 ;
	3'h1 :
		rl_a30_t5 = RG_rl_a30_d9_c1 ;
	3'h2 :
		rl_a30_t5 = RG_rl_a30_d9_c0 ;
	3'h3 :
		rl_a30_t5 = RG_rl_a30_d9_c0 ;
	3'h4 :
		rl_a30_t5 = RG_rl_a30_d9_c0 ;
	3'h5 :
		rl_a30_t5 = RG_rl_a30_d9_c0 ;
	3'h6 :
		rl_a30_t5 = RG_rl_a30_d9_c0 ;
	3'h7 :
		rl_a30_t5 = RG_rl_a30_d9_c0 ;
	default :
		rl_a30_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a31_d9_c1 or RG_rl_a31_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a31_t5 = RG_rl_a31_d9_c0 ;
	3'h1 :
		rl_a31_t5 = RG_rl_a31_d9_c1 ;
	3'h2 :
		rl_a31_t5 = RG_rl_a31_d9_c0 ;
	3'h3 :
		rl_a31_t5 = RG_rl_a31_d9_c0 ;
	3'h4 :
		rl_a31_t5 = RG_rl_a31_d9_c0 ;
	3'h5 :
		rl_a31_t5 = RG_rl_a31_d9_c0 ;
	3'h6 :
		rl_a31_t5 = RG_rl_a31_d9_c0 ;
	3'h7 :
		rl_a31_t5 = RG_rl_a31_d9_c0 ;
	default :
		rl_a31_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a32_d9_c2 or RG_rl_a32_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a32_t5 = RG_rl_a32_d9_c0 ;
	3'h1 :
		rl_a32_t5 = RG_rl_a32_d9_c0 ;
	3'h2 :
		rl_a32_t5 = RG_rl_a32_d9_c2 ;
	3'h3 :
		rl_a32_t5 = RG_rl_a32_d9_c0 ;
	3'h4 :
		rl_a32_t5 = RG_rl_a32_d9_c0 ;
	3'h5 :
		rl_a32_t5 = RG_rl_a32_d9_c0 ;
	3'h6 :
		rl_a32_t5 = RG_rl_a32_d9_c0 ;
	3'h7 :
		rl_a32_t5 = RG_rl_a32_d9_c0 ;
	default :
		rl_a32_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a33_d9_c2 or RG_rl_a33_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a33_t5 = RG_rl_a33_d9_c0 ;
	3'h1 :
		rl_a33_t5 = RG_rl_a33_d9_c0 ;
	3'h2 :
		rl_a33_t5 = RG_rl_a33_d9_c2 ;
	3'h3 :
		rl_a33_t5 = RG_rl_a33_d9_c0 ;
	3'h4 :
		rl_a33_t5 = RG_rl_a33_d9_c0 ;
	3'h5 :
		rl_a33_t5 = RG_rl_a33_d9_c0 ;
	3'h6 :
		rl_a33_t5 = RG_rl_a33_d9_c0 ;
	3'h7 :
		rl_a33_t5 = RG_rl_a33_d9_c0 ;
	default :
		rl_a33_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a34_d9_c2 or RG_rl_a34_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a34_t5 = RG_rl_a34_d9_c0 ;
	3'h1 :
		rl_a34_t5 = RG_rl_a34_d9_c0 ;
	3'h2 :
		rl_a34_t5 = RG_rl_a34_d9_c2 ;
	3'h3 :
		rl_a34_t5 = RG_rl_a34_d9_c0 ;
	3'h4 :
		rl_a34_t5 = RG_rl_a34_d9_c0 ;
	3'h5 :
		rl_a34_t5 = RG_rl_a34_d9_c0 ;
	3'h6 :
		rl_a34_t5 = RG_rl_a34_d9_c0 ;
	3'h7 :
		rl_a34_t5 = RG_rl_a34_d9_c0 ;
	default :
		rl_a34_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a35_d9_c2 or RG_rl_a35_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a35_t5 = RG_rl_a35_d9_c0 ;
	3'h1 :
		rl_a35_t5 = RG_rl_a35_d9_c0 ;
	3'h2 :
		rl_a35_t5 = RG_rl_a35_d9_c2 ;
	3'h3 :
		rl_a35_t5 = RG_rl_a35_d9_c0 ;
	3'h4 :
		rl_a35_t5 = RG_rl_a35_d9_c0 ;
	3'h5 :
		rl_a35_t5 = RG_rl_a35_d9_c0 ;
	3'h6 :
		rl_a35_t5 = RG_rl_a35_d9_c0 ;
	3'h7 :
		rl_a35_t5 = RG_rl_a35_d9_c0 ;
	default :
		rl_a35_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a36_d9_c2 or RG_rl_a36_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a36_t5 = RG_rl_a36_d9_c0 ;
	3'h1 :
		rl_a36_t5 = RG_rl_a36_d9_c0 ;
	3'h2 :
		rl_a36_t5 = RG_rl_a36_d9_c2 ;
	3'h3 :
		rl_a36_t5 = RG_rl_a36_d9_c0 ;
	3'h4 :
		rl_a36_t5 = RG_rl_a36_d9_c0 ;
	3'h5 :
		rl_a36_t5 = RG_rl_a36_d9_c0 ;
	3'h6 :
		rl_a36_t5 = RG_rl_a36_d9_c0 ;
	3'h7 :
		rl_a36_t5 = RG_rl_a36_d9_c0 ;
	default :
		rl_a36_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a37_d9_c2 or RG_rl_a37_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a37_t5 = RG_rl_a37_d9_c0 ;
	3'h1 :
		rl_a37_t5 = RG_rl_a37_d9_c0 ;
	3'h2 :
		rl_a37_t5 = RG_rl_a37_d9_c2 ;
	3'h3 :
		rl_a37_t5 = RG_rl_a37_d9_c0 ;
	3'h4 :
		rl_a37_t5 = RG_rl_a37_d9_c0 ;
	3'h5 :
		rl_a37_t5 = RG_rl_a37_d9_c0 ;
	3'h6 :
		rl_a37_t5 = RG_rl_a37_d9_c0 ;
	3'h7 :
		rl_a37_t5 = RG_rl_a37_d9_c0 ;
	default :
		rl_a37_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a38_d9_c2 or RG_rl_a38_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a38_t5 = RG_rl_a38_d9_c0 ;
	3'h1 :
		rl_a38_t5 = RG_rl_a38_d9_c0 ;
	3'h2 :
		rl_a38_t5 = RG_rl_a38_d9_c2 ;
	3'h3 :
		rl_a38_t5 = RG_rl_a38_d9_c0 ;
	3'h4 :
		rl_a38_t5 = RG_rl_a38_d9_c0 ;
	3'h5 :
		rl_a38_t5 = RG_rl_a38_d9_c0 ;
	3'h6 :
		rl_a38_t5 = RG_rl_a38_d9_c0 ;
	3'h7 :
		rl_a38_t5 = RG_rl_a38_d9_c0 ;
	default :
		rl_a38_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a39_d9_c2 or RG_rl_a39_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a39_t5 = RG_rl_a39_d9_c0 ;
	3'h1 :
		rl_a39_t5 = RG_rl_a39_d9_c0 ;
	3'h2 :
		rl_a39_t5 = RG_rl_a39_d9_c2 ;
	3'h3 :
		rl_a39_t5 = RG_rl_a39_d9_c0 ;
	3'h4 :
		rl_a39_t5 = RG_rl_a39_d9_c0 ;
	3'h5 :
		rl_a39_t5 = RG_rl_a39_d9_c0 ;
	3'h6 :
		rl_a39_t5 = RG_rl_a39_d9_c0 ;
	3'h7 :
		rl_a39_t5 = RG_rl_a39_d9_c0 ;
	default :
		rl_a39_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a40_d9_c2 or RG_rl_a40_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a40_t5 = RG_rl_a40_d9_c0 ;
	3'h1 :
		rl_a40_t5 = RG_rl_a40_d9_c0 ;
	3'h2 :
		rl_a40_t5 = RG_rl_a40_d9_c2 ;
	3'h3 :
		rl_a40_t5 = RG_rl_a40_d9_c0 ;
	3'h4 :
		rl_a40_t5 = RG_rl_a40_d9_c0 ;
	3'h5 :
		rl_a40_t5 = RG_rl_a40_d9_c0 ;
	3'h6 :
		rl_a40_t5 = RG_rl_a40_d9_c0 ;
	3'h7 :
		rl_a40_t5 = RG_rl_a40_d9_c0 ;
	default :
		rl_a40_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a41_d9_c2 or RG_rl_a41_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a41_t5 = RG_rl_a41_d9_c0 ;
	3'h1 :
		rl_a41_t5 = RG_rl_a41_d9_c0 ;
	3'h2 :
		rl_a41_t5 = RG_rl_a41_d9_c2 ;
	3'h3 :
		rl_a41_t5 = RG_rl_a41_d9_c0 ;
	3'h4 :
		rl_a41_t5 = RG_rl_a41_d9_c0 ;
	3'h5 :
		rl_a41_t5 = RG_rl_a41_d9_c0 ;
	3'h6 :
		rl_a41_t5 = RG_rl_a41_d9_c0 ;
	3'h7 :
		rl_a41_t5 = RG_rl_a41_d9_c0 ;
	default :
		rl_a41_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a42_d9_c2 or RG_rl_a42_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a42_t5 = RG_rl_a42_d9_c0 ;
	3'h1 :
		rl_a42_t5 = RG_rl_a42_d9_c0 ;
	3'h2 :
		rl_a42_t5 = RG_rl_a42_d9_c2 ;
	3'h3 :
		rl_a42_t5 = RG_rl_a42_d9_c0 ;
	3'h4 :
		rl_a42_t5 = RG_rl_a42_d9_c0 ;
	3'h5 :
		rl_a42_t5 = RG_rl_a42_d9_c0 ;
	3'h6 :
		rl_a42_t5 = RG_rl_a42_d9_c0 ;
	3'h7 :
		rl_a42_t5 = RG_rl_a42_d9_c0 ;
	default :
		rl_a42_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a43_d9_c2 or RG_rl_a43_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a43_t5 = RG_rl_a43_d9_c0 ;
	3'h1 :
		rl_a43_t5 = RG_rl_a43_d9_c0 ;
	3'h2 :
		rl_a43_t5 = RG_rl_a43_d9_c2 ;
	3'h3 :
		rl_a43_t5 = RG_rl_a43_d9_c0 ;
	3'h4 :
		rl_a43_t5 = RG_rl_a43_d9_c0 ;
	3'h5 :
		rl_a43_t5 = RG_rl_a43_d9_c0 ;
	3'h6 :
		rl_a43_t5 = RG_rl_a43_d9_c0 ;
	3'h7 :
		rl_a43_t5 = RG_rl_a43_d9_c0 ;
	default :
		rl_a43_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a44_d9_c2 or RG_rl_a44_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a44_t5 = RG_rl_a44_d9_c0 ;
	3'h1 :
		rl_a44_t5 = RG_rl_a44_d9_c0 ;
	3'h2 :
		rl_a44_t5 = RG_rl_a44_d9_c2 ;
	3'h3 :
		rl_a44_t5 = RG_rl_a44_d9_c0 ;
	3'h4 :
		rl_a44_t5 = RG_rl_a44_d9_c0 ;
	3'h5 :
		rl_a44_t5 = RG_rl_a44_d9_c0 ;
	3'h6 :
		rl_a44_t5 = RG_rl_a44_d9_c0 ;
	3'h7 :
		rl_a44_t5 = RG_rl_a44_d9_c0 ;
	default :
		rl_a44_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a45_d9_c2 or RG_rl_a45_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a45_t5 = RG_rl_a45_d9_c0 ;
	3'h1 :
		rl_a45_t5 = RG_rl_a45_d9_c0 ;
	3'h2 :
		rl_a45_t5 = RG_rl_a45_d9_c2 ;
	3'h3 :
		rl_a45_t5 = RG_rl_a45_d9_c0 ;
	3'h4 :
		rl_a45_t5 = RG_rl_a45_d9_c0 ;
	3'h5 :
		rl_a45_t5 = RG_rl_a45_d9_c0 ;
	3'h6 :
		rl_a45_t5 = RG_rl_a45_d9_c0 ;
	3'h7 :
		rl_a45_t5 = RG_rl_a45_d9_c0 ;
	default :
		rl_a45_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a46_d9_c2 or RG_rl_a46_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a46_t5 = RG_rl_a46_d9_c0 ;
	3'h1 :
		rl_a46_t5 = RG_rl_a46_d9_c0 ;
	3'h2 :
		rl_a46_t5 = RG_rl_a46_d9_c2 ;
	3'h3 :
		rl_a46_t5 = RG_rl_a46_d9_c0 ;
	3'h4 :
		rl_a46_t5 = RG_rl_a46_d9_c0 ;
	3'h5 :
		rl_a46_t5 = RG_rl_a46_d9_c0 ;
	3'h6 :
		rl_a46_t5 = RG_rl_a46_d9_c0 ;
	3'h7 :
		rl_a46_t5 = RG_rl_a46_d9_c0 ;
	default :
		rl_a46_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a47_d9_c2 or RG_rl_a47_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a47_t5 = RG_rl_a47_d9_c0 ;
	3'h1 :
		rl_a47_t5 = RG_rl_a47_d9_c0 ;
	3'h2 :
		rl_a47_t5 = RG_rl_a47_d9_c2 ;
	3'h3 :
		rl_a47_t5 = RG_rl_a47_d9_c0 ;
	3'h4 :
		rl_a47_t5 = RG_rl_a47_d9_c0 ;
	3'h5 :
		rl_a47_t5 = RG_rl_a47_d9_c0 ;
	3'h6 :
		rl_a47_t5 = RG_rl_a47_d9_c0 ;
	3'h7 :
		rl_a47_t5 = RG_rl_a47_d9_c0 ;
	default :
		rl_a47_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a48_d9_c3 or RG_rl_a48_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a48_t5 = RG_rl_a48_d9_c0 ;
	3'h1 :
		rl_a48_t5 = RG_rl_a48_d9_c0 ;
	3'h2 :
		rl_a48_t5 = RG_rl_a48_d9_c0 ;
	3'h3 :
		rl_a48_t5 = RG_rl_a48_d9_c3 ;
	3'h4 :
		rl_a48_t5 = RG_rl_a48_d9_c0 ;
	3'h5 :
		rl_a48_t5 = RG_rl_a48_d9_c0 ;
	3'h6 :
		rl_a48_t5 = RG_rl_a48_d9_c0 ;
	3'h7 :
		rl_a48_t5 = RG_rl_a48_d9_c0 ;
	default :
		rl_a48_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a49_d9_c3 or RG_rl_a49_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a49_t5 = RG_rl_a49_d9_c0 ;
	3'h1 :
		rl_a49_t5 = RG_rl_a49_d9_c0 ;
	3'h2 :
		rl_a49_t5 = RG_rl_a49_d9_c0 ;
	3'h3 :
		rl_a49_t5 = RG_rl_a49_d9_c3 ;
	3'h4 :
		rl_a49_t5 = RG_rl_a49_d9_c0 ;
	3'h5 :
		rl_a49_t5 = RG_rl_a49_d9_c0 ;
	3'h6 :
		rl_a49_t5 = RG_rl_a49_d9_c0 ;
	3'h7 :
		rl_a49_t5 = RG_rl_a49_d9_c0 ;
	default :
		rl_a49_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a50_d9_c3 or RG_rl_a50_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a50_t5 = RG_rl_a50_d9_c0 ;
	3'h1 :
		rl_a50_t5 = RG_rl_a50_d9_c0 ;
	3'h2 :
		rl_a50_t5 = RG_rl_a50_d9_c0 ;
	3'h3 :
		rl_a50_t5 = RG_rl_a50_d9_c3 ;
	3'h4 :
		rl_a50_t5 = RG_rl_a50_d9_c0 ;
	3'h5 :
		rl_a50_t5 = RG_rl_a50_d9_c0 ;
	3'h6 :
		rl_a50_t5 = RG_rl_a50_d9_c0 ;
	3'h7 :
		rl_a50_t5 = RG_rl_a50_d9_c0 ;
	default :
		rl_a50_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a51_d9_c3 or RG_rl_a51_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a51_t5 = RG_rl_a51_d9_c0 ;
	3'h1 :
		rl_a51_t5 = RG_rl_a51_d9_c0 ;
	3'h2 :
		rl_a51_t5 = RG_rl_a51_d9_c0 ;
	3'h3 :
		rl_a51_t5 = RG_rl_a51_d9_c3 ;
	3'h4 :
		rl_a51_t5 = RG_rl_a51_d9_c0 ;
	3'h5 :
		rl_a51_t5 = RG_rl_a51_d9_c0 ;
	3'h6 :
		rl_a51_t5 = RG_rl_a51_d9_c0 ;
	3'h7 :
		rl_a51_t5 = RG_rl_a51_d9_c0 ;
	default :
		rl_a51_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a52_d9_c3 or RG_rl_a52_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a52_t5 = RG_rl_a52_d9_c0 ;
	3'h1 :
		rl_a52_t5 = RG_rl_a52_d9_c0 ;
	3'h2 :
		rl_a52_t5 = RG_rl_a52_d9_c0 ;
	3'h3 :
		rl_a52_t5 = RG_rl_a52_d9_c3 ;
	3'h4 :
		rl_a52_t5 = RG_rl_a52_d9_c0 ;
	3'h5 :
		rl_a52_t5 = RG_rl_a52_d9_c0 ;
	3'h6 :
		rl_a52_t5 = RG_rl_a52_d9_c0 ;
	3'h7 :
		rl_a52_t5 = RG_rl_a52_d9_c0 ;
	default :
		rl_a52_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a53_d9_c3 or RG_rl_a53_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a53_t5 = RG_rl_a53_d9_c0 ;
	3'h1 :
		rl_a53_t5 = RG_rl_a53_d9_c0 ;
	3'h2 :
		rl_a53_t5 = RG_rl_a53_d9_c0 ;
	3'h3 :
		rl_a53_t5 = RG_rl_a53_d9_c3 ;
	3'h4 :
		rl_a53_t5 = RG_rl_a53_d9_c0 ;
	3'h5 :
		rl_a53_t5 = RG_rl_a53_d9_c0 ;
	3'h6 :
		rl_a53_t5 = RG_rl_a53_d9_c0 ;
	3'h7 :
		rl_a53_t5 = RG_rl_a53_d9_c0 ;
	default :
		rl_a53_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a54_d9_c3 or RG_rl_a54_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a54_t5 = RG_rl_a54_d9_c0 ;
	3'h1 :
		rl_a54_t5 = RG_rl_a54_d9_c0 ;
	3'h2 :
		rl_a54_t5 = RG_rl_a54_d9_c0 ;
	3'h3 :
		rl_a54_t5 = RG_rl_a54_d9_c3 ;
	3'h4 :
		rl_a54_t5 = RG_rl_a54_d9_c0 ;
	3'h5 :
		rl_a54_t5 = RG_rl_a54_d9_c0 ;
	3'h6 :
		rl_a54_t5 = RG_rl_a54_d9_c0 ;
	3'h7 :
		rl_a54_t5 = RG_rl_a54_d9_c0 ;
	default :
		rl_a54_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a55_d9_c3 or RG_rl_a55_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a55_t5 = RG_rl_a55_d9_c0 ;
	3'h1 :
		rl_a55_t5 = RG_rl_a55_d9_c0 ;
	3'h2 :
		rl_a55_t5 = RG_rl_a55_d9_c0 ;
	3'h3 :
		rl_a55_t5 = RG_rl_a55_d9_c3 ;
	3'h4 :
		rl_a55_t5 = RG_rl_a55_d9_c0 ;
	3'h5 :
		rl_a55_t5 = RG_rl_a55_d9_c0 ;
	3'h6 :
		rl_a55_t5 = RG_rl_a55_d9_c0 ;
	3'h7 :
		rl_a55_t5 = RG_rl_a55_d9_c0 ;
	default :
		rl_a55_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a56_d9_c3 or RG_rl_a56_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a56_t5 = RG_rl_a56_d9_c0 ;
	3'h1 :
		rl_a56_t5 = RG_rl_a56_d9_c0 ;
	3'h2 :
		rl_a56_t5 = RG_rl_a56_d9_c0 ;
	3'h3 :
		rl_a56_t5 = RG_rl_a56_d9_c3 ;
	3'h4 :
		rl_a56_t5 = RG_rl_a56_d9_c0 ;
	3'h5 :
		rl_a56_t5 = RG_rl_a56_d9_c0 ;
	3'h6 :
		rl_a56_t5 = RG_rl_a56_d9_c0 ;
	3'h7 :
		rl_a56_t5 = RG_rl_a56_d9_c0 ;
	default :
		rl_a56_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a57_d9_c3 or RG_rl_a57_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a57_t5 = RG_rl_a57_d9_c0 ;
	3'h1 :
		rl_a57_t5 = RG_rl_a57_d9_c0 ;
	3'h2 :
		rl_a57_t5 = RG_rl_a57_d9_c0 ;
	3'h3 :
		rl_a57_t5 = RG_rl_a57_d9_c3 ;
	3'h4 :
		rl_a57_t5 = RG_rl_a57_d9_c0 ;
	3'h5 :
		rl_a57_t5 = RG_rl_a57_d9_c0 ;
	3'h6 :
		rl_a57_t5 = RG_rl_a57_d9_c0 ;
	3'h7 :
		rl_a57_t5 = RG_rl_a57_d9_c0 ;
	default :
		rl_a57_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a58_d9_c3 or RG_rl_a58_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a58_t5 = RG_rl_a58_d9_c0 ;
	3'h1 :
		rl_a58_t5 = RG_rl_a58_d9_c0 ;
	3'h2 :
		rl_a58_t5 = RG_rl_a58_d9_c0 ;
	3'h3 :
		rl_a58_t5 = RG_rl_a58_d9_c3 ;
	3'h4 :
		rl_a58_t5 = RG_rl_a58_d9_c0 ;
	3'h5 :
		rl_a58_t5 = RG_rl_a58_d9_c0 ;
	3'h6 :
		rl_a58_t5 = RG_rl_a58_d9_c0 ;
	3'h7 :
		rl_a58_t5 = RG_rl_a58_d9_c0 ;
	default :
		rl_a58_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a59_d9_c3 or RG_rl_a59_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a59_t5 = RG_rl_a59_d9_c0 ;
	3'h1 :
		rl_a59_t5 = RG_rl_a59_d9_c0 ;
	3'h2 :
		rl_a59_t5 = RG_rl_a59_d9_c0 ;
	3'h3 :
		rl_a59_t5 = RG_rl_a59_d9_c3 ;
	3'h4 :
		rl_a59_t5 = RG_rl_a59_d9_c0 ;
	3'h5 :
		rl_a59_t5 = RG_rl_a59_d9_c0 ;
	3'h6 :
		rl_a59_t5 = RG_rl_a59_d9_c0 ;
	3'h7 :
		rl_a59_t5 = RG_rl_a59_d9_c0 ;
	default :
		rl_a59_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a60_d9_c3 or RG_rl_a60_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a60_t5 = RG_rl_a60_d9_c0 ;
	3'h1 :
		rl_a60_t5 = RG_rl_a60_d9_c0 ;
	3'h2 :
		rl_a60_t5 = RG_rl_a60_d9_c0 ;
	3'h3 :
		rl_a60_t5 = RG_rl_a60_d9_c3 ;
	3'h4 :
		rl_a60_t5 = RG_rl_a60_d9_c0 ;
	3'h5 :
		rl_a60_t5 = RG_rl_a60_d9_c0 ;
	3'h6 :
		rl_a60_t5 = RG_rl_a60_d9_c0 ;
	3'h7 :
		rl_a60_t5 = RG_rl_a60_d9_c0 ;
	default :
		rl_a60_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a61_d9_c3 or RG_rl_a61_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a61_t5 = RG_rl_a61_d9_c0 ;
	3'h1 :
		rl_a61_t5 = RG_rl_a61_d9_c0 ;
	3'h2 :
		rl_a61_t5 = RG_rl_a61_d9_c0 ;
	3'h3 :
		rl_a61_t5 = RG_rl_a61_d9_c3 ;
	3'h4 :
		rl_a61_t5 = RG_rl_a61_d9_c0 ;
	3'h5 :
		rl_a61_t5 = RG_rl_a61_d9_c0 ;
	3'h6 :
		rl_a61_t5 = RG_rl_a61_d9_c0 ;
	3'h7 :
		rl_a61_t5 = RG_rl_a61_d9_c0 ;
	default :
		rl_a61_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a62_d9_c3 or RG_rl_a62_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a62_t5 = RG_rl_a62_d9_c0 ;
	3'h1 :
		rl_a62_t5 = RG_rl_a62_d9_c0 ;
	3'h2 :
		rl_a62_t5 = RG_rl_a62_d9_c0 ;
	3'h3 :
		rl_a62_t5 = RG_rl_a62_d9_c3 ;
	3'h4 :
		rl_a62_t5 = RG_rl_a62_d9_c0 ;
	3'h5 :
		rl_a62_t5 = RG_rl_a62_d9_c0 ;
	3'h6 :
		rl_a62_t5 = RG_rl_a62_d9_c0 ;
	3'h7 :
		rl_a62_t5 = RG_rl_a62_d9_c0 ;
	default :
		rl_a62_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a63_d9_c3 or RG_rl_a63_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a63_t5 = RG_rl_a63_d9_c0 ;
	3'h1 :
		rl_a63_t5 = RG_rl_a63_d9_c0 ;
	3'h2 :
		rl_a63_t5 = RG_rl_a63_d9_c0 ;
	3'h3 :
		rl_a63_t5 = RG_rl_a63_d9_c3 ;
	3'h4 :
		rl_a63_t5 = RG_rl_a63_d9_c0 ;
	3'h5 :
		rl_a63_t5 = RG_rl_a63_d9_c0 ;
	3'h6 :
		rl_a63_t5 = RG_rl_a63_d9_c0 ;
	3'h7 :
		rl_a63_t5 = RG_rl_a63_d9_c0 ;
	default :
		rl_a63_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a64_d9_c4 or RG_rl_a64_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a64_t5 = RG_rl_a64_d9_c0 ;
	3'h1 :
		rl_a64_t5 = RG_rl_a64_d9_c0 ;
	3'h2 :
		rl_a64_t5 = RG_rl_a64_d9_c0 ;
	3'h3 :
		rl_a64_t5 = RG_rl_a64_d9_c0 ;
	3'h4 :
		rl_a64_t5 = RG_rl_a64_d9_c4 ;
	3'h5 :
		rl_a64_t5 = RG_rl_a64_d9_c0 ;
	3'h6 :
		rl_a64_t5 = RG_rl_a64_d9_c0 ;
	3'h7 :
		rl_a64_t5 = RG_rl_a64_d9_c0 ;
	default :
		rl_a64_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a65_d9_c4 or RG_rl_a65_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a65_t5 = RG_rl_a65_d9_c0 ;
	3'h1 :
		rl_a65_t5 = RG_rl_a65_d9_c0 ;
	3'h2 :
		rl_a65_t5 = RG_rl_a65_d9_c0 ;
	3'h3 :
		rl_a65_t5 = RG_rl_a65_d9_c0 ;
	3'h4 :
		rl_a65_t5 = RG_rl_a65_d9_c4 ;
	3'h5 :
		rl_a65_t5 = RG_rl_a65_d9_c0 ;
	3'h6 :
		rl_a65_t5 = RG_rl_a65_d9_c0 ;
	3'h7 :
		rl_a65_t5 = RG_rl_a65_d9_c0 ;
	default :
		rl_a65_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a66_d9_c4 or RG_rl_a66_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a66_t5 = RG_rl_a66_d9_c0 ;
	3'h1 :
		rl_a66_t5 = RG_rl_a66_d9_c0 ;
	3'h2 :
		rl_a66_t5 = RG_rl_a66_d9_c0 ;
	3'h3 :
		rl_a66_t5 = RG_rl_a66_d9_c0 ;
	3'h4 :
		rl_a66_t5 = RG_rl_a66_d9_c4 ;
	3'h5 :
		rl_a66_t5 = RG_rl_a66_d9_c0 ;
	3'h6 :
		rl_a66_t5 = RG_rl_a66_d9_c0 ;
	3'h7 :
		rl_a66_t5 = RG_rl_a66_d9_c0 ;
	default :
		rl_a66_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a67_d9_c4 or RG_rl_a67_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a67_t5 = RG_rl_a67_d9_c0 ;
	3'h1 :
		rl_a67_t5 = RG_rl_a67_d9_c0 ;
	3'h2 :
		rl_a67_t5 = RG_rl_a67_d9_c0 ;
	3'h3 :
		rl_a67_t5 = RG_rl_a67_d9_c0 ;
	3'h4 :
		rl_a67_t5 = RG_rl_a67_d9_c4 ;
	3'h5 :
		rl_a67_t5 = RG_rl_a67_d9_c0 ;
	3'h6 :
		rl_a67_t5 = RG_rl_a67_d9_c0 ;
	3'h7 :
		rl_a67_t5 = RG_rl_a67_d9_c0 ;
	default :
		rl_a67_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a68_d9_c4 or RG_rl_a68_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a68_t5 = RG_rl_a68_d9_c0 ;
	3'h1 :
		rl_a68_t5 = RG_rl_a68_d9_c0 ;
	3'h2 :
		rl_a68_t5 = RG_rl_a68_d9_c0 ;
	3'h3 :
		rl_a68_t5 = RG_rl_a68_d9_c0 ;
	3'h4 :
		rl_a68_t5 = RG_rl_a68_d9_c4 ;
	3'h5 :
		rl_a68_t5 = RG_rl_a68_d9_c0 ;
	3'h6 :
		rl_a68_t5 = RG_rl_a68_d9_c0 ;
	3'h7 :
		rl_a68_t5 = RG_rl_a68_d9_c0 ;
	default :
		rl_a68_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a69_d9_c4 or RG_rl_a69_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a69_t5 = RG_rl_a69_d9_c0 ;
	3'h1 :
		rl_a69_t5 = RG_rl_a69_d9_c0 ;
	3'h2 :
		rl_a69_t5 = RG_rl_a69_d9_c0 ;
	3'h3 :
		rl_a69_t5 = RG_rl_a69_d9_c0 ;
	3'h4 :
		rl_a69_t5 = RG_rl_a69_d9_c4 ;
	3'h5 :
		rl_a69_t5 = RG_rl_a69_d9_c0 ;
	3'h6 :
		rl_a69_t5 = RG_rl_a69_d9_c0 ;
	3'h7 :
		rl_a69_t5 = RG_rl_a69_d9_c0 ;
	default :
		rl_a69_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a70_d9_c4 or RG_rl_a70_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a70_t5 = RG_rl_a70_d9_c0 ;
	3'h1 :
		rl_a70_t5 = RG_rl_a70_d9_c0 ;
	3'h2 :
		rl_a70_t5 = RG_rl_a70_d9_c0 ;
	3'h3 :
		rl_a70_t5 = RG_rl_a70_d9_c0 ;
	3'h4 :
		rl_a70_t5 = RG_rl_a70_d9_c4 ;
	3'h5 :
		rl_a70_t5 = RG_rl_a70_d9_c0 ;
	3'h6 :
		rl_a70_t5 = RG_rl_a70_d9_c0 ;
	3'h7 :
		rl_a70_t5 = RG_rl_a70_d9_c0 ;
	default :
		rl_a70_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a71_d9_c4 or RG_rl_a71_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a71_t5 = RG_rl_a71_d9_c0 ;
	3'h1 :
		rl_a71_t5 = RG_rl_a71_d9_c0 ;
	3'h2 :
		rl_a71_t5 = RG_rl_a71_d9_c0 ;
	3'h3 :
		rl_a71_t5 = RG_rl_a71_d9_c0 ;
	3'h4 :
		rl_a71_t5 = RG_rl_a71_d9_c4 ;
	3'h5 :
		rl_a71_t5 = RG_rl_a71_d9_c0 ;
	3'h6 :
		rl_a71_t5 = RG_rl_a71_d9_c0 ;
	3'h7 :
		rl_a71_t5 = RG_rl_a71_d9_c0 ;
	default :
		rl_a71_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a72_d9_c4 or RG_rl_a72_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a72_t5 = RG_rl_a72_d9_c0 ;
	3'h1 :
		rl_a72_t5 = RG_rl_a72_d9_c0 ;
	3'h2 :
		rl_a72_t5 = RG_rl_a72_d9_c0 ;
	3'h3 :
		rl_a72_t5 = RG_rl_a72_d9_c0 ;
	3'h4 :
		rl_a72_t5 = RG_rl_a72_d9_c4 ;
	3'h5 :
		rl_a72_t5 = RG_rl_a72_d9_c0 ;
	3'h6 :
		rl_a72_t5 = RG_rl_a72_d9_c0 ;
	3'h7 :
		rl_a72_t5 = RG_rl_a72_d9_c0 ;
	default :
		rl_a72_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a73_d9_c4 or RG_rl_a73_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a73_t5 = RG_rl_a73_d9_c0 ;
	3'h1 :
		rl_a73_t5 = RG_rl_a73_d9_c0 ;
	3'h2 :
		rl_a73_t5 = RG_rl_a73_d9_c0 ;
	3'h3 :
		rl_a73_t5 = RG_rl_a73_d9_c0 ;
	3'h4 :
		rl_a73_t5 = RG_rl_a73_d9_c4 ;
	3'h5 :
		rl_a73_t5 = RG_rl_a73_d9_c0 ;
	3'h6 :
		rl_a73_t5 = RG_rl_a73_d9_c0 ;
	3'h7 :
		rl_a73_t5 = RG_rl_a73_d9_c0 ;
	default :
		rl_a73_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a74_d9_c4 or RG_rl_a74_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a74_t5 = RG_rl_a74_d9_c0 ;
	3'h1 :
		rl_a74_t5 = RG_rl_a74_d9_c0 ;
	3'h2 :
		rl_a74_t5 = RG_rl_a74_d9_c0 ;
	3'h3 :
		rl_a74_t5 = RG_rl_a74_d9_c0 ;
	3'h4 :
		rl_a74_t5 = RG_rl_a74_d9_c4 ;
	3'h5 :
		rl_a74_t5 = RG_rl_a74_d9_c0 ;
	3'h6 :
		rl_a74_t5 = RG_rl_a74_d9_c0 ;
	3'h7 :
		rl_a74_t5 = RG_rl_a74_d9_c0 ;
	default :
		rl_a74_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a75_d9_c4 or RG_rl_a75_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a75_t5 = RG_rl_a75_d9_c0 ;
	3'h1 :
		rl_a75_t5 = RG_rl_a75_d9_c0 ;
	3'h2 :
		rl_a75_t5 = RG_rl_a75_d9_c0 ;
	3'h3 :
		rl_a75_t5 = RG_rl_a75_d9_c0 ;
	3'h4 :
		rl_a75_t5 = RG_rl_a75_d9_c4 ;
	3'h5 :
		rl_a75_t5 = RG_rl_a75_d9_c0 ;
	3'h6 :
		rl_a75_t5 = RG_rl_a75_d9_c0 ;
	3'h7 :
		rl_a75_t5 = RG_rl_a75_d9_c0 ;
	default :
		rl_a75_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a76_d9_c4 or RG_rl_a76_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a76_t5 = RG_rl_a76_d9_c0 ;
	3'h1 :
		rl_a76_t5 = RG_rl_a76_d9_c0 ;
	3'h2 :
		rl_a76_t5 = RG_rl_a76_d9_c0 ;
	3'h3 :
		rl_a76_t5 = RG_rl_a76_d9_c0 ;
	3'h4 :
		rl_a76_t5 = RG_rl_a76_d9_c4 ;
	3'h5 :
		rl_a76_t5 = RG_rl_a76_d9_c0 ;
	3'h6 :
		rl_a76_t5 = RG_rl_a76_d9_c0 ;
	3'h7 :
		rl_a76_t5 = RG_rl_a76_d9_c0 ;
	default :
		rl_a76_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a77_d9_c4 or RG_rl_a77_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a77_t5 = RG_rl_a77_d9_c0 ;
	3'h1 :
		rl_a77_t5 = RG_rl_a77_d9_c0 ;
	3'h2 :
		rl_a77_t5 = RG_rl_a77_d9_c0 ;
	3'h3 :
		rl_a77_t5 = RG_rl_a77_d9_c0 ;
	3'h4 :
		rl_a77_t5 = RG_rl_a77_d9_c4 ;
	3'h5 :
		rl_a77_t5 = RG_rl_a77_d9_c0 ;
	3'h6 :
		rl_a77_t5 = RG_rl_a77_d9_c0 ;
	3'h7 :
		rl_a77_t5 = RG_rl_a77_d9_c0 ;
	default :
		rl_a77_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a78_d9_c4 or RG_rl_a78_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a78_t5 = RG_rl_a78_d9_c0 ;
	3'h1 :
		rl_a78_t5 = RG_rl_a78_d9_c0 ;
	3'h2 :
		rl_a78_t5 = RG_rl_a78_d9_c0 ;
	3'h3 :
		rl_a78_t5 = RG_rl_a78_d9_c0 ;
	3'h4 :
		rl_a78_t5 = RG_rl_a78_d9_c4 ;
	3'h5 :
		rl_a78_t5 = RG_rl_a78_d9_c0 ;
	3'h6 :
		rl_a78_t5 = RG_rl_a78_d9_c0 ;
	3'h7 :
		rl_a78_t5 = RG_rl_a78_d9_c0 ;
	default :
		rl_a78_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a79_d9_c4 or RG_rl_a79_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a79_t5 = RG_rl_a79_d9_c0 ;
	3'h1 :
		rl_a79_t5 = RG_rl_a79_d9_c0 ;
	3'h2 :
		rl_a79_t5 = RG_rl_a79_d9_c0 ;
	3'h3 :
		rl_a79_t5 = RG_rl_a79_d9_c0 ;
	3'h4 :
		rl_a79_t5 = RG_rl_a79_d9_c4 ;
	3'h5 :
		rl_a79_t5 = RG_rl_a79_d9_c0 ;
	3'h6 :
		rl_a79_t5 = RG_rl_a79_d9_c0 ;
	3'h7 :
		rl_a79_t5 = RG_rl_a79_d9_c0 ;
	default :
		rl_a79_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a80_d9_c5 or RG_rl_a80_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a80_t5 = RG_rl_a80_d9_c0 ;
	3'h1 :
		rl_a80_t5 = RG_rl_a80_d9_c0 ;
	3'h2 :
		rl_a80_t5 = RG_rl_a80_d9_c0 ;
	3'h3 :
		rl_a80_t5 = RG_rl_a80_d9_c0 ;
	3'h4 :
		rl_a80_t5 = RG_rl_a80_d9_c0 ;
	3'h5 :
		rl_a80_t5 = RG_rl_a80_d9_c5 ;
	3'h6 :
		rl_a80_t5 = RG_rl_a80_d9_c0 ;
	3'h7 :
		rl_a80_t5 = RG_rl_a80_d9_c0 ;
	default :
		rl_a80_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a81_d9_c5 or RG_rl_a81_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a81_t5 = RG_rl_a81_d9_c0 ;
	3'h1 :
		rl_a81_t5 = RG_rl_a81_d9_c0 ;
	3'h2 :
		rl_a81_t5 = RG_rl_a81_d9_c0 ;
	3'h3 :
		rl_a81_t5 = RG_rl_a81_d9_c0 ;
	3'h4 :
		rl_a81_t5 = RG_rl_a81_d9_c0 ;
	3'h5 :
		rl_a81_t5 = RG_rl_a81_d9_c5 ;
	3'h6 :
		rl_a81_t5 = RG_rl_a81_d9_c0 ;
	3'h7 :
		rl_a81_t5 = RG_rl_a81_d9_c0 ;
	default :
		rl_a81_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a82_d9_c5 or RG_rl_a82_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a82_t5 = RG_rl_a82_d9_c0 ;
	3'h1 :
		rl_a82_t5 = RG_rl_a82_d9_c0 ;
	3'h2 :
		rl_a82_t5 = RG_rl_a82_d9_c0 ;
	3'h3 :
		rl_a82_t5 = RG_rl_a82_d9_c0 ;
	3'h4 :
		rl_a82_t5 = RG_rl_a82_d9_c0 ;
	3'h5 :
		rl_a82_t5 = RG_rl_a82_d9_c5 ;
	3'h6 :
		rl_a82_t5 = RG_rl_a82_d9_c0 ;
	3'h7 :
		rl_a82_t5 = RG_rl_a82_d9_c0 ;
	default :
		rl_a82_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a83_d9_c5 or RG_rl_a83_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a83_t5 = RG_rl_a83_d9_c0 ;
	3'h1 :
		rl_a83_t5 = RG_rl_a83_d9_c0 ;
	3'h2 :
		rl_a83_t5 = RG_rl_a83_d9_c0 ;
	3'h3 :
		rl_a83_t5 = RG_rl_a83_d9_c0 ;
	3'h4 :
		rl_a83_t5 = RG_rl_a83_d9_c0 ;
	3'h5 :
		rl_a83_t5 = RG_rl_a83_d9_c5 ;
	3'h6 :
		rl_a83_t5 = RG_rl_a83_d9_c0 ;
	3'h7 :
		rl_a83_t5 = RG_rl_a83_d9_c0 ;
	default :
		rl_a83_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a84_d9_c5 or RG_rl_a84_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a84_t5 = RG_rl_a84_d9_c0 ;
	3'h1 :
		rl_a84_t5 = RG_rl_a84_d9_c0 ;
	3'h2 :
		rl_a84_t5 = RG_rl_a84_d9_c0 ;
	3'h3 :
		rl_a84_t5 = RG_rl_a84_d9_c0 ;
	3'h4 :
		rl_a84_t5 = RG_rl_a84_d9_c0 ;
	3'h5 :
		rl_a84_t5 = RG_rl_a84_d9_c5 ;
	3'h6 :
		rl_a84_t5 = RG_rl_a84_d9_c0 ;
	3'h7 :
		rl_a84_t5 = RG_rl_a84_d9_c0 ;
	default :
		rl_a84_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a85_d9_c5 or RG_rl_a85_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a85_t5 = RG_rl_a85_d9_c0 ;
	3'h1 :
		rl_a85_t5 = RG_rl_a85_d9_c0 ;
	3'h2 :
		rl_a85_t5 = RG_rl_a85_d9_c0 ;
	3'h3 :
		rl_a85_t5 = RG_rl_a85_d9_c0 ;
	3'h4 :
		rl_a85_t5 = RG_rl_a85_d9_c0 ;
	3'h5 :
		rl_a85_t5 = RG_rl_a85_d9_c5 ;
	3'h6 :
		rl_a85_t5 = RG_rl_a85_d9_c0 ;
	3'h7 :
		rl_a85_t5 = RG_rl_a85_d9_c0 ;
	default :
		rl_a85_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a86_d9_c5 or RG_rl_a86_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a86_t5 = RG_rl_a86_d9_c0 ;
	3'h1 :
		rl_a86_t5 = RG_rl_a86_d9_c0 ;
	3'h2 :
		rl_a86_t5 = RG_rl_a86_d9_c0 ;
	3'h3 :
		rl_a86_t5 = RG_rl_a86_d9_c0 ;
	3'h4 :
		rl_a86_t5 = RG_rl_a86_d9_c0 ;
	3'h5 :
		rl_a86_t5 = RG_rl_a86_d9_c5 ;
	3'h6 :
		rl_a86_t5 = RG_rl_a86_d9_c0 ;
	3'h7 :
		rl_a86_t5 = RG_rl_a86_d9_c0 ;
	default :
		rl_a86_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a87_d9_c5 or RG_rl_a87_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a87_t5 = RG_rl_a87_d9_c0 ;
	3'h1 :
		rl_a87_t5 = RG_rl_a87_d9_c0 ;
	3'h2 :
		rl_a87_t5 = RG_rl_a87_d9_c0 ;
	3'h3 :
		rl_a87_t5 = RG_rl_a87_d9_c0 ;
	3'h4 :
		rl_a87_t5 = RG_rl_a87_d9_c0 ;
	3'h5 :
		rl_a87_t5 = RG_rl_a87_d9_c5 ;
	3'h6 :
		rl_a87_t5 = RG_rl_a87_d9_c0 ;
	3'h7 :
		rl_a87_t5 = RG_rl_a87_d9_c0 ;
	default :
		rl_a87_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a88_d9_c5 or RG_rl_a88_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a88_t5 = RG_rl_a88_d9_c0 ;
	3'h1 :
		rl_a88_t5 = RG_rl_a88_d9_c0 ;
	3'h2 :
		rl_a88_t5 = RG_rl_a88_d9_c0 ;
	3'h3 :
		rl_a88_t5 = RG_rl_a88_d9_c0 ;
	3'h4 :
		rl_a88_t5 = RG_rl_a88_d9_c0 ;
	3'h5 :
		rl_a88_t5 = RG_rl_a88_d9_c5 ;
	3'h6 :
		rl_a88_t5 = RG_rl_a88_d9_c0 ;
	3'h7 :
		rl_a88_t5 = RG_rl_a88_d9_c0 ;
	default :
		rl_a88_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a89_d9_c5 or RG_rl_a89_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a89_t5 = RG_rl_a89_d9_c0 ;
	3'h1 :
		rl_a89_t5 = RG_rl_a89_d9_c0 ;
	3'h2 :
		rl_a89_t5 = RG_rl_a89_d9_c0 ;
	3'h3 :
		rl_a89_t5 = RG_rl_a89_d9_c0 ;
	3'h4 :
		rl_a89_t5 = RG_rl_a89_d9_c0 ;
	3'h5 :
		rl_a89_t5 = RG_rl_a89_d9_c5 ;
	3'h6 :
		rl_a89_t5 = RG_rl_a89_d9_c0 ;
	3'h7 :
		rl_a89_t5 = RG_rl_a89_d9_c0 ;
	default :
		rl_a89_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a90_d9_c5 or RG_rl_a90_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a90_t5 = RG_rl_a90_d9_c0 ;
	3'h1 :
		rl_a90_t5 = RG_rl_a90_d9_c0 ;
	3'h2 :
		rl_a90_t5 = RG_rl_a90_d9_c0 ;
	3'h3 :
		rl_a90_t5 = RG_rl_a90_d9_c0 ;
	3'h4 :
		rl_a90_t5 = RG_rl_a90_d9_c0 ;
	3'h5 :
		rl_a90_t5 = RG_rl_a90_d9_c5 ;
	3'h6 :
		rl_a90_t5 = RG_rl_a90_d9_c0 ;
	3'h7 :
		rl_a90_t5 = RG_rl_a90_d9_c0 ;
	default :
		rl_a90_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a91_d9_c5 or RG_rl_a91_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a91_t5 = RG_rl_a91_d9_c0 ;
	3'h1 :
		rl_a91_t5 = RG_rl_a91_d9_c0 ;
	3'h2 :
		rl_a91_t5 = RG_rl_a91_d9_c0 ;
	3'h3 :
		rl_a91_t5 = RG_rl_a91_d9_c0 ;
	3'h4 :
		rl_a91_t5 = RG_rl_a91_d9_c0 ;
	3'h5 :
		rl_a91_t5 = RG_rl_a91_d9_c5 ;
	3'h6 :
		rl_a91_t5 = RG_rl_a91_d9_c0 ;
	3'h7 :
		rl_a91_t5 = RG_rl_a91_d9_c0 ;
	default :
		rl_a91_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a92_d9_c5 or RG_rl_a92_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a92_t5 = RG_rl_a92_d9_c0 ;
	3'h1 :
		rl_a92_t5 = RG_rl_a92_d9_c0 ;
	3'h2 :
		rl_a92_t5 = RG_rl_a92_d9_c0 ;
	3'h3 :
		rl_a92_t5 = RG_rl_a92_d9_c0 ;
	3'h4 :
		rl_a92_t5 = RG_rl_a92_d9_c0 ;
	3'h5 :
		rl_a92_t5 = RG_rl_a92_d9_c5 ;
	3'h6 :
		rl_a92_t5 = RG_rl_a92_d9_c0 ;
	3'h7 :
		rl_a92_t5 = RG_rl_a92_d9_c0 ;
	default :
		rl_a92_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a93_d9_c5 or RG_rl_a93_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a93_t5 = RG_rl_a93_d9_c0 ;
	3'h1 :
		rl_a93_t5 = RG_rl_a93_d9_c0 ;
	3'h2 :
		rl_a93_t5 = RG_rl_a93_d9_c0 ;
	3'h3 :
		rl_a93_t5 = RG_rl_a93_d9_c0 ;
	3'h4 :
		rl_a93_t5 = RG_rl_a93_d9_c0 ;
	3'h5 :
		rl_a93_t5 = RG_rl_a93_d9_c5 ;
	3'h6 :
		rl_a93_t5 = RG_rl_a93_d9_c0 ;
	3'h7 :
		rl_a93_t5 = RG_rl_a93_d9_c0 ;
	default :
		rl_a93_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a94_d9_c5 or RG_rl_a94_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a94_t5 = RG_rl_a94_d9_c0 ;
	3'h1 :
		rl_a94_t5 = RG_rl_a94_d9_c0 ;
	3'h2 :
		rl_a94_t5 = RG_rl_a94_d9_c0 ;
	3'h3 :
		rl_a94_t5 = RG_rl_a94_d9_c0 ;
	3'h4 :
		rl_a94_t5 = RG_rl_a94_d9_c0 ;
	3'h5 :
		rl_a94_t5 = RG_rl_a94_d9_c5 ;
	3'h6 :
		rl_a94_t5 = RG_rl_a94_d9_c0 ;
	3'h7 :
		rl_a94_t5 = RG_rl_a94_d9_c0 ;
	default :
		rl_a94_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a95_d9_c5 or RG_rl_a95_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a95_t5 = RG_rl_a95_d9_c0 ;
	3'h1 :
		rl_a95_t5 = RG_rl_a95_d9_c0 ;
	3'h2 :
		rl_a95_t5 = RG_rl_a95_d9_c0 ;
	3'h3 :
		rl_a95_t5 = RG_rl_a95_d9_c0 ;
	3'h4 :
		rl_a95_t5 = RG_rl_a95_d9_c0 ;
	3'h5 :
		rl_a95_t5 = RG_rl_a95_d9_c5 ;
	3'h6 :
		rl_a95_t5 = RG_rl_a95_d9_c0 ;
	3'h7 :
		rl_a95_t5 = RG_rl_a95_d9_c0 ;
	default :
		rl_a95_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a96_d9_c6 or RG_rl_a96_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a96_t5 = RG_rl_a96_d9_c0 ;
	3'h1 :
		rl_a96_t5 = RG_rl_a96_d9_c0 ;
	3'h2 :
		rl_a96_t5 = RG_rl_a96_d9_c0 ;
	3'h3 :
		rl_a96_t5 = RG_rl_a96_d9_c0 ;
	3'h4 :
		rl_a96_t5 = RG_rl_a96_d9_c0 ;
	3'h5 :
		rl_a96_t5 = RG_rl_a96_d9_c0 ;
	3'h6 :
		rl_a96_t5 = RG_rl_a96_d9_c6 ;
	3'h7 :
		rl_a96_t5 = RG_rl_a96_d9_c0 ;
	default :
		rl_a96_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a97_d9_c6 or RG_rl_a97_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a97_t5 = RG_rl_a97_d9_c0 ;
	3'h1 :
		rl_a97_t5 = RG_rl_a97_d9_c0 ;
	3'h2 :
		rl_a97_t5 = RG_rl_a97_d9_c0 ;
	3'h3 :
		rl_a97_t5 = RG_rl_a97_d9_c0 ;
	3'h4 :
		rl_a97_t5 = RG_rl_a97_d9_c0 ;
	3'h5 :
		rl_a97_t5 = RG_rl_a97_d9_c0 ;
	3'h6 :
		rl_a97_t5 = RG_rl_a97_d9_c6 ;
	3'h7 :
		rl_a97_t5 = RG_rl_a97_d9_c0 ;
	default :
		rl_a97_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a98_d9_c6 or RG_rl_a98_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a98_t5 = RG_rl_a98_d9_c0 ;
	3'h1 :
		rl_a98_t5 = RG_rl_a98_d9_c0 ;
	3'h2 :
		rl_a98_t5 = RG_rl_a98_d9_c0 ;
	3'h3 :
		rl_a98_t5 = RG_rl_a98_d9_c0 ;
	3'h4 :
		rl_a98_t5 = RG_rl_a98_d9_c0 ;
	3'h5 :
		rl_a98_t5 = RG_rl_a98_d9_c0 ;
	3'h6 :
		rl_a98_t5 = RG_rl_a98_d9_c6 ;
	3'h7 :
		rl_a98_t5 = RG_rl_a98_d9_c0 ;
	default :
		rl_a98_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a99_d9_c6 or RG_rl_a99_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a99_t5 = RG_rl_a99_d9_c0 ;
	3'h1 :
		rl_a99_t5 = RG_rl_a99_d9_c0 ;
	3'h2 :
		rl_a99_t5 = RG_rl_a99_d9_c0 ;
	3'h3 :
		rl_a99_t5 = RG_rl_a99_d9_c0 ;
	3'h4 :
		rl_a99_t5 = RG_rl_a99_d9_c0 ;
	3'h5 :
		rl_a99_t5 = RG_rl_a99_d9_c0 ;
	3'h6 :
		rl_a99_t5 = RG_rl_a99_d9_c6 ;
	3'h7 :
		rl_a99_t5 = RG_rl_a99_d9_c0 ;
	default :
		rl_a99_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a100_d9_c6 or RG_rl_a100_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a100_t5 = RG_rl_a100_d9_c0 ;
	3'h1 :
		rl_a100_t5 = RG_rl_a100_d9_c0 ;
	3'h2 :
		rl_a100_t5 = RG_rl_a100_d9_c0 ;
	3'h3 :
		rl_a100_t5 = RG_rl_a100_d9_c0 ;
	3'h4 :
		rl_a100_t5 = RG_rl_a100_d9_c0 ;
	3'h5 :
		rl_a100_t5 = RG_rl_a100_d9_c0 ;
	3'h6 :
		rl_a100_t5 = RG_rl_a100_d9_c6 ;
	3'h7 :
		rl_a100_t5 = RG_rl_a100_d9_c0 ;
	default :
		rl_a100_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a101_d9_c6 or RG_rl_a101_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a101_t5 = RG_rl_a101_d9_c0 ;
	3'h1 :
		rl_a101_t5 = RG_rl_a101_d9_c0 ;
	3'h2 :
		rl_a101_t5 = RG_rl_a101_d9_c0 ;
	3'h3 :
		rl_a101_t5 = RG_rl_a101_d9_c0 ;
	3'h4 :
		rl_a101_t5 = RG_rl_a101_d9_c0 ;
	3'h5 :
		rl_a101_t5 = RG_rl_a101_d9_c0 ;
	3'h6 :
		rl_a101_t5 = RG_rl_a101_d9_c6 ;
	3'h7 :
		rl_a101_t5 = RG_rl_a101_d9_c0 ;
	default :
		rl_a101_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a102_d9_c6 or RG_rl_a102_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a102_t5 = RG_rl_a102_d9_c0 ;
	3'h1 :
		rl_a102_t5 = RG_rl_a102_d9_c0 ;
	3'h2 :
		rl_a102_t5 = RG_rl_a102_d9_c0 ;
	3'h3 :
		rl_a102_t5 = RG_rl_a102_d9_c0 ;
	3'h4 :
		rl_a102_t5 = RG_rl_a102_d9_c0 ;
	3'h5 :
		rl_a102_t5 = RG_rl_a102_d9_c0 ;
	3'h6 :
		rl_a102_t5 = RG_rl_a102_d9_c6 ;
	3'h7 :
		rl_a102_t5 = RG_rl_a102_d9_c0 ;
	default :
		rl_a102_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a103_d9_c6 or RG_rl_a103_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a103_t5 = RG_rl_a103_d9_c0 ;
	3'h1 :
		rl_a103_t5 = RG_rl_a103_d9_c0 ;
	3'h2 :
		rl_a103_t5 = RG_rl_a103_d9_c0 ;
	3'h3 :
		rl_a103_t5 = RG_rl_a103_d9_c0 ;
	3'h4 :
		rl_a103_t5 = RG_rl_a103_d9_c0 ;
	3'h5 :
		rl_a103_t5 = RG_rl_a103_d9_c0 ;
	3'h6 :
		rl_a103_t5 = RG_rl_a103_d9_c6 ;
	3'h7 :
		rl_a103_t5 = RG_rl_a103_d9_c0 ;
	default :
		rl_a103_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a104_d9_c6 or RG_rl_a104_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a104_t5 = RG_rl_a104_d9_c0 ;
	3'h1 :
		rl_a104_t5 = RG_rl_a104_d9_c0 ;
	3'h2 :
		rl_a104_t5 = RG_rl_a104_d9_c0 ;
	3'h3 :
		rl_a104_t5 = RG_rl_a104_d9_c0 ;
	3'h4 :
		rl_a104_t5 = RG_rl_a104_d9_c0 ;
	3'h5 :
		rl_a104_t5 = RG_rl_a104_d9_c0 ;
	3'h6 :
		rl_a104_t5 = RG_rl_a104_d9_c6 ;
	3'h7 :
		rl_a104_t5 = RG_rl_a104_d9_c0 ;
	default :
		rl_a104_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a105_d9_c6 or RG_rl_a105_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a105_t5 = RG_rl_a105_d9_c0 ;
	3'h1 :
		rl_a105_t5 = RG_rl_a105_d9_c0 ;
	3'h2 :
		rl_a105_t5 = RG_rl_a105_d9_c0 ;
	3'h3 :
		rl_a105_t5 = RG_rl_a105_d9_c0 ;
	3'h4 :
		rl_a105_t5 = RG_rl_a105_d9_c0 ;
	3'h5 :
		rl_a105_t5 = RG_rl_a105_d9_c0 ;
	3'h6 :
		rl_a105_t5 = RG_rl_a105_d9_c6 ;
	3'h7 :
		rl_a105_t5 = RG_rl_a105_d9_c0 ;
	default :
		rl_a105_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a106_d9_c6 or RG_rl_a106_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a106_t5 = RG_rl_a106_d9_c0 ;
	3'h1 :
		rl_a106_t5 = RG_rl_a106_d9_c0 ;
	3'h2 :
		rl_a106_t5 = RG_rl_a106_d9_c0 ;
	3'h3 :
		rl_a106_t5 = RG_rl_a106_d9_c0 ;
	3'h4 :
		rl_a106_t5 = RG_rl_a106_d9_c0 ;
	3'h5 :
		rl_a106_t5 = RG_rl_a106_d9_c0 ;
	3'h6 :
		rl_a106_t5 = RG_rl_a106_d9_c6 ;
	3'h7 :
		rl_a106_t5 = RG_rl_a106_d9_c0 ;
	default :
		rl_a106_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a107_d9_c6 or RG_rl_a107_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a107_t5 = RG_rl_a107_d9_c0 ;
	3'h1 :
		rl_a107_t5 = RG_rl_a107_d9_c0 ;
	3'h2 :
		rl_a107_t5 = RG_rl_a107_d9_c0 ;
	3'h3 :
		rl_a107_t5 = RG_rl_a107_d9_c0 ;
	3'h4 :
		rl_a107_t5 = RG_rl_a107_d9_c0 ;
	3'h5 :
		rl_a107_t5 = RG_rl_a107_d9_c0 ;
	3'h6 :
		rl_a107_t5 = RG_rl_a107_d9_c6 ;
	3'h7 :
		rl_a107_t5 = RG_rl_a107_d9_c0 ;
	default :
		rl_a107_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a108_d9_c6 or RG_rl_a108_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a108_t5 = RG_rl_a108_d9_c0 ;
	3'h1 :
		rl_a108_t5 = RG_rl_a108_d9_c0 ;
	3'h2 :
		rl_a108_t5 = RG_rl_a108_d9_c0 ;
	3'h3 :
		rl_a108_t5 = RG_rl_a108_d9_c0 ;
	3'h4 :
		rl_a108_t5 = RG_rl_a108_d9_c0 ;
	3'h5 :
		rl_a108_t5 = RG_rl_a108_d9_c0 ;
	3'h6 :
		rl_a108_t5 = RG_rl_a108_d9_c6 ;
	3'h7 :
		rl_a108_t5 = RG_rl_a108_d9_c0 ;
	default :
		rl_a108_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a109_d9_c6 or RG_rl_a109_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a109_t5 = RG_rl_a109_d9_c0 ;
	3'h1 :
		rl_a109_t5 = RG_rl_a109_d9_c0 ;
	3'h2 :
		rl_a109_t5 = RG_rl_a109_d9_c0 ;
	3'h3 :
		rl_a109_t5 = RG_rl_a109_d9_c0 ;
	3'h4 :
		rl_a109_t5 = RG_rl_a109_d9_c0 ;
	3'h5 :
		rl_a109_t5 = RG_rl_a109_d9_c0 ;
	3'h6 :
		rl_a109_t5 = RG_rl_a109_d9_c6 ;
	3'h7 :
		rl_a109_t5 = RG_rl_a109_d9_c0 ;
	default :
		rl_a109_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a110_d9_c6 or RG_rl_a110_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a110_t5 = RG_rl_a110_d9_c0 ;
	3'h1 :
		rl_a110_t5 = RG_rl_a110_d9_c0 ;
	3'h2 :
		rl_a110_t5 = RG_rl_a110_d9_c0 ;
	3'h3 :
		rl_a110_t5 = RG_rl_a110_d9_c0 ;
	3'h4 :
		rl_a110_t5 = RG_rl_a110_d9_c0 ;
	3'h5 :
		rl_a110_t5 = RG_rl_a110_d9_c0 ;
	3'h6 :
		rl_a110_t5 = RG_rl_a110_d9_c6 ;
	3'h7 :
		rl_a110_t5 = RG_rl_a110_d9_c0 ;
	default :
		rl_a110_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a111_d9_c6 or RG_rl_a111_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a111_t5 = RG_rl_a111_d9_c0 ;
	3'h1 :
		rl_a111_t5 = RG_rl_a111_d9_c0 ;
	3'h2 :
		rl_a111_t5 = RG_rl_a111_d9_c0 ;
	3'h3 :
		rl_a111_t5 = RG_rl_a111_d9_c0 ;
	3'h4 :
		rl_a111_t5 = RG_rl_a111_d9_c0 ;
	3'h5 :
		rl_a111_t5 = RG_rl_a111_d9_c0 ;
	3'h6 :
		rl_a111_t5 = RG_rl_a111_d9_c6 ;
	3'h7 :
		rl_a111_t5 = RG_rl_a111_d9_c0 ;
	default :
		rl_a111_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a112_d9_c7 or RG_rl_a112_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a112_t5 = RG_rl_a112_d9_c0 ;
	3'h1 :
		rl_a112_t5 = RG_rl_a112_d9_c0 ;
	3'h2 :
		rl_a112_t5 = RG_rl_a112_d9_c0 ;
	3'h3 :
		rl_a112_t5 = RG_rl_a112_d9_c0 ;
	3'h4 :
		rl_a112_t5 = RG_rl_a112_d9_c0 ;
	3'h5 :
		rl_a112_t5 = RG_rl_a112_d9_c0 ;
	3'h6 :
		rl_a112_t5 = RG_rl_a112_d9_c0 ;
	3'h7 :
		rl_a112_t5 = RG_rl_a112_d9_c7 ;
	default :
		rl_a112_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a113_d9_c7 or RG_rl_a113_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a113_t5 = RG_rl_a113_d9_c0 ;
	3'h1 :
		rl_a113_t5 = RG_rl_a113_d9_c0 ;
	3'h2 :
		rl_a113_t5 = RG_rl_a113_d9_c0 ;
	3'h3 :
		rl_a113_t5 = RG_rl_a113_d9_c0 ;
	3'h4 :
		rl_a113_t5 = RG_rl_a113_d9_c0 ;
	3'h5 :
		rl_a113_t5 = RG_rl_a113_d9_c0 ;
	3'h6 :
		rl_a113_t5 = RG_rl_a113_d9_c0 ;
	3'h7 :
		rl_a113_t5 = RG_rl_a113_d9_c7 ;
	default :
		rl_a113_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a114_d9_c7 or RG_rl_a114_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a114_t5 = RG_rl_a114_d9_c0 ;
	3'h1 :
		rl_a114_t5 = RG_rl_a114_d9_c0 ;
	3'h2 :
		rl_a114_t5 = RG_rl_a114_d9_c0 ;
	3'h3 :
		rl_a114_t5 = RG_rl_a114_d9_c0 ;
	3'h4 :
		rl_a114_t5 = RG_rl_a114_d9_c0 ;
	3'h5 :
		rl_a114_t5 = RG_rl_a114_d9_c0 ;
	3'h6 :
		rl_a114_t5 = RG_rl_a114_d9_c0 ;
	3'h7 :
		rl_a114_t5 = RG_rl_a114_d9_c7 ;
	default :
		rl_a114_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a115_d9_c7 or RG_rl_a115_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a115_t5 = RG_rl_a115_d9_c0 ;
	3'h1 :
		rl_a115_t5 = RG_rl_a115_d9_c0 ;
	3'h2 :
		rl_a115_t5 = RG_rl_a115_d9_c0 ;
	3'h3 :
		rl_a115_t5 = RG_rl_a115_d9_c0 ;
	3'h4 :
		rl_a115_t5 = RG_rl_a115_d9_c0 ;
	3'h5 :
		rl_a115_t5 = RG_rl_a115_d9_c0 ;
	3'h6 :
		rl_a115_t5 = RG_rl_a115_d9_c0 ;
	3'h7 :
		rl_a115_t5 = RG_rl_a115_d9_c7 ;
	default :
		rl_a115_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a116_d9_c7 or RG_rl_a116_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a116_t5 = RG_rl_a116_d9_c0 ;
	3'h1 :
		rl_a116_t5 = RG_rl_a116_d9_c0 ;
	3'h2 :
		rl_a116_t5 = RG_rl_a116_d9_c0 ;
	3'h3 :
		rl_a116_t5 = RG_rl_a116_d9_c0 ;
	3'h4 :
		rl_a116_t5 = RG_rl_a116_d9_c0 ;
	3'h5 :
		rl_a116_t5 = RG_rl_a116_d9_c0 ;
	3'h6 :
		rl_a116_t5 = RG_rl_a116_d9_c0 ;
	3'h7 :
		rl_a116_t5 = RG_rl_a116_d9_c7 ;
	default :
		rl_a116_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a117_d9_c7 or RG_rl_a117_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a117_t5 = RG_rl_a117_d9_c0 ;
	3'h1 :
		rl_a117_t5 = RG_rl_a117_d9_c0 ;
	3'h2 :
		rl_a117_t5 = RG_rl_a117_d9_c0 ;
	3'h3 :
		rl_a117_t5 = RG_rl_a117_d9_c0 ;
	3'h4 :
		rl_a117_t5 = RG_rl_a117_d9_c0 ;
	3'h5 :
		rl_a117_t5 = RG_rl_a117_d9_c0 ;
	3'h6 :
		rl_a117_t5 = RG_rl_a117_d9_c0 ;
	3'h7 :
		rl_a117_t5 = RG_rl_a117_d9_c7 ;
	default :
		rl_a117_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a118_d9_c7 or RG_rl_a118_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a118_t5 = RG_rl_a118_d9_c0 ;
	3'h1 :
		rl_a118_t5 = RG_rl_a118_d9_c0 ;
	3'h2 :
		rl_a118_t5 = RG_rl_a118_d9_c0 ;
	3'h3 :
		rl_a118_t5 = RG_rl_a118_d9_c0 ;
	3'h4 :
		rl_a118_t5 = RG_rl_a118_d9_c0 ;
	3'h5 :
		rl_a118_t5 = RG_rl_a118_d9_c0 ;
	3'h6 :
		rl_a118_t5 = RG_rl_a118_d9_c0 ;
	3'h7 :
		rl_a118_t5 = RG_rl_a118_d9_c7 ;
	default :
		rl_a118_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a119_d9_c7 or RG_rl_a119_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a119_t5 = RG_rl_a119_d9_c0 ;
	3'h1 :
		rl_a119_t5 = RG_rl_a119_d9_c0 ;
	3'h2 :
		rl_a119_t5 = RG_rl_a119_d9_c0 ;
	3'h3 :
		rl_a119_t5 = RG_rl_a119_d9_c0 ;
	3'h4 :
		rl_a119_t5 = RG_rl_a119_d9_c0 ;
	3'h5 :
		rl_a119_t5 = RG_rl_a119_d9_c0 ;
	3'h6 :
		rl_a119_t5 = RG_rl_a119_d9_c0 ;
	3'h7 :
		rl_a119_t5 = RG_rl_a119_d9_c7 ;
	default :
		rl_a119_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a120_d9_c7 or RG_rl_a120_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a120_t5 = RG_rl_a120_d9_c0 ;
	3'h1 :
		rl_a120_t5 = RG_rl_a120_d9_c0 ;
	3'h2 :
		rl_a120_t5 = RG_rl_a120_d9_c0 ;
	3'h3 :
		rl_a120_t5 = RG_rl_a120_d9_c0 ;
	3'h4 :
		rl_a120_t5 = RG_rl_a120_d9_c0 ;
	3'h5 :
		rl_a120_t5 = RG_rl_a120_d9_c0 ;
	3'h6 :
		rl_a120_t5 = RG_rl_a120_d9_c0 ;
	3'h7 :
		rl_a120_t5 = RG_rl_a120_d9_c7 ;
	default :
		rl_a120_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a121_d9_c7 or RG_rl_a121_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a121_t5 = RG_rl_a121_d9_c0 ;
	3'h1 :
		rl_a121_t5 = RG_rl_a121_d9_c0 ;
	3'h2 :
		rl_a121_t5 = RG_rl_a121_d9_c0 ;
	3'h3 :
		rl_a121_t5 = RG_rl_a121_d9_c0 ;
	3'h4 :
		rl_a121_t5 = RG_rl_a121_d9_c0 ;
	3'h5 :
		rl_a121_t5 = RG_rl_a121_d9_c0 ;
	3'h6 :
		rl_a121_t5 = RG_rl_a121_d9_c0 ;
	3'h7 :
		rl_a121_t5 = RG_rl_a121_d9_c7 ;
	default :
		rl_a121_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a122_d9_c7 or RG_rl_a122_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a122_t5 = RG_rl_a122_d9_c0 ;
	3'h1 :
		rl_a122_t5 = RG_rl_a122_d9_c0 ;
	3'h2 :
		rl_a122_t5 = RG_rl_a122_d9_c0 ;
	3'h3 :
		rl_a122_t5 = RG_rl_a122_d9_c0 ;
	3'h4 :
		rl_a122_t5 = RG_rl_a122_d9_c0 ;
	3'h5 :
		rl_a122_t5 = RG_rl_a122_d9_c0 ;
	3'h6 :
		rl_a122_t5 = RG_rl_a122_d9_c0 ;
	3'h7 :
		rl_a122_t5 = RG_rl_a122_d9_c7 ;
	default :
		rl_a122_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a123_d9_c7 or RG_rl_a123_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a123_t5 = RG_rl_a123_d9_c0 ;
	3'h1 :
		rl_a123_t5 = RG_rl_a123_d9_c0 ;
	3'h2 :
		rl_a123_t5 = RG_rl_a123_d9_c0 ;
	3'h3 :
		rl_a123_t5 = RG_rl_a123_d9_c0 ;
	3'h4 :
		rl_a123_t5 = RG_rl_a123_d9_c0 ;
	3'h5 :
		rl_a123_t5 = RG_rl_a123_d9_c0 ;
	3'h6 :
		rl_a123_t5 = RG_rl_a123_d9_c0 ;
	3'h7 :
		rl_a123_t5 = RG_rl_a123_d9_c7 ;
	default :
		rl_a123_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a124_d9_c7 or RG_rl_a124_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a124_t5 = RG_rl_a124_d9_c0 ;
	3'h1 :
		rl_a124_t5 = RG_rl_a124_d9_c0 ;
	3'h2 :
		rl_a124_t5 = RG_rl_a124_d9_c0 ;
	3'h3 :
		rl_a124_t5 = RG_rl_a124_d9_c0 ;
	3'h4 :
		rl_a124_t5 = RG_rl_a124_d9_c0 ;
	3'h5 :
		rl_a124_t5 = RG_rl_a124_d9_c0 ;
	3'h6 :
		rl_a124_t5 = RG_rl_a124_d9_c0 ;
	3'h7 :
		rl_a124_t5 = RG_rl_a124_d9_c7 ;
	default :
		rl_a124_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a125_d9_c7 or RG_rl_a125_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a125_t5 = RG_rl_a125_d9_c0 ;
	3'h1 :
		rl_a125_t5 = RG_rl_a125_d9_c0 ;
	3'h2 :
		rl_a125_t5 = RG_rl_a125_d9_c0 ;
	3'h3 :
		rl_a125_t5 = RG_rl_a125_d9_c0 ;
	3'h4 :
		rl_a125_t5 = RG_rl_a125_d9_c0 ;
	3'h5 :
		rl_a125_t5 = RG_rl_a125_d9_c0 ;
	3'h6 :
		rl_a125_t5 = RG_rl_a125_d9_c0 ;
	3'h7 :
		rl_a125_t5 = RG_rl_a125_d9_c7 ;
	default :
		rl_a125_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a126_d9_c7 or RG_rl_a126_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a126_t5 = RG_rl_a126_d9_c0 ;
	3'h1 :
		rl_a126_t5 = RG_rl_a126_d9_c0 ;
	3'h2 :
		rl_a126_t5 = RG_rl_a126_d9_c0 ;
	3'h3 :
		rl_a126_t5 = RG_rl_a126_d9_c0 ;
	3'h4 :
		rl_a126_t5 = RG_rl_a126_d9_c0 ;
	3'h5 :
		rl_a126_t5 = RG_rl_a126_d9_c0 ;
	3'h6 :
		rl_a126_t5 = RG_rl_a126_d9_c0 ;
	3'h7 :
		rl_a126_t5 = RG_rl_a126_d9_c7 ;
	default :
		rl_a126_t5 = 9'hx ;
	endcase
always @ ( RG_rl_a127_d9_c7 or RG_rl_a127_d9_c0 or RG_k_01 )
	case ( RG_k_01 [6:4] )
	3'h0 :
		rl_a127_t5 = RG_rl_a127_d9_c0 ;
	3'h1 :
		rl_a127_t5 = RG_rl_a127_d9_c0 ;
	3'h2 :
		rl_a127_t5 = RG_rl_a127_d9_c0 ;
	3'h3 :
		rl_a127_t5 = RG_rl_a127_d9_c0 ;
	3'h4 :
		rl_a127_t5 = RG_rl_a127_d9_c0 ;
	3'h5 :
		rl_a127_t5 = RG_rl_a127_d9_c0 ;
	3'h6 :
		rl_a127_t5 = RG_rl_a127_d9_c0 ;
	3'h7 :
		rl_a127_t5 = RG_rl_a127_d9_c7 ;
	default :
		rl_a127_t5 = 9'hx ;
	endcase
assign	M_190 = ~|rl_a00_t4 ;	// line#=../rle.cpp:77,78
assign	M_191 = ~|rl_a01_t4 ;	// line#=../rle.cpp:77,78
assign	M_192 = ~|rl_a02_t4 ;	// line#=../rle.cpp:77,78
assign	M_193 = ~|rl_a03_t4 ;	// line#=../rle.cpp:77,78
assign	M_194 = ~|rl_a04_t4 ;	// line#=../rle.cpp:77,78
assign	M_195 = ~|rl_a05_t4 ;	// line#=../rle.cpp:77,78
assign	M_196 = ~|rl_a06_t4 ;	// line#=../rle.cpp:77,78
assign	M_197 = ~|rl_a07_t4 ;	// line#=../rle.cpp:77,78
assign	M_198 = ~|rl_a08_t4 ;	// line#=../rle.cpp:77,78
assign	M_199 = ~|rl_a09_t4 ;	// line#=../rle.cpp:77,78
assign	M_200 = ~|rl_a10_t4 ;	// line#=../rle.cpp:77,78
assign	M_201 = ~|rl_a11_t4 ;	// line#=../rle.cpp:77,78
assign	M_202 = ~|rl_a12_t4 ;	// line#=../rle.cpp:77,78
assign	M_203 = ~|rl_a13_t4 ;	// line#=../rle.cpp:77,78
assign	M_204 = ~|rl_a14_t4 ;	// line#=../rle.cpp:77,78
assign	M_205 = ~|rl_a15_t4 ;	// line#=../rle.cpp:77,78
always @ ( M_205 or M_204 or M_203 or M_202 or M_201 or M_200 or M_199 or M_198 or 
	M_197 or M_196 or M_195 or M_194 or M_193 or M_192 or M_191 or M_190 or 
	decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot [3:0] )
	4'h0 :
		RG_M_14_d10_c0_t = M_190 ;	// line#=../rle.cpp:77,78
	4'h1 :
		RG_M_14_d10_c0_t = M_191 ;	// line#=../rle.cpp:77,78
	4'h2 :
		RG_M_14_d10_c0_t = M_192 ;	// line#=../rle.cpp:77,78
	4'h3 :
		RG_M_14_d10_c0_t = M_193 ;	// line#=../rle.cpp:77,78
	4'h4 :
		RG_M_14_d10_c0_t = M_194 ;	// line#=../rle.cpp:77,78
	4'h5 :
		RG_M_14_d10_c0_t = M_195 ;	// line#=../rle.cpp:77,78
	4'h6 :
		RG_M_14_d10_c0_t = M_196 ;	// line#=../rle.cpp:77,78
	4'h7 :
		RG_M_14_d10_c0_t = M_197 ;	// line#=../rle.cpp:77,78
	4'h8 :
		RG_M_14_d10_c0_t = M_198 ;	// line#=../rle.cpp:77,78
	4'h9 :
		RG_M_14_d10_c0_t = M_199 ;	// line#=../rle.cpp:77,78
	4'ha :
		RG_M_14_d10_c0_t = M_200 ;	// line#=../rle.cpp:77,78
	4'hb :
		RG_M_14_d10_c0_t = M_201 ;	// line#=../rle.cpp:77,78
	4'hc :
		RG_M_14_d10_c0_t = M_202 ;	// line#=../rle.cpp:77,78
	4'hd :
		RG_M_14_d10_c0_t = M_203 ;	// line#=../rle.cpp:77,78
	4'he :
		RG_M_14_d10_c0_t = M_204 ;	// line#=../rle.cpp:77,78
	4'hf :
		RG_M_14_d10_c0_t = M_205 ;	// line#=../rle.cpp:77,78
	default :
		RG_M_14_d10_c0_t = 1'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_M_14_d10_c0 <= RG_M_14_d10_c0_t ;	// line#=../rle.cpp:77,78
assign	M_206 = ~|rl_a16_t4 ;	// line#=../rle.cpp:77,78
assign	M_207 = ~|rl_a17_t4 ;	// line#=../rle.cpp:77,78
assign	M_208 = ~|rl_a18_t4 ;	// line#=../rle.cpp:77,78
assign	M_209 = ~|rl_a19_t4 ;	// line#=../rle.cpp:77,78
assign	M_210 = ~|rl_a20_t4 ;	// line#=../rle.cpp:77,78
assign	M_211 = ~|rl_a21_t4 ;	// line#=../rle.cpp:77,78
assign	M_212 = ~|rl_a22_t4 ;	// line#=../rle.cpp:77,78
assign	M_213 = ~|rl_a23_t4 ;	// line#=../rle.cpp:77,78
assign	M_214 = ~|rl_a24_t4 ;	// line#=../rle.cpp:77,78
assign	M_215 = ~|rl_a25_t4 ;	// line#=../rle.cpp:77,78
assign	M_216 = ~|rl_a26_t4 ;	// line#=../rle.cpp:77,78
assign	M_217 = ~|rl_a27_t4 ;	// line#=../rle.cpp:77,78
assign	M_218 = ~|rl_a28_t4 ;	// line#=../rle.cpp:77,78
assign	M_219 = ~|rl_a29_t4 ;	// line#=../rle.cpp:77,78
assign	M_220 = ~|rl_a30_t4 ;	// line#=../rle.cpp:77,78
assign	M_221 = ~|rl_a31_t4 ;	// line#=../rle.cpp:77,78
always @ ( M_221 or M_220 or M_219 or M_218 or M_217 or M_216 or M_215 or M_214 or 
	M_213 or M_212 or M_211 or M_210 or M_209 or M_208 or M_207 or M_206 or 
	decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot [3:0] )
	4'h0 :
		RG_M_14_d10_c1_t = M_206 ;	// line#=../rle.cpp:77,78
	4'h1 :
		RG_M_14_d10_c1_t = M_207 ;	// line#=../rle.cpp:77,78
	4'h2 :
		RG_M_14_d10_c1_t = M_208 ;	// line#=../rle.cpp:77,78
	4'h3 :
		RG_M_14_d10_c1_t = M_209 ;	// line#=../rle.cpp:77,78
	4'h4 :
		RG_M_14_d10_c1_t = M_210 ;	// line#=../rle.cpp:77,78
	4'h5 :
		RG_M_14_d10_c1_t = M_211 ;	// line#=../rle.cpp:77,78
	4'h6 :
		RG_M_14_d10_c1_t = M_212 ;	// line#=../rle.cpp:77,78
	4'h7 :
		RG_M_14_d10_c1_t = M_213 ;	// line#=../rle.cpp:77,78
	4'h8 :
		RG_M_14_d10_c1_t = M_214 ;	// line#=../rle.cpp:77,78
	4'h9 :
		RG_M_14_d10_c1_t = M_215 ;	// line#=../rle.cpp:77,78
	4'ha :
		RG_M_14_d10_c1_t = M_216 ;	// line#=../rle.cpp:77,78
	4'hb :
		RG_M_14_d10_c1_t = M_217 ;	// line#=../rle.cpp:77,78
	4'hc :
		RG_M_14_d10_c1_t = M_218 ;	// line#=../rle.cpp:77,78
	4'hd :
		RG_M_14_d10_c1_t = M_219 ;	// line#=../rle.cpp:77,78
	4'he :
		RG_M_14_d10_c1_t = M_220 ;	// line#=../rle.cpp:77,78
	4'hf :
		RG_M_14_d10_c1_t = M_221 ;	// line#=../rle.cpp:77,78
	default :
		RG_M_14_d10_c1_t = 1'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_M_14_d10_c1 <= RG_M_14_d10_c1_t ;	// line#=../rle.cpp:77,78
assign	M_222 = ~|rl_a32_t4 ;	// line#=../rle.cpp:77,78
assign	M_223 = ~|rl_a33_t4 ;	// line#=../rle.cpp:77,78
assign	M_224 = ~|rl_a34_t4 ;	// line#=../rle.cpp:77,78
assign	M_225 = ~|rl_a35_t4 ;	// line#=../rle.cpp:77,78
assign	M_226 = ~|rl_a36_t4 ;	// line#=../rle.cpp:77,78
assign	M_227 = ~|rl_a37_t4 ;	// line#=../rle.cpp:77,78
assign	M_228 = ~|rl_a38_t4 ;	// line#=../rle.cpp:77,78
assign	M_229 = ~|rl_a39_t4 ;	// line#=../rle.cpp:77,78
assign	M_230 = ~|rl_a40_t4 ;	// line#=../rle.cpp:77,78
assign	M_231 = ~|rl_a41_t4 ;	// line#=../rle.cpp:77,78
assign	M_232 = ~|rl_a42_t4 ;	// line#=../rle.cpp:77,78
assign	M_233 = ~|rl_a43_t4 ;	// line#=../rle.cpp:77,78
assign	M_234 = ~|rl_a44_t4 ;	// line#=../rle.cpp:77,78
assign	M_235 = ~|rl_a45_t4 ;	// line#=../rle.cpp:77,78
assign	M_236 = ~|rl_a46_t4 ;	// line#=../rle.cpp:77,78
assign	M_237 = ~|rl_a47_t4 ;	// line#=../rle.cpp:77,78
always @ ( M_237 or M_236 or M_235 or M_234 or M_233 or M_232 or M_231 or M_230 or 
	M_229 or M_228 or M_227 or M_226 or M_225 or M_224 or M_223 or M_222 or 
	decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot [3:0] )
	4'h0 :
		RG_M_14_d10_c2_t = M_222 ;	// line#=../rle.cpp:77,78
	4'h1 :
		RG_M_14_d10_c2_t = M_223 ;	// line#=../rle.cpp:77,78
	4'h2 :
		RG_M_14_d10_c2_t = M_224 ;	// line#=../rle.cpp:77,78
	4'h3 :
		RG_M_14_d10_c2_t = M_225 ;	// line#=../rle.cpp:77,78
	4'h4 :
		RG_M_14_d10_c2_t = M_226 ;	// line#=../rle.cpp:77,78
	4'h5 :
		RG_M_14_d10_c2_t = M_227 ;	// line#=../rle.cpp:77,78
	4'h6 :
		RG_M_14_d10_c2_t = M_228 ;	// line#=../rle.cpp:77,78
	4'h7 :
		RG_M_14_d10_c2_t = M_229 ;	// line#=../rle.cpp:77,78
	4'h8 :
		RG_M_14_d10_c2_t = M_230 ;	// line#=../rle.cpp:77,78
	4'h9 :
		RG_M_14_d10_c2_t = M_231 ;	// line#=../rle.cpp:77,78
	4'ha :
		RG_M_14_d10_c2_t = M_232 ;	// line#=../rle.cpp:77,78
	4'hb :
		RG_M_14_d10_c2_t = M_233 ;	// line#=../rle.cpp:77,78
	4'hc :
		RG_M_14_d10_c2_t = M_234 ;	// line#=../rle.cpp:77,78
	4'hd :
		RG_M_14_d10_c2_t = M_235 ;	// line#=../rle.cpp:77,78
	4'he :
		RG_M_14_d10_c2_t = M_236 ;	// line#=../rle.cpp:77,78
	4'hf :
		RG_M_14_d10_c2_t = M_237 ;	// line#=../rle.cpp:77,78
	default :
		RG_M_14_d10_c2_t = 1'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_M_14_d10_c2 <= RG_M_14_d10_c2_t ;	// line#=../rle.cpp:77,78
assign	M_238 = ~|rl_a48_t4 ;	// line#=../rle.cpp:77,78
assign	M_239 = ~|rl_a49_t4 ;	// line#=../rle.cpp:77,78
assign	M_240 = ~|rl_a50_t4 ;	// line#=../rle.cpp:77,78
assign	M_241 = ~|rl_a51_t4 ;	// line#=../rle.cpp:77,78
assign	M_242 = ~|rl_a52_t4 ;	// line#=../rle.cpp:77,78
assign	M_243 = ~|rl_a53_t4 ;	// line#=../rle.cpp:77,78
assign	M_244 = ~|rl_a54_t4 ;	// line#=../rle.cpp:77,78
assign	M_245 = ~|rl_a55_t4 ;	// line#=../rle.cpp:77,78
assign	M_246 = ~|rl_a56_t4 ;	// line#=../rle.cpp:77,78
assign	M_247 = ~|rl_a57_t4 ;	// line#=../rle.cpp:77,78
assign	M_248 = ~|rl_a58_t4 ;	// line#=../rle.cpp:77,78
assign	M_249 = ~|rl_a59_t4 ;	// line#=../rle.cpp:77,78
assign	M_250 = ~|rl_a60_t4 ;	// line#=../rle.cpp:77,78
assign	M_251 = ~|rl_a61_t4 ;	// line#=../rle.cpp:77,78
assign	M_252 = ~|rl_a62_t4 ;	// line#=../rle.cpp:77,78
assign	M_253 = ~|rl_a63_t4 ;	// line#=../rle.cpp:77,78
always @ ( M_253 or M_252 or M_251 or M_250 or M_249 or M_248 or M_247 or M_246 or 
	M_245 or M_244 or M_243 or M_242 or M_241 or M_240 or M_239 or M_238 or 
	decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot [3:0] )
	4'h0 :
		RG_M_14_d10_c3_t = M_238 ;	// line#=../rle.cpp:77,78
	4'h1 :
		RG_M_14_d10_c3_t = M_239 ;	// line#=../rle.cpp:77,78
	4'h2 :
		RG_M_14_d10_c3_t = M_240 ;	// line#=../rle.cpp:77,78
	4'h3 :
		RG_M_14_d10_c3_t = M_241 ;	// line#=../rle.cpp:77,78
	4'h4 :
		RG_M_14_d10_c3_t = M_242 ;	// line#=../rle.cpp:77,78
	4'h5 :
		RG_M_14_d10_c3_t = M_243 ;	// line#=../rle.cpp:77,78
	4'h6 :
		RG_M_14_d10_c3_t = M_244 ;	// line#=../rle.cpp:77,78
	4'h7 :
		RG_M_14_d10_c3_t = M_245 ;	// line#=../rle.cpp:77,78
	4'h8 :
		RG_M_14_d10_c3_t = M_246 ;	// line#=../rle.cpp:77,78
	4'h9 :
		RG_M_14_d10_c3_t = M_247 ;	// line#=../rle.cpp:77,78
	4'ha :
		RG_M_14_d10_c3_t = M_248 ;	// line#=../rle.cpp:77,78
	4'hb :
		RG_M_14_d10_c3_t = M_249 ;	// line#=../rle.cpp:77,78
	4'hc :
		RG_M_14_d10_c3_t = M_250 ;	// line#=../rle.cpp:77,78
	4'hd :
		RG_M_14_d10_c3_t = M_251 ;	// line#=../rle.cpp:77,78
	4'he :
		RG_M_14_d10_c3_t = M_252 ;	// line#=../rle.cpp:77,78
	4'hf :
		RG_M_14_d10_c3_t = M_253 ;	// line#=../rle.cpp:77,78
	default :
		RG_M_14_d10_c3_t = 1'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_M_14_d10_c3 <= RG_M_14_d10_c3_t ;	// line#=../rle.cpp:77,78
assign	M_254 = ~|rl_a64_t4 ;	// line#=../rle.cpp:77,78
assign	M_255 = ~|rl_a65_t4 ;	// line#=../rle.cpp:77,78
assign	M_256 = ~|rl_a66_t4 ;	// line#=../rle.cpp:77,78
assign	M_257 = ~|rl_a67_t4 ;	// line#=../rle.cpp:77,78
assign	M_258 = ~|rl_a68_t4 ;	// line#=../rle.cpp:77,78
assign	M_259 = ~|rl_a69_t4 ;	// line#=../rle.cpp:77,78
assign	M_260 = ~|rl_a70_t4 ;	// line#=../rle.cpp:77,78
assign	M_261 = ~|rl_a71_t4 ;	// line#=../rle.cpp:77,78
assign	M_262 = ~|rl_a72_t4 ;	// line#=../rle.cpp:77,78
assign	M_263 = ~|rl_a73_t4 ;	// line#=../rle.cpp:77,78
assign	M_264 = ~|rl_a74_t4 ;	// line#=../rle.cpp:77,78
assign	M_265 = ~|rl_a75_t4 ;	// line#=../rle.cpp:77,78
assign	M_266 = ~|rl_a76_t4 ;	// line#=../rle.cpp:77,78
assign	M_267 = ~|rl_a77_t4 ;	// line#=../rle.cpp:77,78
assign	M_268 = ~|rl_a78_t4 ;	// line#=../rle.cpp:77,78
assign	M_269 = ~|rl_a79_t4 ;	// line#=../rle.cpp:77,78
always @ ( M_269 or M_268 or M_267 or M_266 or M_265 or M_264 or M_263 or M_262 or 
	M_261 or M_260 or M_259 or M_258 or M_257 or M_256 or M_255 or M_254 or 
	decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot [3:0] )
	4'h0 :
		RG_M_14_d10_c4_t = M_254 ;	// line#=../rle.cpp:77,78
	4'h1 :
		RG_M_14_d10_c4_t = M_255 ;	// line#=../rle.cpp:77,78
	4'h2 :
		RG_M_14_d10_c4_t = M_256 ;	// line#=../rle.cpp:77,78
	4'h3 :
		RG_M_14_d10_c4_t = M_257 ;	// line#=../rle.cpp:77,78
	4'h4 :
		RG_M_14_d10_c4_t = M_258 ;	// line#=../rle.cpp:77,78
	4'h5 :
		RG_M_14_d10_c4_t = M_259 ;	// line#=../rle.cpp:77,78
	4'h6 :
		RG_M_14_d10_c4_t = M_260 ;	// line#=../rle.cpp:77,78
	4'h7 :
		RG_M_14_d10_c4_t = M_261 ;	// line#=../rle.cpp:77,78
	4'h8 :
		RG_M_14_d10_c4_t = M_262 ;	// line#=../rle.cpp:77,78
	4'h9 :
		RG_M_14_d10_c4_t = M_263 ;	// line#=../rle.cpp:77,78
	4'ha :
		RG_M_14_d10_c4_t = M_264 ;	// line#=../rle.cpp:77,78
	4'hb :
		RG_M_14_d10_c4_t = M_265 ;	// line#=../rle.cpp:77,78
	4'hc :
		RG_M_14_d10_c4_t = M_266 ;	// line#=../rle.cpp:77,78
	4'hd :
		RG_M_14_d10_c4_t = M_267 ;	// line#=../rle.cpp:77,78
	4'he :
		RG_M_14_d10_c4_t = M_268 ;	// line#=../rle.cpp:77,78
	4'hf :
		RG_M_14_d10_c4_t = M_269 ;	// line#=../rle.cpp:77,78
	default :
		RG_M_14_d10_c4_t = 1'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_M_14_d10_c4 <= RG_M_14_d10_c4_t ;	// line#=../rle.cpp:77,78
assign	M_270 = ~|rl_a80_t4 ;	// line#=../rle.cpp:77,78
assign	M_271 = ~|rl_a81_t4 ;	// line#=../rle.cpp:77,78
assign	M_272 = ~|rl_a82_t4 ;	// line#=../rle.cpp:77,78
assign	M_273 = ~|rl_a83_t4 ;	// line#=../rle.cpp:77,78
assign	M_274 = ~|rl_a84_t4 ;	// line#=../rle.cpp:77,78
assign	M_275 = ~|rl_a85_t4 ;	// line#=../rle.cpp:77,78
assign	M_276 = ~|rl_a86_t4 ;	// line#=../rle.cpp:77,78
assign	M_277 = ~|rl_a87_t4 ;	// line#=../rle.cpp:77,78
assign	M_278 = ~|rl_a88_t4 ;	// line#=../rle.cpp:77,78
assign	M_279 = ~|rl_a89_t4 ;	// line#=../rle.cpp:77,78
assign	M_280 = ~|rl_a90_t4 ;	// line#=../rle.cpp:77,78
assign	M_281 = ~|rl_a91_t4 ;	// line#=../rle.cpp:77,78
assign	M_282 = ~|rl_a92_t4 ;	// line#=../rle.cpp:77,78
assign	M_283 = ~|rl_a93_t4 ;	// line#=../rle.cpp:77,78
assign	M_284 = ~|rl_a94_t4 ;	// line#=../rle.cpp:77,78
assign	M_285 = ~|rl_a95_t4 ;	// line#=../rle.cpp:77,78
always @ ( M_285 or M_284 or M_283 or M_282 or M_281 or M_280 or M_279 or M_278 or 
	M_277 or M_276 or M_275 or M_274 or M_273 or M_272 or M_271 or M_270 or 
	decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot [3:0] )
	4'h0 :
		RG_M_14_d10_c5_t = M_270 ;	// line#=../rle.cpp:77,78
	4'h1 :
		RG_M_14_d10_c5_t = M_271 ;	// line#=../rle.cpp:77,78
	4'h2 :
		RG_M_14_d10_c5_t = M_272 ;	// line#=../rle.cpp:77,78
	4'h3 :
		RG_M_14_d10_c5_t = M_273 ;	// line#=../rle.cpp:77,78
	4'h4 :
		RG_M_14_d10_c5_t = M_274 ;	// line#=../rle.cpp:77,78
	4'h5 :
		RG_M_14_d10_c5_t = M_275 ;	// line#=../rle.cpp:77,78
	4'h6 :
		RG_M_14_d10_c5_t = M_276 ;	// line#=../rle.cpp:77,78
	4'h7 :
		RG_M_14_d10_c5_t = M_277 ;	// line#=../rle.cpp:77,78
	4'h8 :
		RG_M_14_d10_c5_t = M_278 ;	// line#=../rle.cpp:77,78
	4'h9 :
		RG_M_14_d10_c5_t = M_279 ;	// line#=../rle.cpp:77,78
	4'ha :
		RG_M_14_d10_c5_t = M_280 ;	// line#=../rle.cpp:77,78
	4'hb :
		RG_M_14_d10_c5_t = M_281 ;	// line#=../rle.cpp:77,78
	4'hc :
		RG_M_14_d10_c5_t = M_282 ;	// line#=../rle.cpp:77,78
	4'hd :
		RG_M_14_d10_c5_t = M_283 ;	// line#=../rle.cpp:77,78
	4'he :
		RG_M_14_d10_c5_t = M_284 ;	// line#=../rle.cpp:77,78
	4'hf :
		RG_M_14_d10_c5_t = M_285 ;	// line#=../rle.cpp:77,78
	default :
		RG_M_14_d10_c5_t = 1'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_M_14_d10_c5 <= RG_M_14_d10_c5_t ;	// line#=../rle.cpp:77,78
assign	M_286 = ~|rl_a96_t4 ;	// line#=../rle.cpp:77,78
assign	M_287 = ~|rl_a97_t4 ;	// line#=../rle.cpp:77,78
assign	M_288 = ~|rl_a98_t4 ;	// line#=../rle.cpp:77,78
assign	M_289 = ~|rl_a99_t4 ;	// line#=../rle.cpp:77,78
assign	M_290 = ~|rl_a100_t4 ;	// line#=../rle.cpp:77,78
assign	M_291 = ~|rl_a101_t4 ;	// line#=../rle.cpp:77,78
assign	M_292 = ~|rl_a102_t4 ;	// line#=../rle.cpp:77,78
assign	M_293 = ~|rl_a103_t4 ;	// line#=../rle.cpp:77,78
assign	M_294 = ~|rl_a104_t4 ;	// line#=../rle.cpp:77,78
assign	M_295 = ~|rl_a105_t4 ;	// line#=../rle.cpp:77,78
assign	M_296 = ~|rl_a106_t4 ;	// line#=../rle.cpp:77,78
assign	M_297 = ~|rl_a107_t4 ;	// line#=../rle.cpp:77,78
assign	M_298 = ~|rl_a108_t4 ;	// line#=../rle.cpp:77,78
assign	M_299 = ~|rl_a109_t4 ;	// line#=../rle.cpp:77,78
assign	M_300 = ~|rl_a110_t4 ;	// line#=../rle.cpp:77,78
assign	M_301 = ~|rl_a111_t4 ;	// line#=../rle.cpp:77,78
always @ ( M_301 or M_300 or M_299 or M_298 or M_297 or M_296 or M_295 or M_294 or 
	M_293 or M_292 or M_291 or M_290 or M_289 or M_288 or M_287 or M_286 or 
	decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot [3:0] )
	4'h0 :
		RG_M_14_d10_c6_t = M_286 ;	// line#=../rle.cpp:77,78
	4'h1 :
		RG_M_14_d10_c6_t = M_287 ;	// line#=../rle.cpp:77,78
	4'h2 :
		RG_M_14_d10_c6_t = M_288 ;	// line#=../rle.cpp:77,78
	4'h3 :
		RG_M_14_d10_c6_t = M_289 ;	// line#=../rle.cpp:77,78
	4'h4 :
		RG_M_14_d10_c6_t = M_290 ;	// line#=../rle.cpp:77,78
	4'h5 :
		RG_M_14_d10_c6_t = M_291 ;	// line#=../rle.cpp:77,78
	4'h6 :
		RG_M_14_d10_c6_t = M_292 ;	// line#=../rle.cpp:77,78
	4'h7 :
		RG_M_14_d10_c6_t = M_293 ;	// line#=../rle.cpp:77,78
	4'h8 :
		RG_M_14_d10_c6_t = M_294 ;	// line#=../rle.cpp:77,78
	4'h9 :
		RG_M_14_d10_c6_t = M_295 ;	// line#=../rle.cpp:77,78
	4'ha :
		RG_M_14_d10_c6_t = M_296 ;	// line#=../rle.cpp:77,78
	4'hb :
		RG_M_14_d10_c6_t = M_297 ;	// line#=../rle.cpp:77,78
	4'hc :
		RG_M_14_d10_c6_t = M_298 ;	// line#=../rle.cpp:77,78
	4'hd :
		RG_M_14_d10_c6_t = M_299 ;	// line#=../rle.cpp:77,78
	4'he :
		RG_M_14_d10_c6_t = M_300 ;	// line#=../rle.cpp:77,78
	4'hf :
		RG_M_14_d10_c6_t = M_301 ;	// line#=../rle.cpp:77,78
	default :
		RG_M_14_d10_c6_t = 1'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_M_14_d10_c6 <= RG_M_14_d10_c6_t ;	// line#=../rle.cpp:77,78
assign	M_302 = ~|rl_a112_t4 ;	// line#=../rle.cpp:77,78
assign	M_303 = ~|rl_a113_t4 ;	// line#=../rle.cpp:77,78
assign	M_304 = ~|rl_a114_t4 ;	// line#=../rle.cpp:77,78
assign	M_305 = ~|rl_a115_t4 ;	// line#=../rle.cpp:77,78
assign	M_306 = ~|rl_a116_t4 ;	// line#=../rle.cpp:77,78
assign	M_307 = ~|rl_a117_t4 ;	// line#=../rle.cpp:77,78
assign	M_308 = ~|rl_a118_t4 ;	// line#=../rle.cpp:77,78
assign	M_309 = ~|rl_a119_t4 ;	// line#=../rle.cpp:77,78
assign	M_310 = ~|rl_a120_t4 ;	// line#=../rle.cpp:77,78
assign	M_311 = ~|rl_a121_t4 ;	// line#=../rle.cpp:77,78
assign	M_312 = ~|rl_a122_t4 ;	// line#=../rle.cpp:77,78
assign	M_313 = ~|rl_a123_t4 ;	// line#=../rle.cpp:77,78
assign	M_314 = ~|rl_a124_t4 ;	// line#=../rle.cpp:77,78
assign	M_315 = ~|rl_a125_t4 ;	// line#=../rle.cpp:77,78
assign	M_316 = ~|rl_a126_t4 ;	// line#=../rle.cpp:77,78
assign	M_317 = ~|rl_a127_t4 ;	// line#=../rle.cpp:77,78
always @ ( M_317 or M_316 or M_315 or M_314 or M_313 or M_312 or M_311 or M_310 or 
	M_309 or M_308 or M_307 or M_306 or M_305 or M_304 or M_303 or M_302 or 
	decr8u_71ot )	// line#=../rle.cpp:77,78
	case ( decr8u_71ot [3:0] )
	4'h0 :
		RG_M_14_d10_c7_t = M_302 ;	// line#=../rle.cpp:77,78
	4'h1 :
		RG_M_14_d10_c7_t = M_303 ;	// line#=../rle.cpp:77,78
	4'h2 :
		RG_M_14_d10_c7_t = M_304 ;	// line#=../rle.cpp:77,78
	4'h3 :
		RG_M_14_d10_c7_t = M_305 ;	// line#=../rle.cpp:77,78
	4'h4 :
		RG_M_14_d10_c7_t = M_306 ;	// line#=../rle.cpp:77,78
	4'h5 :
		RG_M_14_d10_c7_t = M_307 ;	// line#=../rle.cpp:77,78
	4'h6 :
		RG_M_14_d10_c7_t = M_308 ;	// line#=../rle.cpp:77,78
	4'h7 :
		RG_M_14_d10_c7_t = M_309 ;	// line#=../rle.cpp:77,78
	4'h8 :
		RG_M_14_d10_c7_t = M_310 ;	// line#=../rle.cpp:77,78
	4'h9 :
		RG_M_14_d10_c7_t = M_311 ;	// line#=../rle.cpp:77,78
	4'ha :
		RG_M_14_d10_c7_t = M_312 ;	// line#=../rle.cpp:77,78
	4'hb :
		RG_M_14_d10_c7_t = M_313 ;	// line#=../rle.cpp:77,78
	4'hc :
		RG_M_14_d10_c7_t = M_314 ;	// line#=../rle.cpp:77,78
	4'hd :
		RG_M_14_d10_c7_t = M_315 ;	// line#=../rle.cpp:77,78
	4'he :
		RG_M_14_d10_c7_t = M_316 ;	// line#=../rle.cpp:77,78
	4'hf :
		RG_M_14_d10_c7_t = M_317 ;	// line#=../rle.cpp:77,78
	default :
		RG_M_14_d10_c7_t = 1'hx ;
	endcase
always @ ( posedge clk )	// line#=../rle.cpp:77,78
	RG_M_14_d10_c7 <= RG_M_14_d10_c7_t ;	// line#=../rle.cpp:77,78
always @ ( RG_M_14_d10_c7 or RG_M_14_d10_c6 or RG_M_14_d10_c5 or RG_M_14_d10_c4 or 
	RG_M_14_d10_c3 or RG_M_14_d10_c2 or RG_M_14_d10_c1 or RG_M_14_d10_c0 or 
	RG_323 )
	case ( RG_323 [6:4] )
	3'h0 :
		M_14_t128 = RG_M_14_d10_c0 ;
	3'h1 :
		M_14_t128 = RG_M_14_d10_c1 ;
	3'h2 :
		M_14_t128 = RG_M_14_d10_c2 ;
	3'h3 :
		M_14_t128 = RG_M_14_d10_c3 ;
	3'h4 :
		M_14_t128 = RG_M_14_d10_c4 ;
	3'h5 :
		M_14_t128 = RG_M_14_d10_c5 ;
	3'h6 :
		M_14_t128 = RG_M_14_d10_c6 ;
	3'h7 :
		M_14_t128 = RG_M_14_d10_c7 ;
	default :
		M_14_t128 = 1'hx ;
	endcase
always @ ( RG_rl_127 or RG_rl_126 or RG_rl_125 or RG_rl_124 or RG_rl_123 or RG_rl_122 or 
	RG_rl_121 or RG_rl_120 or RG_rl_119 or RG_rl_118 or RG_rl_117 or RG_rl_116 or 
	RG_rl_115 or RG_rl_114 or RG_rl_113 or RG_rl_112 or RG_rl_111 or RG_rl_110 or 
	RG_rl_109 or RG_rl_108 or RG_rl_107 or RG_rl_106 or RG_rl_105 or RG_rl_104 or 
	RG_rl_103 or RG_rl_102 or RG_rl_101 or RG_rl_100 or RG_rl_99 or RG_rl_98 or 
	RG_rl_97 or RG_rl_96 or RG_rl_95 or RG_rl_94 or RG_rl_93 or RG_rl_92 or 
	RG_rl_91 or RG_rl_90 or RG_rl_89 or RG_rl_88 or RG_rl_87 or RG_rl_86 or 
	RG_rl_85 or RG_rl_84 or RG_rl_83 or RG_rl_82 or RG_rl_81 or RG_rl_80 or 
	RG_rl_79 or RG_rl_78 or RG_rl_77 or RG_rl_76 or RG_rl_75 or RG_rl_74 or 
	RG_rl_73 or RG_rl_72 or RG_rl_71 or RG_rl_70 or RG_rl_69 or RG_rl_68 or 
	RG_rl_67 or RG_rl_66 or RG_rl_65 or RG_rl_64 or RG_rl_63 or RG_rl_62 or 
	RG_rl_61 or RG_rl_60 or RG_rl_59 or RG_rl_58 or RG_rl_57 or RG_rl_56 or 
	RG_rl_55 or RG_rl_54 or RG_rl_53 or RG_rl_52 or RG_rl_51 or RG_rl_50 or 
	RG_rl_49 or RG_rl_48 or RG_rl_47 or RG_rl_46 or RG_rl_45 or RG_rl_44 or 
	RG_rl_43 or RG_rl_42 or RG_rl_41 or RG_rl_40 or RG_rl_39 or RG_rl_38 or 
	RG_rl_37 or RG_rl_36 or RG_rl_35 or RG_rl_34 or RG_rl_33 or RG_rl_32 or 
	RG_rl_31 or RG_rl_30 or RG_rl_29 or RG_rl_28 or RG_rl_27 or RG_rl_26 or 
	RG_rl_25 or RG_rl_24 or RG_rl_23 or RG_rl_22 or RG_rl_21 or RG_rl_20 or 
	RG_rl_19 or RG_rl_18 or RG_rl_17 or RG_rl_16 or RG_rl_15 or RG_rl_14 or 
	RG_rl_13 or RG_rl_12 or RG_rl_11 or RG_rl_10 or RG_rl_9 or RG_rl_8 or RG_rl_7 or 
	RG_rl_6 or RG_rl_5 or RG_rl_4 or RG_rl_3 or RG_rl_2 or RG_rl_1 or RG_rl or 
	sub8u_71ot )	// line#=../rle.cpp:83,84
	case ( sub8u_71ot )
	7'h00 :
		M_15_t128 = ~|{ RG_rl [8:4] , ~RG_rl [3:0] } ;	// line#=../rle.cpp:83,84
	7'h01 :
		M_15_t128 = ~|{ RG_rl_1 [8:4] , ~RG_rl_1 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h02 :
		M_15_t128 = ~|{ RG_rl_2 [8:4] , ~RG_rl_2 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h03 :
		M_15_t128 = ~|{ RG_rl_3 [8:4] , ~RG_rl_3 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h04 :
		M_15_t128 = ~|{ RG_rl_4 [8:4] , ~RG_rl_4 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h05 :
		M_15_t128 = ~|{ RG_rl_5 [8:4] , ~RG_rl_5 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h06 :
		M_15_t128 = ~|{ RG_rl_6 [8:4] , ~RG_rl_6 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h07 :
		M_15_t128 = ~|{ RG_rl_7 [8:4] , ~RG_rl_7 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h08 :
		M_15_t128 = ~|{ RG_rl_8 [8:4] , ~RG_rl_8 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h09 :
		M_15_t128 = ~|{ RG_rl_9 [8:4] , ~RG_rl_9 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0a :
		M_15_t128 = ~|{ RG_rl_10 [8:4] , ~RG_rl_10 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0b :
		M_15_t128 = ~|{ RG_rl_11 [8:4] , ~RG_rl_11 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0c :
		M_15_t128 = ~|{ RG_rl_12 [8:4] , ~RG_rl_12 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0d :
		M_15_t128 = ~|{ RG_rl_13 [8:4] , ~RG_rl_13 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0e :
		M_15_t128 = ~|{ RG_rl_14 [8:4] , ~RG_rl_14 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h0f :
		M_15_t128 = ~|{ RG_rl_15 [8:4] , ~RG_rl_15 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h10 :
		M_15_t128 = ~|{ RG_rl_16 [8:4] , ~RG_rl_16 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h11 :
		M_15_t128 = ~|{ RG_rl_17 [8:4] , ~RG_rl_17 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h12 :
		M_15_t128 = ~|{ RG_rl_18 [8:4] , ~RG_rl_18 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h13 :
		M_15_t128 = ~|{ RG_rl_19 [8:4] , ~RG_rl_19 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h14 :
		M_15_t128 = ~|{ RG_rl_20 [8:4] , ~RG_rl_20 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h15 :
		M_15_t128 = ~|{ RG_rl_21 [8:4] , ~RG_rl_21 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h16 :
		M_15_t128 = ~|{ RG_rl_22 [8:4] , ~RG_rl_22 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h17 :
		M_15_t128 = ~|{ RG_rl_23 [8:4] , ~RG_rl_23 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h18 :
		M_15_t128 = ~|{ RG_rl_24 [8:4] , ~RG_rl_24 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h19 :
		M_15_t128 = ~|{ RG_rl_25 [8:4] , ~RG_rl_25 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1a :
		M_15_t128 = ~|{ RG_rl_26 [8:4] , ~RG_rl_26 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1b :
		M_15_t128 = ~|{ RG_rl_27 [8:4] , ~RG_rl_27 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1c :
		M_15_t128 = ~|{ RG_rl_28 [8:4] , ~RG_rl_28 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1d :
		M_15_t128 = ~|{ RG_rl_29 [8:4] , ~RG_rl_29 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1e :
		M_15_t128 = ~|{ RG_rl_30 [8:4] , ~RG_rl_30 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h1f :
		M_15_t128 = ~|{ RG_rl_31 [8:4] , ~RG_rl_31 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h20 :
		M_15_t128 = ~|{ RG_rl_32 [8:4] , ~RG_rl_32 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h21 :
		M_15_t128 = ~|{ RG_rl_33 [8:4] , ~RG_rl_33 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h22 :
		M_15_t128 = ~|{ RG_rl_34 [8:4] , ~RG_rl_34 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h23 :
		M_15_t128 = ~|{ RG_rl_35 [8:4] , ~RG_rl_35 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h24 :
		M_15_t128 = ~|{ RG_rl_36 [8:4] , ~RG_rl_36 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h25 :
		M_15_t128 = ~|{ RG_rl_37 [8:4] , ~RG_rl_37 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h26 :
		M_15_t128 = ~|{ RG_rl_38 [8:4] , ~RG_rl_38 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h27 :
		M_15_t128 = ~|{ RG_rl_39 [8:4] , ~RG_rl_39 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h28 :
		M_15_t128 = ~|{ RG_rl_40 [8:4] , ~RG_rl_40 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h29 :
		M_15_t128 = ~|{ RG_rl_41 [8:4] , ~RG_rl_41 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2a :
		M_15_t128 = ~|{ RG_rl_42 [8:4] , ~RG_rl_42 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2b :
		M_15_t128 = ~|{ RG_rl_43 [8:4] , ~RG_rl_43 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2c :
		M_15_t128 = ~|{ RG_rl_44 [8:4] , ~RG_rl_44 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2d :
		M_15_t128 = ~|{ RG_rl_45 [8:4] , ~RG_rl_45 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2e :
		M_15_t128 = ~|{ RG_rl_46 [8:4] , ~RG_rl_46 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h2f :
		M_15_t128 = ~|{ RG_rl_47 [8:4] , ~RG_rl_47 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h30 :
		M_15_t128 = ~|{ RG_rl_48 [8:4] , ~RG_rl_48 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h31 :
		M_15_t128 = ~|{ RG_rl_49 [8:4] , ~RG_rl_49 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h32 :
		M_15_t128 = ~|{ RG_rl_50 [8:4] , ~RG_rl_50 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h33 :
		M_15_t128 = ~|{ RG_rl_51 [8:4] , ~RG_rl_51 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h34 :
		M_15_t128 = ~|{ RG_rl_52 [8:4] , ~RG_rl_52 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h35 :
		M_15_t128 = ~|{ RG_rl_53 [8:4] , ~RG_rl_53 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h36 :
		M_15_t128 = ~|{ RG_rl_54 [8:4] , ~RG_rl_54 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h37 :
		M_15_t128 = ~|{ RG_rl_55 [8:4] , ~RG_rl_55 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h38 :
		M_15_t128 = ~|{ RG_rl_56 [8:4] , ~RG_rl_56 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h39 :
		M_15_t128 = ~|{ RG_rl_57 [8:4] , ~RG_rl_57 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3a :
		M_15_t128 = ~|{ RG_rl_58 [8:4] , ~RG_rl_58 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3b :
		M_15_t128 = ~|{ RG_rl_59 [8:4] , ~RG_rl_59 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3c :
		M_15_t128 = ~|{ RG_rl_60 [8:4] , ~RG_rl_60 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3d :
		M_15_t128 = ~|{ RG_rl_61 [8:4] , ~RG_rl_61 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3e :
		M_15_t128 = ~|{ RG_rl_62 [8:4] , ~RG_rl_62 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h3f :
		M_15_t128 = ~|{ RG_rl_63 [8:4] , ~RG_rl_63 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h40 :
		M_15_t128 = ~|{ RG_rl_64 [8:4] , ~RG_rl_64 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h41 :
		M_15_t128 = ~|{ RG_rl_65 [8:4] , ~RG_rl_65 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h42 :
		M_15_t128 = ~|{ RG_rl_66 [8:4] , ~RG_rl_66 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h43 :
		M_15_t128 = ~|{ RG_rl_67 [8:4] , ~RG_rl_67 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h44 :
		M_15_t128 = ~|{ RG_rl_68 [8:4] , ~RG_rl_68 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h45 :
		M_15_t128 = ~|{ RG_rl_69 [8:4] , ~RG_rl_69 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h46 :
		M_15_t128 = ~|{ RG_rl_70 [8:4] , ~RG_rl_70 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h47 :
		M_15_t128 = ~|{ RG_rl_71 [8:4] , ~RG_rl_71 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h48 :
		M_15_t128 = ~|{ RG_rl_72 [8:4] , ~RG_rl_72 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h49 :
		M_15_t128 = ~|{ RG_rl_73 [8:4] , ~RG_rl_73 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4a :
		M_15_t128 = ~|{ RG_rl_74 [8:4] , ~RG_rl_74 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4b :
		M_15_t128 = ~|{ RG_rl_75 [8:4] , ~RG_rl_75 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4c :
		M_15_t128 = ~|{ RG_rl_76 [8:4] , ~RG_rl_76 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4d :
		M_15_t128 = ~|{ RG_rl_77 [8:4] , ~RG_rl_77 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4e :
		M_15_t128 = ~|{ RG_rl_78 [8:4] , ~RG_rl_78 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h4f :
		M_15_t128 = ~|{ RG_rl_79 [8:4] , ~RG_rl_79 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h50 :
		M_15_t128 = ~|{ RG_rl_80 [8:4] , ~RG_rl_80 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h51 :
		M_15_t128 = ~|{ RG_rl_81 [8:4] , ~RG_rl_81 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h52 :
		M_15_t128 = ~|{ RG_rl_82 [8:4] , ~RG_rl_82 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h53 :
		M_15_t128 = ~|{ RG_rl_83 [8:4] , ~RG_rl_83 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h54 :
		M_15_t128 = ~|{ RG_rl_84 [8:4] , ~RG_rl_84 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h55 :
		M_15_t128 = ~|{ RG_rl_85 [8:4] , ~RG_rl_85 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h56 :
		M_15_t128 = ~|{ RG_rl_86 [8:4] , ~RG_rl_86 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h57 :
		M_15_t128 = ~|{ RG_rl_87 [8:4] , ~RG_rl_87 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h58 :
		M_15_t128 = ~|{ RG_rl_88 [8:4] , ~RG_rl_88 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h59 :
		M_15_t128 = ~|{ RG_rl_89 [8:4] , ~RG_rl_89 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5a :
		M_15_t128 = ~|{ RG_rl_90 [8:4] , ~RG_rl_90 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5b :
		M_15_t128 = ~|{ RG_rl_91 [8:4] , ~RG_rl_91 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5c :
		M_15_t128 = ~|{ RG_rl_92 [8:4] , ~RG_rl_92 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5d :
		M_15_t128 = ~|{ RG_rl_93 [8:4] , ~RG_rl_93 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5e :
		M_15_t128 = ~|{ RG_rl_94 [8:4] , ~RG_rl_94 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h5f :
		M_15_t128 = ~|{ RG_rl_95 [8:4] , ~RG_rl_95 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h60 :
		M_15_t128 = ~|{ RG_rl_96 [8:4] , ~RG_rl_96 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h61 :
		M_15_t128 = ~|{ RG_rl_97 [8:4] , ~RG_rl_97 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h62 :
		M_15_t128 = ~|{ RG_rl_98 [8:4] , ~RG_rl_98 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h63 :
		M_15_t128 = ~|{ RG_rl_99 [8:4] , ~RG_rl_99 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h64 :
		M_15_t128 = ~|{ RG_rl_100 [8:4] , ~RG_rl_100 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h65 :
		M_15_t128 = ~|{ RG_rl_101 [8:4] , ~RG_rl_101 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h66 :
		M_15_t128 = ~|{ RG_rl_102 [8:4] , ~RG_rl_102 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h67 :
		M_15_t128 = ~|{ RG_rl_103 [8:4] , ~RG_rl_103 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h68 :
		M_15_t128 = ~|{ RG_rl_104 [8:4] , ~RG_rl_104 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h69 :
		M_15_t128 = ~|{ RG_rl_105 [8:4] , ~RG_rl_105 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6a :
		M_15_t128 = ~|{ RG_rl_106 [8:4] , ~RG_rl_106 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6b :
		M_15_t128 = ~|{ RG_rl_107 [8:4] , ~RG_rl_107 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6c :
		M_15_t128 = ~|{ RG_rl_108 [8:4] , ~RG_rl_108 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6d :
		M_15_t128 = ~|{ RG_rl_109 [8:4] , ~RG_rl_109 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6e :
		M_15_t128 = ~|{ RG_rl_110 [8:4] , ~RG_rl_110 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h6f :
		M_15_t128 = ~|{ RG_rl_111 [8:4] , ~RG_rl_111 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h70 :
		M_15_t128 = ~|{ RG_rl_112 [8:4] , ~RG_rl_112 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h71 :
		M_15_t128 = ~|{ RG_rl_113 [8:4] , ~RG_rl_113 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h72 :
		M_15_t128 = ~|{ RG_rl_114 [8:4] , ~RG_rl_114 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h73 :
		M_15_t128 = ~|{ RG_rl_115 [8:4] , ~RG_rl_115 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h74 :
		M_15_t128 = ~|{ RG_rl_116 [8:4] , ~RG_rl_116 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h75 :
		M_15_t128 = ~|{ RG_rl_117 [8:4] , ~RG_rl_117 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h76 :
		M_15_t128 = ~|{ RG_rl_118 [8:4] , ~RG_rl_118 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h77 :
		M_15_t128 = ~|{ RG_rl_119 [8:4] , ~RG_rl_119 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h78 :
		M_15_t128 = ~|{ RG_rl_120 [8:4] , ~RG_rl_120 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h79 :
		M_15_t128 = ~|{ RG_rl_121 [8:4] , ~RG_rl_121 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7a :
		M_15_t128 = ~|{ RG_rl_122 [8:4] , ~RG_rl_122 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7b :
		M_15_t128 = ~|{ RG_rl_123 [8:4] , ~RG_rl_123 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7c :
		M_15_t128 = ~|{ RG_rl_124 [8:4] , ~RG_rl_124 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7d :
		M_15_t128 = ~|{ RG_rl_125 [8:4] , ~RG_rl_125 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7e :
		M_15_t128 = ~|{ RG_rl_126 [8:4] , ~RG_rl_126 [3:0] } ;	// line#=../rle.cpp:83,84
	7'h7f :
		M_15_t128 = ~|{ RG_rl_127 [8:4] , ~RG_rl_127 [3:0] } ;	// line#=../rle.cpp:83,84
	default :
		M_15_t128 = 1'hx ;
	endcase
jpeg_MEMB9W64 zz ( .RA1(zz_RA1) ,.RD1(zz_RD1) ,.RCLK1(clk) ,.WA2(RG_k_01[5:0]) ,
	.WD2(zz_WD2) ,.WE2(zz_WE2) ,.WCLK2(clk) );	// line#=../rle.h:65
assign	sub12s_91i1 = zz_RD1 ;	// line#=../rle.cpp:52,53
assign	sub12s_91i2 = RG_previous_dc_rl ;	// line#=../rle.cpp:52
assign	lop8u_11i1 = RG_k_01 [5:0] ;	// line#=../rle.cpp:109,110
assign	lop8u_11i2 = 6'h24 ;	// line#=../rle.cpp:109,110
assign	incr4s1i1 = RG_j ;	// line#=../rle.cpp:34
assign	incr8u2i1 = incr8u1ot ;	// line#=../rle.cpp:68,69
assign	incr8u4i1 = incr8u1ot ;	// line#=../rle.cpp:79,80
assign	incr32s3i1 = RG_i_j_01 ;	// line#=../rle.cpp:74
assign	decr8u_71i1 = len1_t3 [6:0] ;	// line#=../rle.cpp:77,78
assign	sub8u_71i1 = RG_len [6:0] ;	// line#=../rle.cpp:83,84
assign	sub8u_71i2 = 3'h4 ;	// line#=../rle.cpp:83,84
assign	sub8u_7_11i1 = RG_len [6:0] ;	// line#=../rle.cpp:83,84
assign	sub8u_7_11i2 = 2'h3 ;	// line#=../rle.cpp:83,84
assign	C_01 = ~|{ ~incr4s1ot [3] , incr4s1ot [2:0] } ;	// line#=../rle.cpp:34,35
assign	U_01 = ( ST1_02d & C_01 ) ;	// line#=../rle.cpp:35
assign	U_05 = ( ST1_03d & lop8u_11ot ) ;	// line#=../rle.cpp:109,110
assign	U_06 = ( ST1_03d & ( ~lop8u_11ot ) ) ;	// line#=../rle.cpp:109,110
assign	U_07 = ( U_05 & M_175 ) ;	// line#=../rle.cpp:111
assign	U_08 = ( U_05 & M_173 ) ;	// line#=../rle.cpp:111
assign	U_09 = ( U_05 & M_177 ) ;	// line#=../rle.cpp:111
assign	U_10 = ( U_05 & M_183 ) ;	// line#=../rle.cpp:111
assign	U_11 = ( U_05 & M_181 ) ;	// line#=../rle.cpp:111
assign	U_12 = ( U_05 & M_185 ) ;	// line#=../rle.cpp:111
assign	U_13 = ( U_05 & M_187 ) ;	// line#=../rle.cpp:111
assign	U_14 = ( U_05 & M_179 ) ;	// line#=../rle.cpp:111
assign	C_02 = ( ( ~|RG_i_k_01 ) & M_189 ) ;	// line#=../rle.cpp:112,113
assign	U_79 = ( U_05 & C_02 ) ;	// line#=../rle.cpp:112,113
assign	U_80 = ( U_05 & ( ~C_02 ) ) ;	// line#=../rle.cpp:112,113
assign	U_81 = ( U_80 & CT_12 ) ;	// line#=../rle.cpp:117,118
assign	U_82 = ( U_80 & ( ~CT_12 ) ) ;	// line#=../rle.cpp:117,118
assign	U_83 = ( U_82 & ( ~FF_d_01 ) ) ;	// line#=../rle.cpp:122,123
assign	U_84 = ( U_82 & FF_d_01 ) ;	// line#=../rle.cpp:122,123
assign	U_87 = ( ST1_04d & ( ~RG_k_01 [6] ) ) ;	// line#=../rle.cpp:140,141
assign	U_88 = ( ST1_04d & RG_k_01 [6] ) ;	// line#=../rle.cpp:140,141
assign	M_175 = ~|RG_i_k_01 [2:0] ;	// line#=../rle.cpp:111,140,141,142
assign	U_89 = ( U_87 & M_175 ) ;	// line#=../rle.cpp:140,141,142
assign	M_173 = ~|( RG_i_k_01 [2:0] ^ 3'h1 ) ;	// line#=../rle.cpp:111,140,141,142
assign	U_90 = ( U_87 & M_173 ) ;	// line#=../rle.cpp:140,141,142
assign	M_177 = ~|( RG_i_k_01 [2:0] ^ 3'h2 ) ;	// line#=../rle.cpp:111,140,141,142
assign	U_91 = ( U_87 & M_177 ) ;	// line#=../rle.cpp:140,141,142
assign	M_183 = ~|( RG_i_k_01 [2:0] ^ 3'h3 ) ;	// line#=../rle.cpp:111,140,141,142
assign	U_92 = ( U_87 & M_183 ) ;	// line#=../rle.cpp:140,141,142
assign	M_181 = ~|( RG_i_k_01 [2:0] ^ 3'h4 ) ;	// line#=../rle.cpp:111,140,141,142
assign	U_93 = ( U_87 & M_181 ) ;	// line#=../rle.cpp:140,141,142
assign	M_185 = ~|( RG_i_k_01 [2:0] ^ 3'h5 ) ;	// line#=../rle.cpp:111,140,141,142
assign	U_94 = ( U_87 & M_185 ) ;	// line#=../rle.cpp:140,141,142
assign	M_187 = ~|( RG_i_k_01 [2:0] ^ 3'h6 ) ;	// line#=../rle.cpp:111,140,141,142
assign	U_95 = ( U_87 & M_187 ) ;	// line#=../rle.cpp:140,141,142
assign	M_179 = ~|( RG_i_k_01 [2:0] ^ 3'h7 ) ;	// line#=../rle.cpp:111,140,141,142
assign	U_96 = ( U_87 & M_179 ) ;	// line#=../rle.cpp:140,141,142
assign	M_189 = ~|{ ( RG_i_j_01 [31] & RG_i_j_01 [0] ) , RG_i_j_01 [0] } ;	// line#=../rle.cpp:112,113,140,141,143
										// ,144
assign	C_05 = ( ( ~|{ RG_i_k_01 [31:3] , ~RG_i_k_01 [2:0] } ) & M_189 ) ;	// line#=../rle.cpp:140,141,143,144
assign	U_161 = ( U_87 & C_05 ) ;	// line#=../rle.cpp:143,144
assign	U_162 = ( U_87 & ( ~C_05 ) ) ;	// line#=../rle.cpp:143,144
assign	U_163 = ( U_162 & CT_17 ) ;	// line#=../rle.cpp:148,149
assign	U_164 = ( U_162 & ( ~CT_17 ) ) ;	// line#=../rle.cpp:148,149
assign	U_165 = ( U_164 & ( ~FF_d_01 ) ) ;	// line#=../rle.cpp:153,154
assign	U_166 = ( U_164 & FF_d_01 ) ;	// line#=../rle.cpp:153,154
assign	U_171 = ( ST1_08d & CT_33 ) ;	// line#=../rle.cpp:61,62
assign	U_172 = ( ST1_08d & ( ~CT_33 ) ) ;	// line#=../rle.cpp:61,62
assign	U_173 = ( U_172 & CT_32 ) ;	// line#=../rle.cpp:66,67
assign	U_174 = ( U_172 & ( ~CT_32 ) ) ;	// line#=../rle.cpp:66,67
assign	U_569 = ( ST1_10d & ( ~M_02_t ) ) ;	// line#=../rle.cpp:77,78
assign	U_570 = ( ST1_10d & M_02_t ) ;	// line#=../rle.cpp:77,78
assign	U_571 = ( ST1_11d & M_03_t128 ) ;	// line#=../rle.cpp:83,84
assign	U_572 = ( ST1_11d & ( ~M_03_t128 ) ) ;	// line#=../rle.cpp:83,84
always @ ( TR_12 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h01 :
		RG_rl_t1 = TR_12 ;
	7'h02 :
		RG_rl_t1 = TR_12 ;
	7'h03 :
		RG_rl_t1 = TR_12 ;
	7'h04 :
		RG_rl_t1 = TR_12 ;
	7'h05 :
		RG_rl_t1 = TR_12 ;
	7'h06 :
		RG_rl_t1 = TR_12 ;
	7'h07 :
		RG_rl_t1 = TR_12 ;
	7'h08 :
		RG_rl_t1 = TR_12 ;
	7'h09 :
		RG_rl_t1 = TR_12 ;
	7'h0a :
		RG_rl_t1 = TR_12 ;
	7'h0b :
		RG_rl_t1 = TR_12 ;
	7'h0c :
		RG_rl_t1 = TR_12 ;
	7'h0d :
		RG_rl_t1 = TR_12 ;
	7'h0e :
		RG_rl_t1 = TR_12 ;
	7'h0f :
		RG_rl_t1 = TR_12 ;
	7'h10 :
		RG_rl_t1 = TR_12 ;
	7'h11 :
		RG_rl_t1 = TR_12 ;
	7'h12 :
		RG_rl_t1 = TR_12 ;
	7'h13 :
		RG_rl_t1 = TR_12 ;
	7'h14 :
		RG_rl_t1 = TR_12 ;
	7'h15 :
		RG_rl_t1 = TR_12 ;
	7'h16 :
		RG_rl_t1 = TR_12 ;
	7'h17 :
		RG_rl_t1 = TR_12 ;
	7'h18 :
		RG_rl_t1 = TR_12 ;
	7'h19 :
		RG_rl_t1 = TR_12 ;
	7'h1a :
		RG_rl_t1 = TR_12 ;
	7'h1b :
		RG_rl_t1 = TR_12 ;
	7'h1c :
		RG_rl_t1 = TR_12 ;
	7'h1d :
		RG_rl_t1 = TR_12 ;
	7'h1e :
		RG_rl_t1 = TR_12 ;
	7'h1f :
		RG_rl_t1 = TR_12 ;
	7'h20 :
		RG_rl_t1 = TR_12 ;
	7'h21 :
		RG_rl_t1 = TR_12 ;
	7'h22 :
		RG_rl_t1 = TR_12 ;
	7'h23 :
		RG_rl_t1 = TR_12 ;
	7'h24 :
		RG_rl_t1 = TR_12 ;
	7'h25 :
		RG_rl_t1 = TR_12 ;
	7'h26 :
		RG_rl_t1 = TR_12 ;
	7'h27 :
		RG_rl_t1 = TR_12 ;
	7'h28 :
		RG_rl_t1 = TR_12 ;
	7'h29 :
		RG_rl_t1 = TR_12 ;
	7'h2a :
		RG_rl_t1 = TR_12 ;
	7'h2b :
		RG_rl_t1 = TR_12 ;
	7'h2c :
		RG_rl_t1 = TR_12 ;
	7'h2d :
		RG_rl_t1 = TR_12 ;
	7'h2e :
		RG_rl_t1 = TR_12 ;
	7'h2f :
		RG_rl_t1 = TR_12 ;
	7'h30 :
		RG_rl_t1 = TR_12 ;
	7'h31 :
		RG_rl_t1 = TR_12 ;
	7'h32 :
		RG_rl_t1 = TR_12 ;
	7'h33 :
		RG_rl_t1 = TR_12 ;
	7'h34 :
		RG_rl_t1 = TR_12 ;
	7'h35 :
		RG_rl_t1 = TR_12 ;
	7'h36 :
		RG_rl_t1 = TR_12 ;
	7'h37 :
		RG_rl_t1 = TR_12 ;
	7'h38 :
		RG_rl_t1 = TR_12 ;
	7'h39 :
		RG_rl_t1 = TR_12 ;
	7'h3a :
		RG_rl_t1 = TR_12 ;
	7'h3b :
		RG_rl_t1 = TR_12 ;
	7'h3c :
		RG_rl_t1 = TR_12 ;
	7'h3d :
		RG_rl_t1 = TR_12 ;
	7'h3e :
		RG_rl_t1 = TR_12 ;
	7'h3f :
		RG_rl_t1 = TR_12 ;
	7'h40 :
		RG_rl_t1 = TR_12 ;
	7'h41 :
		RG_rl_t1 = TR_12 ;
	7'h42 :
		RG_rl_t1 = TR_12 ;
	7'h43 :
		RG_rl_t1 = TR_12 ;
	7'h44 :
		RG_rl_t1 = TR_12 ;
	7'h45 :
		RG_rl_t1 = TR_12 ;
	7'h46 :
		RG_rl_t1 = TR_12 ;
	7'h47 :
		RG_rl_t1 = TR_12 ;
	7'h48 :
		RG_rl_t1 = TR_12 ;
	7'h49 :
		RG_rl_t1 = TR_12 ;
	7'h4a :
		RG_rl_t1 = TR_12 ;
	7'h4b :
		RG_rl_t1 = TR_12 ;
	7'h4c :
		RG_rl_t1 = TR_12 ;
	7'h4d :
		RG_rl_t1 = TR_12 ;
	7'h4e :
		RG_rl_t1 = TR_12 ;
	7'h4f :
		RG_rl_t1 = TR_12 ;
	7'h50 :
		RG_rl_t1 = TR_12 ;
	7'h51 :
		RG_rl_t1 = TR_12 ;
	7'h52 :
		RG_rl_t1 = TR_12 ;
	7'h53 :
		RG_rl_t1 = TR_12 ;
	7'h54 :
		RG_rl_t1 = TR_12 ;
	7'h55 :
		RG_rl_t1 = TR_12 ;
	7'h56 :
		RG_rl_t1 = TR_12 ;
	7'h57 :
		RG_rl_t1 = TR_12 ;
	7'h58 :
		RG_rl_t1 = TR_12 ;
	7'h59 :
		RG_rl_t1 = TR_12 ;
	7'h5a :
		RG_rl_t1 = TR_12 ;
	7'h5b :
		RG_rl_t1 = TR_12 ;
	7'h5c :
		RG_rl_t1 = TR_12 ;
	7'h5d :
		RG_rl_t1 = TR_12 ;
	7'h5e :
		RG_rl_t1 = TR_12 ;
	7'h5f :
		RG_rl_t1 = TR_12 ;
	7'h60 :
		RG_rl_t1 = TR_12 ;
	7'h61 :
		RG_rl_t1 = TR_12 ;
	7'h62 :
		RG_rl_t1 = TR_12 ;
	7'h63 :
		RG_rl_t1 = TR_12 ;
	7'h64 :
		RG_rl_t1 = TR_12 ;
	7'h65 :
		RG_rl_t1 = TR_12 ;
	7'h66 :
		RG_rl_t1 = TR_12 ;
	7'h67 :
		RG_rl_t1 = TR_12 ;
	7'h68 :
		RG_rl_t1 = TR_12 ;
	7'h69 :
		RG_rl_t1 = TR_12 ;
	7'h6a :
		RG_rl_t1 = TR_12 ;
	7'h6b :
		RG_rl_t1 = TR_12 ;
	7'h6c :
		RG_rl_t1 = TR_12 ;
	7'h6d :
		RG_rl_t1 = TR_12 ;
	7'h6e :
		RG_rl_t1 = TR_12 ;
	7'h6f :
		RG_rl_t1 = TR_12 ;
	7'h70 :
		RG_rl_t1 = TR_12 ;
	7'h71 :
		RG_rl_t1 = TR_12 ;
	7'h72 :
		RG_rl_t1 = TR_12 ;
	7'h73 :
		RG_rl_t1 = TR_12 ;
	7'h74 :
		RG_rl_t1 = TR_12 ;
	7'h75 :
		RG_rl_t1 = TR_12 ;
	7'h76 :
		RG_rl_t1 = TR_12 ;
	7'h77 :
		RG_rl_t1 = TR_12 ;
	7'h78 :
		RG_rl_t1 = TR_12 ;
	7'h79 :
		RG_rl_t1 = TR_12 ;
	7'h7a :
		RG_rl_t1 = TR_12 ;
	7'h7b :
		RG_rl_t1 = TR_12 ;
	7'h7c :
		RG_rl_t1 = TR_12 ;
	7'h7d :
		RG_rl_t1 = TR_12 ;
	7'h7e :
		RG_rl_t1 = TR_12 ;
	7'h7f :
		RG_rl_t1 = TR_12 ;
	default :
		RG_rl_t1 = 9'hx ;
	endcase
always @ ( RG_rl_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_184 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_t_c1 = ( U_571 & ( ~|sub8u_71ot ) ) ;	// line#=../rle.cpp:85
	RG_rl_t = ( ( { 9{ U_570 } } & RG_rl_184 )
		| ( { 9{ U_569 } } & RG_rl_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_en = ( U_570 | RG_rl_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_en )
		RG_rl <= RG_rl_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_13 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_1_t1 = TR_13 ;
	7'h01 :
		RG_rl_1_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h02 :
		RG_rl_1_t1 = TR_13 ;
	7'h03 :
		RG_rl_1_t1 = TR_13 ;
	7'h04 :
		RG_rl_1_t1 = TR_13 ;
	7'h05 :
		RG_rl_1_t1 = TR_13 ;
	7'h06 :
		RG_rl_1_t1 = TR_13 ;
	7'h07 :
		RG_rl_1_t1 = TR_13 ;
	7'h08 :
		RG_rl_1_t1 = TR_13 ;
	7'h09 :
		RG_rl_1_t1 = TR_13 ;
	7'h0a :
		RG_rl_1_t1 = TR_13 ;
	7'h0b :
		RG_rl_1_t1 = TR_13 ;
	7'h0c :
		RG_rl_1_t1 = TR_13 ;
	7'h0d :
		RG_rl_1_t1 = TR_13 ;
	7'h0e :
		RG_rl_1_t1 = TR_13 ;
	7'h0f :
		RG_rl_1_t1 = TR_13 ;
	7'h10 :
		RG_rl_1_t1 = TR_13 ;
	7'h11 :
		RG_rl_1_t1 = TR_13 ;
	7'h12 :
		RG_rl_1_t1 = TR_13 ;
	7'h13 :
		RG_rl_1_t1 = TR_13 ;
	7'h14 :
		RG_rl_1_t1 = TR_13 ;
	7'h15 :
		RG_rl_1_t1 = TR_13 ;
	7'h16 :
		RG_rl_1_t1 = TR_13 ;
	7'h17 :
		RG_rl_1_t1 = TR_13 ;
	7'h18 :
		RG_rl_1_t1 = TR_13 ;
	7'h19 :
		RG_rl_1_t1 = TR_13 ;
	7'h1a :
		RG_rl_1_t1 = TR_13 ;
	7'h1b :
		RG_rl_1_t1 = TR_13 ;
	7'h1c :
		RG_rl_1_t1 = TR_13 ;
	7'h1d :
		RG_rl_1_t1 = TR_13 ;
	7'h1e :
		RG_rl_1_t1 = TR_13 ;
	7'h1f :
		RG_rl_1_t1 = TR_13 ;
	7'h20 :
		RG_rl_1_t1 = TR_13 ;
	7'h21 :
		RG_rl_1_t1 = TR_13 ;
	7'h22 :
		RG_rl_1_t1 = TR_13 ;
	7'h23 :
		RG_rl_1_t1 = TR_13 ;
	7'h24 :
		RG_rl_1_t1 = TR_13 ;
	7'h25 :
		RG_rl_1_t1 = TR_13 ;
	7'h26 :
		RG_rl_1_t1 = TR_13 ;
	7'h27 :
		RG_rl_1_t1 = TR_13 ;
	7'h28 :
		RG_rl_1_t1 = TR_13 ;
	7'h29 :
		RG_rl_1_t1 = TR_13 ;
	7'h2a :
		RG_rl_1_t1 = TR_13 ;
	7'h2b :
		RG_rl_1_t1 = TR_13 ;
	7'h2c :
		RG_rl_1_t1 = TR_13 ;
	7'h2d :
		RG_rl_1_t1 = TR_13 ;
	7'h2e :
		RG_rl_1_t1 = TR_13 ;
	7'h2f :
		RG_rl_1_t1 = TR_13 ;
	7'h30 :
		RG_rl_1_t1 = TR_13 ;
	7'h31 :
		RG_rl_1_t1 = TR_13 ;
	7'h32 :
		RG_rl_1_t1 = TR_13 ;
	7'h33 :
		RG_rl_1_t1 = TR_13 ;
	7'h34 :
		RG_rl_1_t1 = TR_13 ;
	7'h35 :
		RG_rl_1_t1 = TR_13 ;
	7'h36 :
		RG_rl_1_t1 = TR_13 ;
	7'h37 :
		RG_rl_1_t1 = TR_13 ;
	7'h38 :
		RG_rl_1_t1 = TR_13 ;
	7'h39 :
		RG_rl_1_t1 = TR_13 ;
	7'h3a :
		RG_rl_1_t1 = TR_13 ;
	7'h3b :
		RG_rl_1_t1 = TR_13 ;
	7'h3c :
		RG_rl_1_t1 = TR_13 ;
	7'h3d :
		RG_rl_1_t1 = TR_13 ;
	7'h3e :
		RG_rl_1_t1 = TR_13 ;
	7'h3f :
		RG_rl_1_t1 = TR_13 ;
	7'h40 :
		RG_rl_1_t1 = TR_13 ;
	7'h41 :
		RG_rl_1_t1 = TR_13 ;
	7'h42 :
		RG_rl_1_t1 = TR_13 ;
	7'h43 :
		RG_rl_1_t1 = TR_13 ;
	7'h44 :
		RG_rl_1_t1 = TR_13 ;
	7'h45 :
		RG_rl_1_t1 = TR_13 ;
	7'h46 :
		RG_rl_1_t1 = TR_13 ;
	7'h47 :
		RG_rl_1_t1 = TR_13 ;
	7'h48 :
		RG_rl_1_t1 = TR_13 ;
	7'h49 :
		RG_rl_1_t1 = TR_13 ;
	7'h4a :
		RG_rl_1_t1 = TR_13 ;
	7'h4b :
		RG_rl_1_t1 = TR_13 ;
	7'h4c :
		RG_rl_1_t1 = TR_13 ;
	7'h4d :
		RG_rl_1_t1 = TR_13 ;
	7'h4e :
		RG_rl_1_t1 = TR_13 ;
	7'h4f :
		RG_rl_1_t1 = TR_13 ;
	7'h50 :
		RG_rl_1_t1 = TR_13 ;
	7'h51 :
		RG_rl_1_t1 = TR_13 ;
	7'h52 :
		RG_rl_1_t1 = TR_13 ;
	7'h53 :
		RG_rl_1_t1 = TR_13 ;
	7'h54 :
		RG_rl_1_t1 = TR_13 ;
	7'h55 :
		RG_rl_1_t1 = TR_13 ;
	7'h56 :
		RG_rl_1_t1 = TR_13 ;
	7'h57 :
		RG_rl_1_t1 = TR_13 ;
	7'h58 :
		RG_rl_1_t1 = TR_13 ;
	7'h59 :
		RG_rl_1_t1 = TR_13 ;
	7'h5a :
		RG_rl_1_t1 = TR_13 ;
	7'h5b :
		RG_rl_1_t1 = TR_13 ;
	7'h5c :
		RG_rl_1_t1 = TR_13 ;
	7'h5d :
		RG_rl_1_t1 = TR_13 ;
	7'h5e :
		RG_rl_1_t1 = TR_13 ;
	7'h5f :
		RG_rl_1_t1 = TR_13 ;
	7'h60 :
		RG_rl_1_t1 = TR_13 ;
	7'h61 :
		RG_rl_1_t1 = TR_13 ;
	7'h62 :
		RG_rl_1_t1 = TR_13 ;
	7'h63 :
		RG_rl_1_t1 = TR_13 ;
	7'h64 :
		RG_rl_1_t1 = TR_13 ;
	7'h65 :
		RG_rl_1_t1 = TR_13 ;
	7'h66 :
		RG_rl_1_t1 = TR_13 ;
	7'h67 :
		RG_rl_1_t1 = TR_13 ;
	7'h68 :
		RG_rl_1_t1 = TR_13 ;
	7'h69 :
		RG_rl_1_t1 = TR_13 ;
	7'h6a :
		RG_rl_1_t1 = TR_13 ;
	7'h6b :
		RG_rl_1_t1 = TR_13 ;
	7'h6c :
		RG_rl_1_t1 = TR_13 ;
	7'h6d :
		RG_rl_1_t1 = TR_13 ;
	7'h6e :
		RG_rl_1_t1 = TR_13 ;
	7'h6f :
		RG_rl_1_t1 = TR_13 ;
	7'h70 :
		RG_rl_1_t1 = TR_13 ;
	7'h71 :
		RG_rl_1_t1 = TR_13 ;
	7'h72 :
		RG_rl_1_t1 = TR_13 ;
	7'h73 :
		RG_rl_1_t1 = TR_13 ;
	7'h74 :
		RG_rl_1_t1 = TR_13 ;
	7'h75 :
		RG_rl_1_t1 = TR_13 ;
	7'h76 :
		RG_rl_1_t1 = TR_13 ;
	7'h77 :
		RG_rl_1_t1 = TR_13 ;
	7'h78 :
		RG_rl_1_t1 = TR_13 ;
	7'h79 :
		RG_rl_1_t1 = TR_13 ;
	7'h7a :
		RG_rl_1_t1 = TR_13 ;
	7'h7b :
		RG_rl_1_t1 = TR_13 ;
	7'h7c :
		RG_rl_1_t1 = TR_13 ;
	7'h7d :
		RG_rl_1_t1 = TR_13 ;
	7'h7e :
		RG_rl_1_t1 = TR_13 ;
	7'h7f :
		RG_rl_1_t1 = TR_13 ;
	default :
		RG_rl_1_t1 = 9'hx ;
	endcase
always @ ( RG_rl_1_t1 or U_569 or sub8u_71ot or U_571 or RG_previous_dc_rl or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_1_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h01 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_1_t = ( ( { 9{ U_570 } } & RG_previous_dc_rl )
		| ( { 9{ U_569 } } & RG_rl_1_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_1_en = ( U_570 | RG_rl_1_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_1_en )
		RG_rl_1 <= RG_rl_1_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_14 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_2_t1 = TR_14 ;
	7'h01 :
		RG_rl_2_t1 = TR_14 ;
	7'h02 :
		RG_rl_2_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h03 :
		RG_rl_2_t1 = TR_14 ;
	7'h04 :
		RG_rl_2_t1 = TR_14 ;
	7'h05 :
		RG_rl_2_t1 = TR_14 ;
	7'h06 :
		RG_rl_2_t1 = TR_14 ;
	7'h07 :
		RG_rl_2_t1 = TR_14 ;
	7'h08 :
		RG_rl_2_t1 = TR_14 ;
	7'h09 :
		RG_rl_2_t1 = TR_14 ;
	7'h0a :
		RG_rl_2_t1 = TR_14 ;
	7'h0b :
		RG_rl_2_t1 = TR_14 ;
	7'h0c :
		RG_rl_2_t1 = TR_14 ;
	7'h0d :
		RG_rl_2_t1 = TR_14 ;
	7'h0e :
		RG_rl_2_t1 = TR_14 ;
	7'h0f :
		RG_rl_2_t1 = TR_14 ;
	7'h10 :
		RG_rl_2_t1 = TR_14 ;
	7'h11 :
		RG_rl_2_t1 = TR_14 ;
	7'h12 :
		RG_rl_2_t1 = TR_14 ;
	7'h13 :
		RG_rl_2_t1 = TR_14 ;
	7'h14 :
		RG_rl_2_t1 = TR_14 ;
	7'h15 :
		RG_rl_2_t1 = TR_14 ;
	7'h16 :
		RG_rl_2_t1 = TR_14 ;
	7'h17 :
		RG_rl_2_t1 = TR_14 ;
	7'h18 :
		RG_rl_2_t1 = TR_14 ;
	7'h19 :
		RG_rl_2_t1 = TR_14 ;
	7'h1a :
		RG_rl_2_t1 = TR_14 ;
	7'h1b :
		RG_rl_2_t1 = TR_14 ;
	7'h1c :
		RG_rl_2_t1 = TR_14 ;
	7'h1d :
		RG_rl_2_t1 = TR_14 ;
	7'h1e :
		RG_rl_2_t1 = TR_14 ;
	7'h1f :
		RG_rl_2_t1 = TR_14 ;
	7'h20 :
		RG_rl_2_t1 = TR_14 ;
	7'h21 :
		RG_rl_2_t1 = TR_14 ;
	7'h22 :
		RG_rl_2_t1 = TR_14 ;
	7'h23 :
		RG_rl_2_t1 = TR_14 ;
	7'h24 :
		RG_rl_2_t1 = TR_14 ;
	7'h25 :
		RG_rl_2_t1 = TR_14 ;
	7'h26 :
		RG_rl_2_t1 = TR_14 ;
	7'h27 :
		RG_rl_2_t1 = TR_14 ;
	7'h28 :
		RG_rl_2_t1 = TR_14 ;
	7'h29 :
		RG_rl_2_t1 = TR_14 ;
	7'h2a :
		RG_rl_2_t1 = TR_14 ;
	7'h2b :
		RG_rl_2_t1 = TR_14 ;
	7'h2c :
		RG_rl_2_t1 = TR_14 ;
	7'h2d :
		RG_rl_2_t1 = TR_14 ;
	7'h2e :
		RG_rl_2_t1 = TR_14 ;
	7'h2f :
		RG_rl_2_t1 = TR_14 ;
	7'h30 :
		RG_rl_2_t1 = TR_14 ;
	7'h31 :
		RG_rl_2_t1 = TR_14 ;
	7'h32 :
		RG_rl_2_t1 = TR_14 ;
	7'h33 :
		RG_rl_2_t1 = TR_14 ;
	7'h34 :
		RG_rl_2_t1 = TR_14 ;
	7'h35 :
		RG_rl_2_t1 = TR_14 ;
	7'h36 :
		RG_rl_2_t1 = TR_14 ;
	7'h37 :
		RG_rl_2_t1 = TR_14 ;
	7'h38 :
		RG_rl_2_t1 = TR_14 ;
	7'h39 :
		RG_rl_2_t1 = TR_14 ;
	7'h3a :
		RG_rl_2_t1 = TR_14 ;
	7'h3b :
		RG_rl_2_t1 = TR_14 ;
	7'h3c :
		RG_rl_2_t1 = TR_14 ;
	7'h3d :
		RG_rl_2_t1 = TR_14 ;
	7'h3e :
		RG_rl_2_t1 = TR_14 ;
	7'h3f :
		RG_rl_2_t1 = TR_14 ;
	7'h40 :
		RG_rl_2_t1 = TR_14 ;
	7'h41 :
		RG_rl_2_t1 = TR_14 ;
	7'h42 :
		RG_rl_2_t1 = TR_14 ;
	7'h43 :
		RG_rl_2_t1 = TR_14 ;
	7'h44 :
		RG_rl_2_t1 = TR_14 ;
	7'h45 :
		RG_rl_2_t1 = TR_14 ;
	7'h46 :
		RG_rl_2_t1 = TR_14 ;
	7'h47 :
		RG_rl_2_t1 = TR_14 ;
	7'h48 :
		RG_rl_2_t1 = TR_14 ;
	7'h49 :
		RG_rl_2_t1 = TR_14 ;
	7'h4a :
		RG_rl_2_t1 = TR_14 ;
	7'h4b :
		RG_rl_2_t1 = TR_14 ;
	7'h4c :
		RG_rl_2_t1 = TR_14 ;
	7'h4d :
		RG_rl_2_t1 = TR_14 ;
	7'h4e :
		RG_rl_2_t1 = TR_14 ;
	7'h4f :
		RG_rl_2_t1 = TR_14 ;
	7'h50 :
		RG_rl_2_t1 = TR_14 ;
	7'h51 :
		RG_rl_2_t1 = TR_14 ;
	7'h52 :
		RG_rl_2_t1 = TR_14 ;
	7'h53 :
		RG_rl_2_t1 = TR_14 ;
	7'h54 :
		RG_rl_2_t1 = TR_14 ;
	7'h55 :
		RG_rl_2_t1 = TR_14 ;
	7'h56 :
		RG_rl_2_t1 = TR_14 ;
	7'h57 :
		RG_rl_2_t1 = TR_14 ;
	7'h58 :
		RG_rl_2_t1 = TR_14 ;
	7'h59 :
		RG_rl_2_t1 = TR_14 ;
	7'h5a :
		RG_rl_2_t1 = TR_14 ;
	7'h5b :
		RG_rl_2_t1 = TR_14 ;
	7'h5c :
		RG_rl_2_t1 = TR_14 ;
	7'h5d :
		RG_rl_2_t1 = TR_14 ;
	7'h5e :
		RG_rl_2_t1 = TR_14 ;
	7'h5f :
		RG_rl_2_t1 = TR_14 ;
	7'h60 :
		RG_rl_2_t1 = TR_14 ;
	7'h61 :
		RG_rl_2_t1 = TR_14 ;
	7'h62 :
		RG_rl_2_t1 = TR_14 ;
	7'h63 :
		RG_rl_2_t1 = TR_14 ;
	7'h64 :
		RG_rl_2_t1 = TR_14 ;
	7'h65 :
		RG_rl_2_t1 = TR_14 ;
	7'h66 :
		RG_rl_2_t1 = TR_14 ;
	7'h67 :
		RG_rl_2_t1 = TR_14 ;
	7'h68 :
		RG_rl_2_t1 = TR_14 ;
	7'h69 :
		RG_rl_2_t1 = TR_14 ;
	7'h6a :
		RG_rl_2_t1 = TR_14 ;
	7'h6b :
		RG_rl_2_t1 = TR_14 ;
	7'h6c :
		RG_rl_2_t1 = TR_14 ;
	7'h6d :
		RG_rl_2_t1 = TR_14 ;
	7'h6e :
		RG_rl_2_t1 = TR_14 ;
	7'h6f :
		RG_rl_2_t1 = TR_14 ;
	7'h70 :
		RG_rl_2_t1 = TR_14 ;
	7'h71 :
		RG_rl_2_t1 = TR_14 ;
	7'h72 :
		RG_rl_2_t1 = TR_14 ;
	7'h73 :
		RG_rl_2_t1 = TR_14 ;
	7'h74 :
		RG_rl_2_t1 = TR_14 ;
	7'h75 :
		RG_rl_2_t1 = TR_14 ;
	7'h76 :
		RG_rl_2_t1 = TR_14 ;
	7'h77 :
		RG_rl_2_t1 = TR_14 ;
	7'h78 :
		RG_rl_2_t1 = TR_14 ;
	7'h79 :
		RG_rl_2_t1 = TR_14 ;
	7'h7a :
		RG_rl_2_t1 = TR_14 ;
	7'h7b :
		RG_rl_2_t1 = TR_14 ;
	7'h7c :
		RG_rl_2_t1 = TR_14 ;
	7'h7d :
		RG_rl_2_t1 = TR_14 ;
	7'h7e :
		RG_rl_2_t1 = TR_14 ;
	7'h7f :
		RG_rl_2_t1 = TR_14 ;
	default :
		RG_rl_2_t1 = 9'hx ;
	endcase
always @ ( RG_rl_2_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_185 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_2_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h02 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_2_t = ( ( { 9{ U_570 } } & RG_rl_185 )
		| ( { 9{ U_569 } } & RG_rl_2_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_2_en = ( U_570 | RG_rl_2_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_2_en )
		RG_rl_2 <= RG_rl_2_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_15 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_3_t1 = TR_15 ;
	7'h01 :
		RG_rl_3_t1 = TR_15 ;
	7'h02 :
		RG_rl_3_t1 = TR_15 ;
	7'h03 :
		RG_rl_3_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h04 :
		RG_rl_3_t1 = TR_15 ;
	7'h05 :
		RG_rl_3_t1 = TR_15 ;
	7'h06 :
		RG_rl_3_t1 = TR_15 ;
	7'h07 :
		RG_rl_3_t1 = TR_15 ;
	7'h08 :
		RG_rl_3_t1 = TR_15 ;
	7'h09 :
		RG_rl_3_t1 = TR_15 ;
	7'h0a :
		RG_rl_3_t1 = TR_15 ;
	7'h0b :
		RG_rl_3_t1 = TR_15 ;
	7'h0c :
		RG_rl_3_t1 = TR_15 ;
	7'h0d :
		RG_rl_3_t1 = TR_15 ;
	7'h0e :
		RG_rl_3_t1 = TR_15 ;
	7'h0f :
		RG_rl_3_t1 = TR_15 ;
	7'h10 :
		RG_rl_3_t1 = TR_15 ;
	7'h11 :
		RG_rl_3_t1 = TR_15 ;
	7'h12 :
		RG_rl_3_t1 = TR_15 ;
	7'h13 :
		RG_rl_3_t1 = TR_15 ;
	7'h14 :
		RG_rl_3_t1 = TR_15 ;
	7'h15 :
		RG_rl_3_t1 = TR_15 ;
	7'h16 :
		RG_rl_3_t1 = TR_15 ;
	7'h17 :
		RG_rl_3_t1 = TR_15 ;
	7'h18 :
		RG_rl_3_t1 = TR_15 ;
	7'h19 :
		RG_rl_3_t1 = TR_15 ;
	7'h1a :
		RG_rl_3_t1 = TR_15 ;
	7'h1b :
		RG_rl_3_t1 = TR_15 ;
	7'h1c :
		RG_rl_3_t1 = TR_15 ;
	7'h1d :
		RG_rl_3_t1 = TR_15 ;
	7'h1e :
		RG_rl_3_t1 = TR_15 ;
	7'h1f :
		RG_rl_3_t1 = TR_15 ;
	7'h20 :
		RG_rl_3_t1 = TR_15 ;
	7'h21 :
		RG_rl_3_t1 = TR_15 ;
	7'h22 :
		RG_rl_3_t1 = TR_15 ;
	7'h23 :
		RG_rl_3_t1 = TR_15 ;
	7'h24 :
		RG_rl_3_t1 = TR_15 ;
	7'h25 :
		RG_rl_3_t1 = TR_15 ;
	7'h26 :
		RG_rl_3_t1 = TR_15 ;
	7'h27 :
		RG_rl_3_t1 = TR_15 ;
	7'h28 :
		RG_rl_3_t1 = TR_15 ;
	7'h29 :
		RG_rl_3_t1 = TR_15 ;
	7'h2a :
		RG_rl_3_t1 = TR_15 ;
	7'h2b :
		RG_rl_3_t1 = TR_15 ;
	7'h2c :
		RG_rl_3_t1 = TR_15 ;
	7'h2d :
		RG_rl_3_t1 = TR_15 ;
	7'h2e :
		RG_rl_3_t1 = TR_15 ;
	7'h2f :
		RG_rl_3_t1 = TR_15 ;
	7'h30 :
		RG_rl_3_t1 = TR_15 ;
	7'h31 :
		RG_rl_3_t1 = TR_15 ;
	7'h32 :
		RG_rl_3_t1 = TR_15 ;
	7'h33 :
		RG_rl_3_t1 = TR_15 ;
	7'h34 :
		RG_rl_3_t1 = TR_15 ;
	7'h35 :
		RG_rl_3_t1 = TR_15 ;
	7'h36 :
		RG_rl_3_t1 = TR_15 ;
	7'h37 :
		RG_rl_3_t1 = TR_15 ;
	7'h38 :
		RG_rl_3_t1 = TR_15 ;
	7'h39 :
		RG_rl_3_t1 = TR_15 ;
	7'h3a :
		RG_rl_3_t1 = TR_15 ;
	7'h3b :
		RG_rl_3_t1 = TR_15 ;
	7'h3c :
		RG_rl_3_t1 = TR_15 ;
	7'h3d :
		RG_rl_3_t1 = TR_15 ;
	7'h3e :
		RG_rl_3_t1 = TR_15 ;
	7'h3f :
		RG_rl_3_t1 = TR_15 ;
	7'h40 :
		RG_rl_3_t1 = TR_15 ;
	7'h41 :
		RG_rl_3_t1 = TR_15 ;
	7'h42 :
		RG_rl_3_t1 = TR_15 ;
	7'h43 :
		RG_rl_3_t1 = TR_15 ;
	7'h44 :
		RG_rl_3_t1 = TR_15 ;
	7'h45 :
		RG_rl_3_t1 = TR_15 ;
	7'h46 :
		RG_rl_3_t1 = TR_15 ;
	7'h47 :
		RG_rl_3_t1 = TR_15 ;
	7'h48 :
		RG_rl_3_t1 = TR_15 ;
	7'h49 :
		RG_rl_3_t1 = TR_15 ;
	7'h4a :
		RG_rl_3_t1 = TR_15 ;
	7'h4b :
		RG_rl_3_t1 = TR_15 ;
	7'h4c :
		RG_rl_3_t1 = TR_15 ;
	7'h4d :
		RG_rl_3_t1 = TR_15 ;
	7'h4e :
		RG_rl_3_t1 = TR_15 ;
	7'h4f :
		RG_rl_3_t1 = TR_15 ;
	7'h50 :
		RG_rl_3_t1 = TR_15 ;
	7'h51 :
		RG_rl_3_t1 = TR_15 ;
	7'h52 :
		RG_rl_3_t1 = TR_15 ;
	7'h53 :
		RG_rl_3_t1 = TR_15 ;
	7'h54 :
		RG_rl_3_t1 = TR_15 ;
	7'h55 :
		RG_rl_3_t1 = TR_15 ;
	7'h56 :
		RG_rl_3_t1 = TR_15 ;
	7'h57 :
		RG_rl_3_t1 = TR_15 ;
	7'h58 :
		RG_rl_3_t1 = TR_15 ;
	7'h59 :
		RG_rl_3_t1 = TR_15 ;
	7'h5a :
		RG_rl_3_t1 = TR_15 ;
	7'h5b :
		RG_rl_3_t1 = TR_15 ;
	7'h5c :
		RG_rl_3_t1 = TR_15 ;
	7'h5d :
		RG_rl_3_t1 = TR_15 ;
	7'h5e :
		RG_rl_3_t1 = TR_15 ;
	7'h5f :
		RG_rl_3_t1 = TR_15 ;
	7'h60 :
		RG_rl_3_t1 = TR_15 ;
	7'h61 :
		RG_rl_3_t1 = TR_15 ;
	7'h62 :
		RG_rl_3_t1 = TR_15 ;
	7'h63 :
		RG_rl_3_t1 = TR_15 ;
	7'h64 :
		RG_rl_3_t1 = TR_15 ;
	7'h65 :
		RG_rl_3_t1 = TR_15 ;
	7'h66 :
		RG_rl_3_t1 = TR_15 ;
	7'h67 :
		RG_rl_3_t1 = TR_15 ;
	7'h68 :
		RG_rl_3_t1 = TR_15 ;
	7'h69 :
		RG_rl_3_t1 = TR_15 ;
	7'h6a :
		RG_rl_3_t1 = TR_15 ;
	7'h6b :
		RG_rl_3_t1 = TR_15 ;
	7'h6c :
		RG_rl_3_t1 = TR_15 ;
	7'h6d :
		RG_rl_3_t1 = TR_15 ;
	7'h6e :
		RG_rl_3_t1 = TR_15 ;
	7'h6f :
		RG_rl_3_t1 = TR_15 ;
	7'h70 :
		RG_rl_3_t1 = TR_15 ;
	7'h71 :
		RG_rl_3_t1 = TR_15 ;
	7'h72 :
		RG_rl_3_t1 = TR_15 ;
	7'h73 :
		RG_rl_3_t1 = TR_15 ;
	7'h74 :
		RG_rl_3_t1 = TR_15 ;
	7'h75 :
		RG_rl_3_t1 = TR_15 ;
	7'h76 :
		RG_rl_3_t1 = TR_15 ;
	7'h77 :
		RG_rl_3_t1 = TR_15 ;
	7'h78 :
		RG_rl_3_t1 = TR_15 ;
	7'h79 :
		RG_rl_3_t1 = TR_15 ;
	7'h7a :
		RG_rl_3_t1 = TR_15 ;
	7'h7b :
		RG_rl_3_t1 = TR_15 ;
	7'h7c :
		RG_rl_3_t1 = TR_15 ;
	7'h7d :
		RG_rl_3_t1 = TR_15 ;
	7'h7e :
		RG_rl_3_t1 = TR_15 ;
	7'h7f :
		RG_rl_3_t1 = TR_15 ;
	default :
		RG_rl_3_t1 = 9'hx ;
	endcase
always @ ( RG_rl_3_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_186 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_3_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h03 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_3_t = ( ( { 9{ U_570 } } & RG_rl_186 )
		| ( { 9{ U_569 } } & RG_rl_3_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_3_en = ( U_570 | RG_rl_3_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_3_en )
		RG_rl_3 <= RG_rl_3_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_16 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_4_t1 = TR_16 ;
	7'h01 :
		RG_rl_4_t1 = TR_16 ;
	7'h02 :
		RG_rl_4_t1 = TR_16 ;
	7'h03 :
		RG_rl_4_t1 = TR_16 ;
	7'h04 :
		RG_rl_4_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h05 :
		RG_rl_4_t1 = TR_16 ;
	7'h06 :
		RG_rl_4_t1 = TR_16 ;
	7'h07 :
		RG_rl_4_t1 = TR_16 ;
	7'h08 :
		RG_rl_4_t1 = TR_16 ;
	7'h09 :
		RG_rl_4_t1 = TR_16 ;
	7'h0a :
		RG_rl_4_t1 = TR_16 ;
	7'h0b :
		RG_rl_4_t1 = TR_16 ;
	7'h0c :
		RG_rl_4_t1 = TR_16 ;
	7'h0d :
		RG_rl_4_t1 = TR_16 ;
	7'h0e :
		RG_rl_4_t1 = TR_16 ;
	7'h0f :
		RG_rl_4_t1 = TR_16 ;
	7'h10 :
		RG_rl_4_t1 = TR_16 ;
	7'h11 :
		RG_rl_4_t1 = TR_16 ;
	7'h12 :
		RG_rl_4_t1 = TR_16 ;
	7'h13 :
		RG_rl_4_t1 = TR_16 ;
	7'h14 :
		RG_rl_4_t1 = TR_16 ;
	7'h15 :
		RG_rl_4_t1 = TR_16 ;
	7'h16 :
		RG_rl_4_t1 = TR_16 ;
	7'h17 :
		RG_rl_4_t1 = TR_16 ;
	7'h18 :
		RG_rl_4_t1 = TR_16 ;
	7'h19 :
		RG_rl_4_t1 = TR_16 ;
	7'h1a :
		RG_rl_4_t1 = TR_16 ;
	7'h1b :
		RG_rl_4_t1 = TR_16 ;
	7'h1c :
		RG_rl_4_t1 = TR_16 ;
	7'h1d :
		RG_rl_4_t1 = TR_16 ;
	7'h1e :
		RG_rl_4_t1 = TR_16 ;
	7'h1f :
		RG_rl_4_t1 = TR_16 ;
	7'h20 :
		RG_rl_4_t1 = TR_16 ;
	7'h21 :
		RG_rl_4_t1 = TR_16 ;
	7'h22 :
		RG_rl_4_t1 = TR_16 ;
	7'h23 :
		RG_rl_4_t1 = TR_16 ;
	7'h24 :
		RG_rl_4_t1 = TR_16 ;
	7'h25 :
		RG_rl_4_t1 = TR_16 ;
	7'h26 :
		RG_rl_4_t1 = TR_16 ;
	7'h27 :
		RG_rl_4_t1 = TR_16 ;
	7'h28 :
		RG_rl_4_t1 = TR_16 ;
	7'h29 :
		RG_rl_4_t1 = TR_16 ;
	7'h2a :
		RG_rl_4_t1 = TR_16 ;
	7'h2b :
		RG_rl_4_t1 = TR_16 ;
	7'h2c :
		RG_rl_4_t1 = TR_16 ;
	7'h2d :
		RG_rl_4_t1 = TR_16 ;
	7'h2e :
		RG_rl_4_t1 = TR_16 ;
	7'h2f :
		RG_rl_4_t1 = TR_16 ;
	7'h30 :
		RG_rl_4_t1 = TR_16 ;
	7'h31 :
		RG_rl_4_t1 = TR_16 ;
	7'h32 :
		RG_rl_4_t1 = TR_16 ;
	7'h33 :
		RG_rl_4_t1 = TR_16 ;
	7'h34 :
		RG_rl_4_t1 = TR_16 ;
	7'h35 :
		RG_rl_4_t1 = TR_16 ;
	7'h36 :
		RG_rl_4_t1 = TR_16 ;
	7'h37 :
		RG_rl_4_t1 = TR_16 ;
	7'h38 :
		RG_rl_4_t1 = TR_16 ;
	7'h39 :
		RG_rl_4_t1 = TR_16 ;
	7'h3a :
		RG_rl_4_t1 = TR_16 ;
	7'h3b :
		RG_rl_4_t1 = TR_16 ;
	7'h3c :
		RG_rl_4_t1 = TR_16 ;
	7'h3d :
		RG_rl_4_t1 = TR_16 ;
	7'h3e :
		RG_rl_4_t1 = TR_16 ;
	7'h3f :
		RG_rl_4_t1 = TR_16 ;
	7'h40 :
		RG_rl_4_t1 = TR_16 ;
	7'h41 :
		RG_rl_4_t1 = TR_16 ;
	7'h42 :
		RG_rl_4_t1 = TR_16 ;
	7'h43 :
		RG_rl_4_t1 = TR_16 ;
	7'h44 :
		RG_rl_4_t1 = TR_16 ;
	7'h45 :
		RG_rl_4_t1 = TR_16 ;
	7'h46 :
		RG_rl_4_t1 = TR_16 ;
	7'h47 :
		RG_rl_4_t1 = TR_16 ;
	7'h48 :
		RG_rl_4_t1 = TR_16 ;
	7'h49 :
		RG_rl_4_t1 = TR_16 ;
	7'h4a :
		RG_rl_4_t1 = TR_16 ;
	7'h4b :
		RG_rl_4_t1 = TR_16 ;
	7'h4c :
		RG_rl_4_t1 = TR_16 ;
	7'h4d :
		RG_rl_4_t1 = TR_16 ;
	7'h4e :
		RG_rl_4_t1 = TR_16 ;
	7'h4f :
		RG_rl_4_t1 = TR_16 ;
	7'h50 :
		RG_rl_4_t1 = TR_16 ;
	7'h51 :
		RG_rl_4_t1 = TR_16 ;
	7'h52 :
		RG_rl_4_t1 = TR_16 ;
	7'h53 :
		RG_rl_4_t1 = TR_16 ;
	7'h54 :
		RG_rl_4_t1 = TR_16 ;
	7'h55 :
		RG_rl_4_t1 = TR_16 ;
	7'h56 :
		RG_rl_4_t1 = TR_16 ;
	7'h57 :
		RG_rl_4_t1 = TR_16 ;
	7'h58 :
		RG_rl_4_t1 = TR_16 ;
	7'h59 :
		RG_rl_4_t1 = TR_16 ;
	7'h5a :
		RG_rl_4_t1 = TR_16 ;
	7'h5b :
		RG_rl_4_t1 = TR_16 ;
	7'h5c :
		RG_rl_4_t1 = TR_16 ;
	7'h5d :
		RG_rl_4_t1 = TR_16 ;
	7'h5e :
		RG_rl_4_t1 = TR_16 ;
	7'h5f :
		RG_rl_4_t1 = TR_16 ;
	7'h60 :
		RG_rl_4_t1 = TR_16 ;
	7'h61 :
		RG_rl_4_t1 = TR_16 ;
	7'h62 :
		RG_rl_4_t1 = TR_16 ;
	7'h63 :
		RG_rl_4_t1 = TR_16 ;
	7'h64 :
		RG_rl_4_t1 = TR_16 ;
	7'h65 :
		RG_rl_4_t1 = TR_16 ;
	7'h66 :
		RG_rl_4_t1 = TR_16 ;
	7'h67 :
		RG_rl_4_t1 = TR_16 ;
	7'h68 :
		RG_rl_4_t1 = TR_16 ;
	7'h69 :
		RG_rl_4_t1 = TR_16 ;
	7'h6a :
		RG_rl_4_t1 = TR_16 ;
	7'h6b :
		RG_rl_4_t1 = TR_16 ;
	7'h6c :
		RG_rl_4_t1 = TR_16 ;
	7'h6d :
		RG_rl_4_t1 = TR_16 ;
	7'h6e :
		RG_rl_4_t1 = TR_16 ;
	7'h6f :
		RG_rl_4_t1 = TR_16 ;
	7'h70 :
		RG_rl_4_t1 = TR_16 ;
	7'h71 :
		RG_rl_4_t1 = TR_16 ;
	7'h72 :
		RG_rl_4_t1 = TR_16 ;
	7'h73 :
		RG_rl_4_t1 = TR_16 ;
	7'h74 :
		RG_rl_4_t1 = TR_16 ;
	7'h75 :
		RG_rl_4_t1 = TR_16 ;
	7'h76 :
		RG_rl_4_t1 = TR_16 ;
	7'h77 :
		RG_rl_4_t1 = TR_16 ;
	7'h78 :
		RG_rl_4_t1 = TR_16 ;
	7'h79 :
		RG_rl_4_t1 = TR_16 ;
	7'h7a :
		RG_rl_4_t1 = TR_16 ;
	7'h7b :
		RG_rl_4_t1 = TR_16 ;
	7'h7c :
		RG_rl_4_t1 = TR_16 ;
	7'h7d :
		RG_rl_4_t1 = TR_16 ;
	7'h7e :
		RG_rl_4_t1 = TR_16 ;
	7'h7f :
		RG_rl_4_t1 = TR_16 ;
	default :
		RG_rl_4_t1 = 9'hx ;
	endcase
always @ ( RG_rl_4_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_187 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_4_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h04 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_4_t = ( ( { 9{ U_570 } } & RG_rl_187 )
		| ( { 9{ U_569 } } & RG_rl_4_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_4_en = ( U_570 | RG_rl_4_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_4_en )
		RG_rl_4 <= RG_rl_4_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_17 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_5_t1 = TR_17 ;
	7'h01 :
		RG_rl_5_t1 = TR_17 ;
	7'h02 :
		RG_rl_5_t1 = TR_17 ;
	7'h03 :
		RG_rl_5_t1 = TR_17 ;
	7'h04 :
		RG_rl_5_t1 = TR_17 ;
	7'h05 :
		RG_rl_5_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h06 :
		RG_rl_5_t1 = TR_17 ;
	7'h07 :
		RG_rl_5_t1 = TR_17 ;
	7'h08 :
		RG_rl_5_t1 = TR_17 ;
	7'h09 :
		RG_rl_5_t1 = TR_17 ;
	7'h0a :
		RG_rl_5_t1 = TR_17 ;
	7'h0b :
		RG_rl_5_t1 = TR_17 ;
	7'h0c :
		RG_rl_5_t1 = TR_17 ;
	7'h0d :
		RG_rl_5_t1 = TR_17 ;
	7'h0e :
		RG_rl_5_t1 = TR_17 ;
	7'h0f :
		RG_rl_5_t1 = TR_17 ;
	7'h10 :
		RG_rl_5_t1 = TR_17 ;
	7'h11 :
		RG_rl_5_t1 = TR_17 ;
	7'h12 :
		RG_rl_5_t1 = TR_17 ;
	7'h13 :
		RG_rl_5_t1 = TR_17 ;
	7'h14 :
		RG_rl_5_t1 = TR_17 ;
	7'h15 :
		RG_rl_5_t1 = TR_17 ;
	7'h16 :
		RG_rl_5_t1 = TR_17 ;
	7'h17 :
		RG_rl_5_t1 = TR_17 ;
	7'h18 :
		RG_rl_5_t1 = TR_17 ;
	7'h19 :
		RG_rl_5_t1 = TR_17 ;
	7'h1a :
		RG_rl_5_t1 = TR_17 ;
	7'h1b :
		RG_rl_5_t1 = TR_17 ;
	7'h1c :
		RG_rl_5_t1 = TR_17 ;
	7'h1d :
		RG_rl_5_t1 = TR_17 ;
	7'h1e :
		RG_rl_5_t1 = TR_17 ;
	7'h1f :
		RG_rl_5_t1 = TR_17 ;
	7'h20 :
		RG_rl_5_t1 = TR_17 ;
	7'h21 :
		RG_rl_5_t1 = TR_17 ;
	7'h22 :
		RG_rl_5_t1 = TR_17 ;
	7'h23 :
		RG_rl_5_t1 = TR_17 ;
	7'h24 :
		RG_rl_5_t1 = TR_17 ;
	7'h25 :
		RG_rl_5_t1 = TR_17 ;
	7'h26 :
		RG_rl_5_t1 = TR_17 ;
	7'h27 :
		RG_rl_5_t1 = TR_17 ;
	7'h28 :
		RG_rl_5_t1 = TR_17 ;
	7'h29 :
		RG_rl_5_t1 = TR_17 ;
	7'h2a :
		RG_rl_5_t1 = TR_17 ;
	7'h2b :
		RG_rl_5_t1 = TR_17 ;
	7'h2c :
		RG_rl_5_t1 = TR_17 ;
	7'h2d :
		RG_rl_5_t1 = TR_17 ;
	7'h2e :
		RG_rl_5_t1 = TR_17 ;
	7'h2f :
		RG_rl_5_t1 = TR_17 ;
	7'h30 :
		RG_rl_5_t1 = TR_17 ;
	7'h31 :
		RG_rl_5_t1 = TR_17 ;
	7'h32 :
		RG_rl_5_t1 = TR_17 ;
	7'h33 :
		RG_rl_5_t1 = TR_17 ;
	7'h34 :
		RG_rl_5_t1 = TR_17 ;
	7'h35 :
		RG_rl_5_t1 = TR_17 ;
	7'h36 :
		RG_rl_5_t1 = TR_17 ;
	7'h37 :
		RG_rl_5_t1 = TR_17 ;
	7'h38 :
		RG_rl_5_t1 = TR_17 ;
	7'h39 :
		RG_rl_5_t1 = TR_17 ;
	7'h3a :
		RG_rl_5_t1 = TR_17 ;
	7'h3b :
		RG_rl_5_t1 = TR_17 ;
	7'h3c :
		RG_rl_5_t1 = TR_17 ;
	7'h3d :
		RG_rl_5_t1 = TR_17 ;
	7'h3e :
		RG_rl_5_t1 = TR_17 ;
	7'h3f :
		RG_rl_5_t1 = TR_17 ;
	7'h40 :
		RG_rl_5_t1 = TR_17 ;
	7'h41 :
		RG_rl_5_t1 = TR_17 ;
	7'h42 :
		RG_rl_5_t1 = TR_17 ;
	7'h43 :
		RG_rl_5_t1 = TR_17 ;
	7'h44 :
		RG_rl_5_t1 = TR_17 ;
	7'h45 :
		RG_rl_5_t1 = TR_17 ;
	7'h46 :
		RG_rl_5_t1 = TR_17 ;
	7'h47 :
		RG_rl_5_t1 = TR_17 ;
	7'h48 :
		RG_rl_5_t1 = TR_17 ;
	7'h49 :
		RG_rl_5_t1 = TR_17 ;
	7'h4a :
		RG_rl_5_t1 = TR_17 ;
	7'h4b :
		RG_rl_5_t1 = TR_17 ;
	7'h4c :
		RG_rl_5_t1 = TR_17 ;
	7'h4d :
		RG_rl_5_t1 = TR_17 ;
	7'h4e :
		RG_rl_5_t1 = TR_17 ;
	7'h4f :
		RG_rl_5_t1 = TR_17 ;
	7'h50 :
		RG_rl_5_t1 = TR_17 ;
	7'h51 :
		RG_rl_5_t1 = TR_17 ;
	7'h52 :
		RG_rl_5_t1 = TR_17 ;
	7'h53 :
		RG_rl_5_t1 = TR_17 ;
	7'h54 :
		RG_rl_5_t1 = TR_17 ;
	7'h55 :
		RG_rl_5_t1 = TR_17 ;
	7'h56 :
		RG_rl_5_t1 = TR_17 ;
	7'h57 :
		RG_rl_5_t1 = TR_17 ;
	7'h58 :
		RG_rl_5_t1 = TR_17 ;
	7'h59 :
		RG_rl_5_t1 = TR_17 ;
	7'h5a :
		RG_rl_5_t1 = TR_17 ;
	7'h5b :
		RG_rl_5_t1 = TR_17 ;
	7'h5c :
		RG_rl_5_t1 = TR_17 ;
	7'h5d :
		RG_rl_5_t1 = TR_17 ;
	7'h5e :
		RG_rl_5_t1 = TR_17 ;
	7'h5f :
		RG_rl_5_t1 = TR_17 ;
	7'h60 :
		RG_rl_5_t1 = TR_17 ;
	7'h61 :
		RG_rl_5_t1 = TR_17 ;
	7'h62 :
		RG_rl_5_t1 = TR_17 ;
	7'h63 :
		RG_rl_5_t1 = TR_17 ;
	7'h64 :
		RG_rl_5_t1 = TR_17 ;
	7'h65 :
		RG_rl_5_t1 = TR_17 ;
	7'h66 :
		RG_rl_5_t1 = TR_17 ;
	7'h67 :
		RG_rl_5_t1 = TR_17 ;
	7'h68 :
		RG_rl_5_t1 = TR_17 ;
	7'h69 :
		RG_rl_5_t1 = TR_17 ;
	7'h6a :
		RG_rl_5_t1 = TR_17 ;
	7'h6b :
		RG_rl_5_t1 = TR_17 ;
	7'h6c :
		RG_rl_5_t1 = TR_17 ;
	7'h6d :
		RG_rl_5_t1 = TR_17 ;
	7'h6e :
		RG_rl_5_t1 = TR_17 ;
	7'h6f :
		RG_rl_5_t1 = TR_17 ;
	7'h70 :
		RG_rl_5_t1 = TR_17 ;
	7'h71 :
		RG_rl_5_t1 = TR_17 ;
	7'h72 :
		RG_rl_5_t1 = TR_17 ;
	7'h73 :
		RG_rl_5_t1 = TR_17 ;
	7'h74 :
		RG_rl_5_t1 = TR_17 ;
	7'h75 :
		RG_rl_5_t1 = TR_17 ;
	7'h76 :
		RG_rl_5_t1 = TR_17 ;
	7'h77 :
		RG_rl_5_t1 = TR_17 ;
	7'h78 :
		RG_rl_5_t1 = TR_17 ;
	7'h79 :
		RG_rl_5_t1 = TR_17 ;
	7'h7a :
		RG_rl_5_t1 = TR_17 ;
	7'h7b :
		RG_rl_5_t1 = TR_17 ;
	7'h7c :
		RG_rl_5_t1 = TR_17 ;
	7'h7d :
		RG_rl_5_t1 = TR_17 ;
	7'h7e :
		RG_rl_5_t1 = TR_17 ;
	7'h7f :
		RG_rl_5_t1 = TR_17 ;
	default :
		RG_rl_5_t1 = 9'hx ;
	endcase
always @ ( RG_rl_5_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_188 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_5_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h05 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_5_t = ( ( { 9{ U_570 } } & RG_rl_188 )
		| ( { 9{ U_569 } } & RG_rl_5_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_5_en = ( U_570 | RG_rl_5_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_5_en )
		RG_rl_5 <= RG_rl_5_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_18 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_6_t1 = TR_18 ;
	7'h01 :
		RG_rl_6_t1 = TR_18 ;
	7'h02 :
		RG_rl_6_t1 = TR_18 ;
	7'h03 :
		RG_rl_6_t1 = TR_18 ;
	7'h04 :
		RG_rl_6_t1 = TR_18 ;
	7'h05 :
		RG_rl_6_t1 = TR_18 ;
	7'h06 :
		RG_rl_6_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h07 :
		RG_rl_6_t1 = TR_18 ;
	7'h08 :
		RG_rl_6_t1 = TR_18 ;
	7'h09 :
		RG_rl_6_t1 = TR_18 ;
	7'h0a :
		RG_rl_6_t1 = TR_18 ;
	7'h0b :
		RG_rl_6_t1 = TR_18 ;
	7'h0c :
		RG_rl_6_t1 = TR_18 ;
	7'h0d :
		RG_rl_6_t1 = TR_18 ;
	7'h0e :
		RG_rl_6_t1 = TR_18 ;
	7'h0f :
		RG_rl_6_t1 = TR_18 ;
	7'h10 :
		RG_rl_6_t1 = TR_18 ;
	7'h11 :
		RG_rl_6_t1 = TR_18 ;
	7'h12 :
		RG_rl_6_t1 = TR_18 ;
	7'h13 :
		RG_rl_6_t1 = TR_18 ;
	7'h14 :
		RG_rl_6_t1 = TR_18 ;
	7'h15 :
		RG_rl_6_t1 = TR_18 ;
	7'h16 :
		RG_rl_6_t1 = TR_18 ;
	7'h17 :
		RG_rl_6_t1 = TR_18 ;
	7'h18 :
		RG_rl_6_t1 = TR_18 ;
	7'h19 :
		RG_rl_6_t1 = TR_18 ;
	7'h1a :
		RG_rl_6_t1 = TR_18 ;
	7'h1b :
		RG_rl_6_t1 = TR_18 ;
	7'h1c :
		RG_rl_6_t1 = TR_18 ;
	7'h1d :
		RG_rl_6_t1 = TR_18 ;
	7'h1e :
		RG_rl_6_t1 = TR_18 ;
	7'h1f :
		RG_rl_6_t1 = TR_18 ;
	7'h20 :
		RG_rl_6_t1 = TR_18 ;
	7'h21 :
		RG_rl_6_t1 = TR_18 ;
	7'h22 :
		RG_rl_6_t1 = TR_18 ;
	7'h23 :
		RG_rl_6_t1 = TR_18 ;
	7'h24 :
		RG_rl_6_t1 = TR_18 ;
	7'h25 :
		RG_rl_6_t1 = TR_18 ;
	7'h26 :
		RG_rl_6_t1 = TR_18 ;
	7'h27 :
		RG_rl_6_t1 = TR_18 ;
	7'h28 :
		RG_rl_6_t1 = TR_18 ;
	7'h29 :
		RG_rl_6_t1 = TR_18 ;
	7'h2a :
		RG_rl_6_t1 = TR_18 ;
	7'h2b :
		RG_rl_6_t1 = TR_18 ;
	7'h2c :
		RG_rl_6_t1 = TR_18 ;
	7'h2d :
		RG_rl_6_t1 = TR_18 ;
	7'h2e :
		RG_rl_6_t1 = TR_18 ;
	7'h2f :
		RG_rl_6_t1 = TR_18 ;
	7'h30 :
		RG_rl_6_t1 = TR_18 ;
	7'h31 :
		RG_rl_6_t1 = TR_18 ;
	7'h32 :
		RG_rl_6_t1 = TR_18 ;
	7'h33 :
		RG_rl_6_t1 = TR_18 ;
	7'h34 :
		RG_rl_6_t1 = TR_18 ;
	7'h35 :
		RG_rl_6_t1 = TR_18 ;
	7'h36 :
		RG_rl_6_t1 = TR_18 ;
	7'h37 :
		RG_rl_6_t1 = TR_18 ;
	7'h38 :
		RG_rl_6_t1 = TR_18 ;
	7'h39 :
		RG_rl_6_t1 = TR_18 ;
	7'h3a :
		RG_rl_6_t1 = TR_18 ;
	7'h3b :
		RG_rl_6_t1 = TR_18 ;
	7'h3c :
		RG_rl_6_t1 = TR_18 ;
	7'h3d :
		RG_rl_6_t1 = TR_18 ;
	7'h3e :
		RG_rl_6_t1 = TR_18 ;
	7'h3f :
		RG_rl_6_t1 = TR_18 ;
	7'h40 :
		RG_rl_6_t1 = TR_18 ;
	7'h41 :
		RG_rl_6_t1 = TR_18 ;
	7'h42 :
		RG_rl_6_t1 = TR_18 ;
	7'h43 :
		RG_rl_6_t1 = TR_18 ;
	7'h44 :
		RG_rl_6_t1 = TR_18 ;
	7'h45 :
		RG_rl_6_t1 = TR_18 ;
	7'h46 :
		RG_rl_6_t1 = TR_18 ;
	7'h47 :
		RG_rl_6_t1 = TR_18 ;
	7'h48 :
		RG_rl_6_t1 = TR_18 ;
	7'h49 :
		RG_rl_6_t1 = TR_18 ;
	7'h4a :
		RG_rl_6_t1 = TR_18 ;
	7'h4b :
		RG_rl_6_t1 = TR_18 ;
	7'h4c :
		RG_rl_6_t1 = TR_18 ;
	7'h4d :
		RG_rl_6_t1 = TR_18 ;
	7'h4e :
		RG_rl_6_t1 = TR_18 ;
	7'h4f :
		RG_rl_6_t1 = TR_18 ;
	7'h50 :
		RG_rl_6_t1 = TR_18 ;
	7'h51 :
		RG_rl_6_t1 = TR_18 ;
	7'h52 :
		RG_rl_6_t1 = TR_18 ;
	7'h53 :
		RG_rl_6_t1 = TR_18 ;
	7'h54 :
		RG_rl_6_t1 = TR_18 ;
	7'h55 :
		RG_rl_6_t1 = TR_18 ;
	7'h56 :
		RG_rl_6_t1 = TR_18 ;
	7'h57 :
		RG_rl_6_t1 = TR_18 ;
	7'h58 :
		RG_rl_6_t1 = TR_18 ;
	7'h59 :
		RG_rl_6_t1 = TR_18 ;
	7'h5a :
		RG_rl_6_t1 = TR_18 ;
	7'h5b :
		RG_rl_6_t1 = TR_18 ;
	7'h5c :
		RG_rl_6_t1 = TR_18 ;
	7'h5d :
		RG_rl_6_t1 = TR_18 ;
	7'h5e :
		RG_rl_6_t1 = TR_18 ;
	7'h5f :
		RG_rl_6_t1 = TR_18 ;
	7'h60 :
		RG_rl_6_t1 = TR_18 ;
	7'h61 :
		RG_rl_6_t1 = TR_18 ;
	7'h62 :
		RG_rl_6_t1 = TR_18 ;
	7'h63 :
		RG_rl_6_t1 = TR_18 ;
	7'h64 :
		RG_rl_6_t1 = TR_18 ;
	7'h65 :
		RG_rl_6_t1 = TR_18 ;
	7'h66 :
		RG_rl_6_t1 = TR_18 ;
	7'h67 :
		RG_rl_6_t1 = TR_18 ;
	7'h68 :
		RG_rl_6_t1 = TR_18 ;
	7'h69 :
		RG_rl_6_t1 = TR_18 ;
	7'h6a :
		RG_rl_6_t1 = TR_18 ;
	7'h6b :
		RG_rl_6_t1 = TR_18 ;
	7'h6c :
		RG_rl_6_t1 = TR_18 ;
	7'h6d :
		RG_rl_6_t1 = TR_18 ;
	7'h6e :
		RG_rl_6_t1 = TR_18 ;
	7'h6f :
		RG_rl_6_t1 = TR_18 ;
	7'h70 :
		RG_rl_6_t1 = TR_18 ;
	7'h71 :
		RG_rl_6_t1 = TR_18 ;
	7'h72 :
		RG_rl_6_t1 = TR_18 ;
	7'h73 :
		RG_rl_6_t1 = TR_18 ;
	7'h74 :
		RG_rl_6_t1 = TR_18 ;
	7'h75 :
		RG_rl_6_t1 = TR_18 ;
	7'h76 :
		RG_rl_6_t1 = TR_18 ;
	7'h77 :
		RG_rl_6_t1 = TR_18 ;
	7'h78 :
		RG_rl_6_t1 = TR_18 ;
	7'h79 :
		RG_rl_6_t1 = TR_18 ;
	7'h7a :
		RG_rl_6_t1 = TR_18 ;
	7'h7b :
		RG_rl_6_t1 = TR_18 ;
	7'h7c :
		RG_rl_6_t1 = TR_18 ;
	7'h7d :
		RG_rl_6_t1 = TR_18 ;
	7'h7e :
		RG_rl_6_t1 = TR_18 ;
	7'h7f :
		RG_rl_6_t1 = TR_18 ;
	default :
		RG_rl_6_t1 = 9'hx ;
	endcase
always @ ( RG_rl_6_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_189 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_6_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h06 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_6_t = ( ( { 9{ U_570 } } & RG_rl_189 )
		| ( { 9{ U_569 } } & RG_rl_6_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_6_en = ( U_570 | RG_rl_6_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_6_en )
		RG_rl_6 <= RG_rl_6_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_19 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_7_t1 = TR_19 ;
	7'h01 :
		RG_rl_7_t1 = TR_19 ;
	7'h02 :
		RG_rl_7_t1 = TR_19 ;
	7'h03 :
		RG_rl_7_t1 = TR_19 ;
	7'h04 :
		RG_rl_7_t1 = TR_19 ;
	7'h05 :
		RG_rl_7_t1 = TR_19 ;
	7'h06 :
		RG_rl_7_t1 = TR_19 ;
	7'h07 :
		RG_rl_7_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h08 :
		RG_rl_7_t1 = TR_19 ;
	7'h09 :
		RG_rl_7_t1 = TR_19 ;
	7'h0a :
		RG_rl_7_t1 = TR_19 ;
	7'h0b :
		RG_rl_7_t1 = TR_19 ;
	7'h0c :
		RG_rl_7_t1 = TR_19 ;
	7'h0d :
		RG_rl_7_t1 = TR_19 ;
	7'h0e :
		RG_rl_7_t1 = TR_19 ;
	7'h0f :
		RG_rl_7_t1 = TR_19 ;
	7'h10 :
		RG_rl_7_t1 = TR_19 ;
	7'h11 :
		RG_rl_7_t1 = TR_19 ;
	7'h12 :
		RG_rl_7_t1 = TR_19 ;
	7'h13 :
		RG_rl_7_t1 = TR_19 ;
	7'h14 :
		RG_rl_7_t1 = TR_19 ;
	7'h15 :
		RG_rl_7_t1 = TR_19 ;
	7'h16 :
		RG_rl_7_t1 = TR_19 ;
	7'h17 :
		RG_rl_7_t1 = TR_19 ;
	7'h18 :
		RG_rl_7_t1 = TR_19 ;
	7'h19 :
		RG_rl_7_t1 = TR_19 ;
	7'h1a :
		RG_rl_7_t1 = TR_19 ;
	7'h1b :
		RG_rl_7_t1 = TR_19 ;
	7'h1c :
		RG_rl_7_t1 = TR_19 ;
	7'h1d :
		RG_rl_7_t1 = TR_19 ;
	7'h1e :
		RG_rl_7_t1 = TR_19 ;
	7'h1f :
		RG_rl_7_t1 = TR_19 ;
	7'h20 :
		RG_rl_7_t1 = TR_19 ;
	7'h21 :
		RG_rl_7_t1 = TR_19 ;
	7'h22 :
		RG_rl_7_t1 = TR_19 ;
	7'h23 :
		RG_rl_7_t1 = TR_19 ;
	7'h24 :
		RG_rl_7_t1 = TR_19 ;
	7'h25 :
		RG_rl_7_t1 = TR_19 ;
	7'h26 :
		RG_rl_7_t1 = TR_19 ;
	7'h27 :
		RG_rl_7_t1 = TR_19 ;
	7'h28 :
		RG_rl_7_t1 = TR_19 ;
	7'h29 :
		RG_rl_7_t1 = TR_19 ;
	7'h2a :
		RG_rl_7_t1 = TR_19 ;
	7'h2b :
		RG_rl_7_t1 = TR_19 ;
	7'h2c :
		RG_rl_7_t1 = TR_19 ;
	7'h2d :
		RG_rl_7_t1 = TR_19 ;
	7'h2e :
		RG_rl_7_t1 = TR_19 ;
	7'h2f :
		RG_rl_7_t1 = TR_19 ;
	7'h30 :
		RG_rl_7_t1 = TR_19 ;
	7'h31 :
		RG_rl_7_t1 = TR_19 ;
	7'h32 :
		RG_rl_7_t1 = TR_19 ;
	7'h33 :
		RG_rl_7_t1 = TR_19 ;
	7'h34 :
		RG_rl_7_t1 = TR_19 ;
	7'h35 :
		RG_rl_7_t1 = TR_19 ;
	7'h36 :
		RG_rl_7_t1 = TR_19 ;
	7'h37 :
		RG_rl_7_t1 = TR_19 ;
	7'h38 :
		RG_rl_7_t1 = TR_19 ;
	7'h39 :
		RG_rl_7_t1 = TR_19 ;
	7'h3a :
		RG_rl_7_t1 = TR_19 ;
	7'h3b :
		RG_rl_7_t1 = TR_19 ;
	7'h3c :
		RG_rl_7_t1 = TR_19 ;
	7'h3d :
		RG_rl_7_t1 = TR_19 ;
	7'h3e :
		RG_rl_7_t1 = TR_19 ;
	7'h3f :
		RG_rl_7_t1 = TR_19 ;
	7'h40 :
		RG_rl_7_t1 = TR_19 ;
	7'h41 :
		RG_rl_7_t1 = TR_19 ;
	7'h42 :
		RG_rl_7_t1 = TR_19 ;
	7'h43 :
		RG_rl_7_t1 = TR_19 ;
	7'h44 :
		RG_rl_7_t1 = TR_19 ;
	7'h45 :
		RG_rl_7_t1 = TR_19 ;
	7'h46 :
		RG_rl_7_t1 = TR_19 ;
	7'h47 :
		RG_rl_7_t1 = TR_19 ;
	7'h48 :
		RG_rl_7_t1 = TR_19 ;
	7'h49 :
		RG_rl_7_t1 = TR_19 ;
	7'h4a :
		RG_rl_7_t1 = TR_19 ;
	7'h4b :
		RG_rl_7_t1 = TR_19 ;
	7'h4c :
		RG_rl_7_t1 = TR_19 ;
	7'h4d :
		RG_rl_7_t1 = TR_19 ;
	7'h4e :
		RG_rl_7_t1 = TR_19 ;
	7'h4f :
		RG_rl_7_t1 = TR_19 ;
	7'h50 :
		RG_rl_7_t1 = TR_19 ;
	7'h51 :
		RG_rl_7_t1 = TR_19 ;
	7'h52 :
		RG_rl_7_t1 = TR_19 ;
	7'h53 :
		RG_rl_7_t1 = TR_19 ;
	7'h54 :
		RG_rl_7_t1 = TR_19 ;
	7'h55 :
		RG_rl_7_t1 = TR_19 ;
	7'h56 :
		RG_rl_7_t1 = TR_19 ;
	7'h57 :
		RG_rl_7_t1 = TR_19 ;
	7'h58 :
		RG_rl_7_t1 = TR_19 ;
	7'h59 :
		RG_rl_7_t1 = TR_19 ;
	7'h5a :
		RG_rl_7_t1 = TR_19 ;
	7'h5b :
		RG_rl_7_t1 = TR_19 ;
	7'h5c :
		RG_rl_7_t1 = TR_19 ;
	7'h5d :
		RG_rl_7_t1 = TR_19 ;
	7'h5e :
		RG_rl_7_t1 = TR_19 ;
	7'h5f :
		RG_rl_7_t1 = TR_19 ;
	7'h60 :
		RG_rl_7_t1 = TR_19 ;
	7'h61 :
		RG_rl_7_t1 = TR_19 ;
	7'h62 :
		RG_rl_7_t1 = TR_19 ;
	7'h63 :
		RG_rl_7_t1 = TR_19 ;
	7'h64 :
		RG_rl_7_t1 = TR_19 ;
	7'h65 :
		RG_rl_7_t1 = TR_19 ;
	7'h66 :
		RG_rl_7_t1 = TR_19 ;
	7'h67 :
		RG_rl_7_t1 = TR_19 ;
	7'h68 :
		RG_rl_7_t1 = TR_19 ;
	7'h69 :
		RG_rl_7_t1 = TR_19 ;
	7'h6a :
		RG_rl_7_t1 = TR_19 ;
	7'h6b :
		RG_rl_7_t1 = TR_19 ;
	7'h6c :
		RG_rl_7_t1 = TR_19 ;
	7'h6d :
		RG_rl_7_t1 = TR_19 ;
	7'h6e :
		RG_rl_7_t1 = TR_19 ;
	7'h6f :
		RG_rl_7_t1 = TR_19 ;
	7'h70 :
		RG_rl_7_t1 = TR_19 ;
	7'h71 :
		RG_rl_7_t1 = TR_19 ;
	7'h72 :
		RG_rl_7_t1 = TR_19 ;
	7'h73 :
		RG_rl_7_t1 = TR_19 ;
	7'h74 :
		RG_rl_7_t1 = TR_19 ;
	7'h75 :
		RG_rl_7_t1 = TR_19 ;
	7'h76 :
		RG_rl_7_t1 = TR_19 ;
	7'h77 :
		RG_rl_7_t1 = TR_19 ;
	7'h78 :
		RG_rl_7_t1 = TR_19 ;
	7'h79 :
		RG_rl_7_t1 = TR_19 ;
	7'h7a :
		RG_rl_7_t1 = TR_19 ;
	7'h7b :
		RG_rl_7_t1 = TR_19 ;
	7'h7c :
		RG_rl_7_t1 = TR_19 ;
	7'h7d :
		RG_rl_7_t1 = TR_19 ;
	7'h7e :
		RG_rl_7_t1 = TR_19 ;
	7'h7f :
		RG_rl_7_t1 = TR_19 ;
	default :
		RG_rl_7_t1 = 9'hx ;
	endcase
always @ ( RG_rl_7_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_190 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_7_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h07 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_7_t = ( ( { 9{ U_570 } } & RG_rl_190 )
		| ( { 9{ U_569 } } & RG_rl_7_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_7_en = ( U_570 | RG_rl_7_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_7_en )
		RG_rl_7 <= RG_rl_7_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_20 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_8_t1 = TR_20 ;
	7'h01 :
		RG_rl_8_t1 = TR_20 ;
	7'h02 :
		RG_rl_8_t1 = TR_20 ;
	7'h03 :
		RG_rl_8_t1 = TR_20 ;
	7'h04 :
		RG_rl_8_t1 = TR_20 ;
	7'h05 :
		RG_rl_8_t1 = TR_20 ;
	7'h06 :
		RG_rl_8_t1 = TR_20 ;
	7'h07 :
		RG_rl_8_t1 = TR_20 ;
	7'h08 :
		RG_rl_8_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h09 :
		RG_rl_8_t1 = TR_20 ;
	7'h0a :
		RG_rl_8_t1 = TR_20 ;
	7'h0b :
		RG_rl_8_t1 = TR_20 ;
	7'h0c :
		RG_rl_8_t1 = TR_20 ;
	7'h0d :
		RG_rl_8_t1 = TR_20 ;
	7'h0e :
		RG_rl_8_t1 = TR_20 ;
	7'h0f :
		RG_rl_8_t1 = TR_20 ;
	7'h10 :
		RG_rl_8_t1 = TR_20 ;
	7'h11 :
		RG_rl_8_t1 = TR_20 ;
	7'h12 :
		RG_rl_8_t1 = TR_20 ;
	7'h13 :
		RG_rl_8_t1 = TR_20 ;
	7'h14 :
		RG_rl_8_t1 = TR_20 ;
	7'h15 :
		RG_rl_8_t1 = TR_20 ;
	7'h16 :
		RG_rl_8_t1 = TR_20 ;
	7'h17 :
		RG_rl_8_t1 = TR_20 ;
	7'h18 :
		RG_rl_8_t1 = TR_20 ;
	7'h19 :
		RG_rl_8_t1 = TR_20 ;
	7'h1a :
		RG_rl_8_t1 = TR_20 ;
	7'h1b :
		RG_rl_8_t1 = TR_20 ;
	7'h1c :
		RG_rl_8_t1 = TR_20 ;
	7'h1d :
		RG_rl_8_t1 = TR_20 ;
	7'h1e :
		RG_rl_8_t1 = TR_20 ;
	7'h1f :
		RG_rl_8_t1 = TR_20 ;
	7'h20 :
		RG_rl_8_t1 = TR_20 ;
	7'h21 :
		RG_rl_8_t1 = TR_20 ;
	7'h22 :
		RG_rl_8_t1 = TR_20 ;
	7'h23 :
		RG_rl_8_t1 = TR_20 ;
	7'h24 :
		RG_rl_8_t1 = TR_20 ;
	7'h25 :
		RG_rl_8_t1 = TR_20 ;
	7'h26 :
		RG_rl_8_t1 = TR_20 ;
	7'h27 :
		RG_rl_8_t1 = TR_20 ;
	7'h28 :
		RG_rl_8_t1 = TR_20 ;
	7'h29 :
		RG_rl_8_t1 = TR_20 ;
	7'h2a :
		RG_rl_8_t1 = TR_20 ;
	7'h2b :
		RG_rl_8_t1 = TR_20 ;
	7'h2c :
		RG_rl_8_t1 = TR_20 ;
	7'h2d :
		RG_rl_8_t1 = TR_20 ;
	7'h2e :
		RG_rl_8_t1 = TR_20 ;
	7'h2f :
		RG_rl_8_t1 = TR_20 ;
	7'h30 :
		RG_rl_8_t1 = TR_20 ;
	7'h31 :
		RG_rl_8_t1 = TR_20 ;
	7'h32 :
		RG_rl_8_t1 = TR_20 ;
	7'h33 :
		RG_rl_8_t1 = TR_20 ;
	7'h34 :
		RG_rl_8_t1 = TR_20 ;
	7'h35 :
		RG_rl_8_t1 = TR_20 ;
	7'h36 :
		RG_rl_8_t1 = TR_20 ;
	7'h37 :
		RG_rl_8_t1 = TR_20 ;
	7'h38 :
		RG_rl_8_t1 = TR_20 ;
	7'h39 :
		RG_rl_8_t1 = TR_20 ;
	7'h3a :
		RG_rl_8_t1 = TR_20 ;
	7'h3b :
		RG_rl_8_t1 = TR_20 ;
	7'h3c :
		RG_rl_8_t1 = TR_20 ;
	7'h3d :
		RG_rl_8_t1 = TR_20 ;
	7'h3e :
		RG_rl_8_t1 = TR_20 ;
	7'h3f :
		RG_rl_8_t1 = TR_20 ;
	7'h40 :
		RG_rl_8_t1 = TR_20 ;
	7'h41 :
		RG_rl_8_t1 = TR_20 ;
	7'h42 :
		RG_rl_8_t1 = TR_20 ;
	7'h43 :
		RG_rl_8_t1 = TR_20 ;
	7'h44 :
		RG_rl_8_t1 = TR_20 ;
	7'h45 :
		RG_rl_8_t1 = TR_20 ;
	7'h46 :
		RG_rl_8_t1 = TR_20 ;
	7'h47 :
		RG_rl_8_t1 = TR_20 ;
	7'h48 :
		RG_rl_8_t1 = TR_20 ;
	7'h49 :
		RG_rl_8_t1 = TR_20 ;
	7'h4a :
		RG_rl_8_t1 = TR_20 ;
	7'h4b :
		RG_rl_8_t1 = TR_20 ;
	7'h4c :
		RG_rl_8_t1 = TR_20 ;
	7'h4d :
		RG_rl_8_t1 = TR_20 ;
	7'h4e :
		RG_rl_8_t1 = TR_20 ;
	7'h4f :
		RG_rl_8_t1 = TR_20 ;
	7'h50 :
		RG_rl_8_t1 = TR_20 ;
	7'h51 :
		RG_rl_8_t1 = TR_20 ;
	7'h52 :
		RG_rl_8_t1 = TR_20 ;
	7'h53 :
		RG_rl_8_t1 = TR_20 ;
	7'h54 :
		RG_rl_8_t1 = TR_20 ;
	7'h55 :
		RG_rl_8_t1 = TR_20 ;
	7'h56 :
		RG_rl_8_t1 = TR_20 ;
	7'h57 :
		RG_rl_8_t1 = TR_20 ;
	7'h58 :
		RG_rl_8_t1 = TR_20 ;
	7'h59 :
		RG_rl_8_t1 = TR_20 ;
	7'h5a :
		RG_rl_8_t1 = TR_20 ;
	7'h5b :
		RG_rl_8_t1 = TR_20 ;
	7'h5c :
		RG_rl_8_t1 = TR_20 ;
	7'h5d :
		RG_rl_8_t1 = TR_20 ;
	7'h5e :
		RG_rl_8_t1 = TR_20 ;
	7'h5f :
		RG_rl_8_t1 = TR_20 ;
	7'h60 :
		RG_rl_8_t1 = TR_20 ;
	7'h61 :
		RG_rl_8_t1 = TR_20 ;
	7'h62 :
		RG_rl_8_t1 = TR_20 ;
	7'h63 :
		RG_rl_8_t1 = TR_20 ;
	7'h64 :
		RG_rl_8_t1 = TR_20 ;
	7'h65 :
		RG_rl_8_t1 = TR_20 ;
	7'h66 :
		RG_rl_8_t1 = TR_20 ;
	7'h67 :
		RG_rl_8_t1 = TR_20 ;
	7'h68 :
		RG_rl_8_t1 = TR_20 ;
	7'h69 :
		RG_rl_8_t1 = TR_20 ;
	7'h6a :
		RG_rl_8_t1 = TR_20 ;
	7'h6b :
		RG_rl_8_t1 = TR_20 ;
	7'h6c :
		RG_rl_8_t1 = TR_20 ;
	7'h6d :
		RG_rl_8_t1 = TR_20 ;
	7'h6e :
		RG_rl_8_t1 = TR_20 ;
	7'h6f :
		RG_rl_8_t1 = TR_20 ;
	7'h70 :
		RG_rl_8_t1 = TR_20 ;
	7'h71 :
		RG_rl_8_t1 = TR_20 ;
	7'h72 :
		RG_rl_8_t1 = TR_20 ;
	7'h73 :
		RG_rl_8_t1 = TR_20 ;
	7'h74 :
		RG_rl_8_t1 = TR_20 ;
	7'h75 :
		RG_rl_8_t1 = TR_20 ;
	7'h76 :
		RG_rl_8_t1 = TR_20 ;
	7'h77 :
		RG_rl_8_t1 = TR_20 ;
	7'h78 :
		RG_rl_8_t1 = TR_20 ;
	7'h79 :
		RG_rl_8_t1 = TR_20 ;
	7'h7a :
		RG_rl_8_t1 = TR_20 ;
	7'h7b :
		RG_rl_8_t1 = TR_20 ;
	7'h7c :
		RG_rl_8_t1 = TR_20 ;
	7'h7d :
		RG_rl_8_t1 = TR_20 ;
	7'h7e :
		RG_rl_8_t1 = TR_20 ;
	7'h7f :
		RG_rl_8_t1 = TR_20 ;
	default :
		RG_rl_8_t1 = 9'hx ;
	endcase
always @ ( RG_rl_8_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_191 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_8_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h08 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_8_t = ( ( { 9{ U_570 } } & RG_rl_191 )
		| ( { 9{ U_569 } } & RG_rl_8_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_8_en = ( U_570 | RG_rl_8_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_8_en )
		RG_rl_8 <= RG_rl_8_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_21 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_9_t1 = TR_21 ;
	7'h01 :
		RG_rl_9_t1 = TR_21 ;
	7'h02 :
		RG_rl_9_t1 = TR_21 ;
	7'h03 :
		RG_rl_9_t1 = TR_21 ;
	7'h04 :
		RG_rl_9_t1 = TR_21 ;
	7'h05 :
		RG_rl_9_t1 = TR_21 ;
	7'h06 :
		RG_rl_9_t1 = TR_21 ;
	7'h07 :
		RG_rl_9_t1 = TR_21 ;
	7'h08 :
		RG_rl_9_t1 = TR_21 ;
	7'h09 :
		RG_rl_9_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0a :
		RG_rl_9_t1 = TR_21 ;
	7'h0b :
		RG_rl_9_t1 = TR_21 ;
	7'h0c :
		RG_rl_9_t1 = TR_21 ;
	7'h0d :
		RG_rl_9_t1 = TR_21 ;
	7'h0e :
		RG_rl_9_t1 = TR_21 ;
	7'h0f :
		RG_rl_9_t1 = TR_21 ;
	7'h10 :
		RG_rl_9_t1 = TR_21 ;
	7'h11 :
		RG_rl_9_t1 = TR_21 ;
	7'h12 :
		RG_rl_9_t1 = TR_21 ;
	7'h13 :
		RG_rl_9_t1 = TR_21 ;
	7'h14 :
		RG_rl_9_t1 = TR_21 ;
	7'h15 :
		RG_rl_9_t1 = TR_21 ;
	7'h16 :
		RG_rl_9_t1 = TR_21 ;
	7'h17 :
		RG_rl_9_t1 = TR_21 ;
	7'h18 :
		RG_rl_9_t1 = TR_21 ;
	7'h19 :
		RG_rl_9_t1 = TR_21 ;
	7'h1a :
		RG_rl_9_t1 = TR_21 ;
	7'h1b :
		RG_rl_9_t1 = TR_21 ;
	7'h1c :
		RG_rl_9_t1 = TR_21 ;
	7'h1d :
		RG_rl_9_t1 = TR_21 ;
	7'h1e :
		RG_rl_9_t1 = TR_21 ;
	7'h1f :
		RG_rl_9_t1 = TR_21 ;
	7'h20 :
		RG_rl_9_t1 = TR_21 ;
	7'h21 :
		RG_rl_9_t1 = TR_21 ;
	7'h22 :
		RG_rl_9_t1 = TR_21 ;
	7'h23 :
		RG_rl_9_t1 = TR_21 ;
	7'h24 :
		RG_rl_9_t1 = TR_21 ;
	7'h25 :
		RG_rl_9_t1 = TR_21 ;
	7'h26 :
		RG_rl_9_t1 = TR_21 ;
	7'h27 :
		RG_rl_9_t1 = TR_21 ;
	7'h28 :
		RG_rl_9_t1 = TR_21 ;
	7'h29 :
		RG_rl_9_t1 = TR_21 ;
	7'h2a :
		RG_rl_9_t1 = TR_21 ;
	7'h2b :
		RG_rl_9_t1 = TR_21 ;
	7'h2c :
		RG_rl_9_t1 = TR_21 ;
	7'h2d :
		RG_rl_9_t1 = TR_21 ;
	7'h2e :
		RG_rl_9_t1 = TR_21 ;
	7'h2f :
		RG_rl_9_t1 = TR_21 ;
	7'h30 :
		RG_rl_9_t1 = TR_21 ;
	7'h31 :
		RG_rl_9_t1 = TR_21 ;
	7'h32 :
		RG_rl_9_t1 = TR_21 ;
	7'h33 :
		RG_rl_9_t1 = TR_21 ;
	7'h34 :
		RG_rl_9_t1 = TR_21 ;
	7'h35 :
		RG_rl_9_t1 = TR_21 ;
	7'h36 :
		RG_rl_9_t1 = TR_21 ;
	7'h37 :
		RG_rl_9_t1 = TR_21 ;
	7'h38 :
		RG_rl_9_t1 = TR_21 ;
	7'h39 :
		RG_rl_9_t1 = TR_21 ;
	7'h3a :
		RG_rl_9_t1 = TR_21 ;
	7'h3b :
		RG_rl_9_t1 = TR_21 ;
	7'h3c :
		RG_rl_9_t1 = TR_21 ;
	7'h3d :
		RG_rl_9_t1 = TR_21 ;
	7'h3e :
		RG_rl_9_t1 = TR_21 ;
	7'h3f :
		RG_rl_9_t1 = TR_21 ;
	7'h40 :
		RG_rl_9_t1 = TR_21 ;
	7'h41 :
		RG_rl_9_t1 = TR_21 ;
	7'h42 :
		RG_rl_9_t1 = TR_21 ;
	7'h43 :
		RG_rl_9_t1 = TR_21 ;
	7'h44 :
		RG_rl_9_t1 = TR_21 ;
	7'h45 :
		RG_rl_9_t1 = TR_21 ;
	7'h46 :
		RG_rl_9_t1 = TR_21 ;
	7'h47 :
		RG_rl_9_t1 = TR_21 ;
	7'h48 :
		RG_rl_9_t1 = TR_21 ;
	7'h49 :
		RG_rl_9_t1 = TR_21 ;
	7'h4a :
		RG_rl_9_t1 = TR_21 ;
	7'h4b :
		RG_rl_9_t1 = TR_21 ;
	7'h4c :
		RG_rl_9_t1 = TR_21 ;
	7'h4d :
		RG_rl_9_t1 = TR_21 ;
	7'h4e :
		RG_rl_9_t1 = TR_21 ;
	7'h4f :
		RG_rl_9_t1 = TR_21 ;
	7'h50 :
		RG_rl_9_t1 = TR_21 ;
	7'h51 :
		RG_rl_9_t1 = TR_21 ;
	7'h52 :
		RG_rl_9_t1 = TR_21 ;
	7'h53 :
		RG_rl_9_t1 = TR_21 ;
	7'h54 :
		RG_rl_9_t1 = TR_21 ;
	7'h55 :
		RG_rl_9_t1 = TR_21 ;
	7'h56 :
		RG_rl_9_t1 = TR_21 ;
	7'h57 :
		RG_rl_9_t1 = TR_21 ;
	7'h58 :
		RG_rl_9_t1 = TR_21 ;
	7'h59 :
		RG_rl_9_t1 = TR_21 ;
	7'h5a :
		RG_rl_9_t1 = TR_21 ;
	7'h5b :
		RG_rl_9_t1 = TR_21 ;
	7'h5c :
		RG_rl_9_t1 = TR_21 ;
	7'h5d :
		RG_rl_9_t1 = TR_21 ;
	7'h5e :
		RG_rl_9_t1 = TR_21 ;
	7'h5f :
		RG_rl_9_t1 = TR_21 ;
	7'h60 :
		RG_rl_9_t1 = TR_21 ;
	7'h61 :
		RG_rl_9_t1 = TR_21 ;
	7'h62 :
		RG_rl_9_t1 = TR_21 ;
	7'h63 :
		RG_rl_9_t1 = TR_21 ;
	7'h64 :
		RG_rl_9_t1 = TR_21 ;
	7'h65 :
		RG_rl_9_t1 = TR_21 ;
	7'h66 :
		RG_rl_9_t1 = TR_21 ;
	7'h67 :
		RG_rl_9_t1 = TR_21 ;
	7'h68 :
		RG_rl_9_t1 = TR_21 ;
	7'h69 :
		RG_rl_9_t1 = TR_21 ;
	7'h6a :
		RG_rl_9_t1 = TR_21 ;
	7'h6b :
		RG_rl_9_t1 = TR_21 ;
	7'h6c :
		RG_rl_9_t1 = TR_21 ;
	7'h6d :
		RG_rl_9_t1 = TR_21 ;
	7'h6e :
		RG_rl_9_t1 = TR_21 ;
	7'h6f :
		RG_rl_9_t1 = TR_21 ;
	7'h70 :
		RG_rl_9_t1 = TR_21 ;
	7'h71 :
		RG_rl_9_t1 = TR_21 ;
	7'h72 :
		RG_rl_9_t1 = TR_21 ;
	7'h73 :
		RG_rl_9_t1 = TR_21 ;
	7'h74 :
		RG_rl_9_t1 = TR_21 ;
	7'h75 :
		RG_rl_9_t1 = TR_21 ;
	7'h76 :
		RG_rl_9_t1 = TR_21 ;
	7'h77 :
		RG_rl_9_t1 = TR_21 ;
	7'h78 :
		RG_rl_9_t1 = TR_21 ;
	7'h79 :
		RG_rl_9_t1 = TR_21 ;
	7'h7a :
		RG_rl_9_t1 = TR_21 ;
	7'h7b :
		RG_rl_9_t1 = TR_21 ;
	7'h7c :
		RG_rl_9_t1 = TR_21 ;
	7'h7d :
		RG_rl_9_t1 = TR_21 ;
	7'h7e :
		RG_rl_9_t1 = TR_21 ;
	7'h7f :
		RG_rl_9_t1 = TR_21 ;
	default :
		RG_rl_9_t1 = 9'hx ;
	endcase
always @ ( RG_rl_9_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_192 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_9_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h09 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_9_t = ( ( { 9{ U_570 } } & RG_rl_192 )
		| ( { 9{ U_569 } } & RG_rl_9_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_9_en = ( U_570 | RG_rl_9_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_9_en )
		RG_rl_9 <= RG_rl_9_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_22 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_10_t1 = TR_22 ;
	7'h01 :
		RG_rl_10_t1 = TR_22 ;
	7'h02 :
		RG_rl_10_t1 = TR_22 ;
	7'h03 :
		RG_rl_10_t1 = TR_22 ;
	7'h04 :
		RG_rl_10_t1 = TR_22 ;
	7'h05 :
		RG_rl_10_t1 = TR_22 ;
	7'h06 :
		RG_rl_10_t1 = TR_22 ;
	7'h07 :
		RG_rl_10_t1 = TR_22 ;
	7'h08 :
		RG_rl_10_t1 = TR_22 ;
	7'h09 :
		RG_rl_10_t1 = TR_22 ;
	7'h0a :
		RG_rl_10_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0b :
		RG_rl_10_t1 = TR_22 ;
	7'h0c :
		RG_rl_10_t1 = TR_22 ;
	7'h0d :
		RG_rl_10_t1 = TR_22 ;
	7'h0e :
		RG_rl_10_t1 = TR_22 ;
	7'h0f :
		RG_rl_10_t1 = TR_22 ;
	7'h10 :
		RG_rl_10_t1 = TR_22 ;
	7'h11 :
		RG_rl_10_t1 = TR_22 ;
	7'h12 :
		RG_rl_10_t1 = TR_22 ;
	7'h13 :
		RG_rl_10_t1 = TR_22 ;
	7'h14 :
		RG_rl_10_t1 = TR_22 ;
	7'h15 :
		RG_rl_10_t1 = TR_22 ;
	7'h16 :
		RG_rl_10_t1 = TR_22 ;
	7'h17 :
		RG_rl_10_t1 = TR_22 ;
	7'h18 :
		RG_rl_10_t1 = TR_22 ;
	7'h19 :
		RG_rl_10_t1 = TR_22 ;
	7'h1a :
		RG_rl_10_t1 = TR_22 ;
	7'h1b :
		RG_rl_10_t1 = TR_22 ;
	7'h1c :
		RG_rl_10_t1 = TR_22 ;
	7'h1d :
		RG_rl_10_t1 = TR_22 ;
	7'h1e :
		RG_rl_10_t1 = TR_22 ;
	7'h1f :
		RG_rl_10_t1 = TR_22 ;
	7'h20 :
		RG_rl_10_t1 = TR_22 ;
	7'h21 :
		RG_rl_10_t1 = TR_22 ;
	7'h22 :
		RG_rl_10_t1 = TR_22 ;
	7'h23 :
		RG_rl_10_t1 = TR_22 ;
	7'h24 :
		RG_rl_10_t1 = TR_22 ;
	7'h25 :
		RG_rl_10_t1 = TR_22 ;
	7'h26 :
		RG_rl_10_t1 = TR_22 ;
	7'h27 :
		RG_rl_10_t1 = TR_22 ;
	7'h28 :
		RG_rl_10_t1 = TR_22 ;
	7'h29 :
		RG_rl_10_t1 = TR_22 ;
	7'h2a :
		RG_rl_10_t1 = TR_22 ;
	7'h2b :
		RG_rl_10_t1 = TR_22 ;
	7'h2c :
		RG_rl_10_t1 = TR_22 ;
	7'h2d :
		RG_rl_10_t1 = TR_22 ;
	7'h2e :
		RG_rl_10_t1 = TR_22 ;
	7'h2f :
		RG_rl_10_t1 = TR_22 ;
	7'h30 :
		RG_rl_10_t1 = TR_22 ;
	7'h31 :
		RG_rl_10_t1 = TR_22 ;
	7'h32 :
		RG_rl_10_t1 = TR_22 ;
	7'h33 :
		RG_rl_10_t1 = TR_22 ;
	7'h34 :
		RG_rl_10_t1 = TR_22 ;
	7'h35 :
		RG_rl_10_t1 = TR_22 ;
	7'h36 :
		RG_rl_10_t1 = TR_22 ;
	7'h37 :
		RG_rl_10_t1 = TR_22 ;
	7'h38 :
		RG_rl_10_t1 = TR_22 ;
	7'h39 :
		RG_rl_10_t1 = TR_22 ;
	7'h3a :
		RG_rl_10_t1 = TR_22 ;
	7'h3b :
		RG_rl_10_t1 = TR_22 ;
	7'h3c :
		RG_rl_10_t1 = TR_22 ;
	7'h3d :
		RG_rl_10_t1 = TR_22 ;
	7'h3e :
		RG_rl_10_t1 = TR_22 ;
	7'h3f :
		RG_rl_10_t1 = TR_22 ;
	7'h40 :
		RG_rl_10_t1 = TR_22 ;
	7'h41 :
		RG_rl_10_t1 = TR_22 ;
	7'h42 :
		RG_rl_10_t1 = TR_22 ;
	7'h43 :
		RG_rl_10_t1 = TR_22 ;
	7'h44 :
		RG_rl_10_t1 = TR_22 ;
	7'h45 :
		RG_rl_10_t1 = TR_22 ;
	7'h46 :
		RG_rl_10_t1 = TR_22 ;
	7'h47 :
		RG_rl_10_t1 = TR_22 ;
	7'h48 :
		RG_rl_10_t1 = TR_22 ;
	7'h49 :
		RG_rl_10_t1 = TR_22 ;
	7'h4a :
		RG_rl_10_t1 = TR_22 ;
	7'h4b :
		RG_rl_10_t1 = TR_22 ;
	7'h4c :
		RG_rl_10_t1 = TR_22 ;
	7'h4d :
		RG_rl_10_t1 = TR_22 ;
	7'h4e :
		RG_rl_10_t1 = TR_22 ;
	7'h4f :
		RG_rl_10_t1 = TR_22 ;
	7'h50 :
		RG_rl_10_t1 = TR_22 ;
	7'h51 :
		RG_rl_10_t1 = TR_22 ;
	7'h52 :
		RG_rl_10_t1 = TR_22 ;
	7'h53 :
		RG_rl_10_t1 = TR_22 ;
	7'h54 :
		RG_rl_10_t1 = TR_22 ;
	7'h55 :
		RG_rl_10_t1 = TR_22 ;
	7'h56 :
		RG_rl_10_t1 = TR_22 ;
	7'h57 :
		RG_rl_10_t1 = TR_22 ;
	7'h58 :
		RG_rl_10_t1 = TR_22 ;
	7'h59 :
		RG_rl_10_t1 = TR_22 ;
	7'h5a :
		RG_rl_10_t1 = TR_22 ;
	7'h5b :
		RG_rl_10_t1 = TR_22 ;
	7'h5c :
		RG_rl_10_t1 = TR_22 ;
	7'h5d :
		RG_rl_10_t1 = TR_22 ;
	7'h5e :
		RG_rl_10_t1 = TR_22 ;
	7'h5f :
		RG_rl_10_t1 = TR_22 ;
	7'h60 :
		RG_rl_10_t1 = TR_22 ;
	7'h61 :
		RG_rl_10_t1 = TR_22 ;
	7'h62 :
		RG_rl_10_t1 = TR_22 ;
	7'h63 :
		RG_rl_10_t1 = TR_22 ;
	7'h64 :
		RG_rl_10_t1 = TR_22 ;
	7'h65 :
		RG_rl_10_t1 = TR_22 ;
	7'h66 :
		RG_rl_10_t1 = TR_22 ;
	7'h67 :
		RG_rl_10_t1 = TR_22 ;
	7'h68 :
		RG_rl_10_t1 = TR_22 ;
	7'h69 :
		RG_rl_10_t1 = TR_22 ;
	7'h6a :
		RG_rl_10_t1 = TR_22 ;
	7'h6b :
		RG_rl_10_t1 = TR_22 ;
	7'h6c :
		RG_rl_10_t1 = TR_22 ;
	7'h6d :
		RG_rl_10_t1 = TR_22 ;
	7'h6e :
		RG_rl_10_t1 = TR_22 ;
	7'h6f :
		RG_rl_10_t1 = TR_22 ;
	7'h70 :
		RG_rl_10_t1 = TR_22 ;
	7'h71 :
		RG_rl_10_t1 = TR_22 ;
	7'h72 :
		RG_rl_10_t1 = TR_22 ;
	7'h73 :
		RG_rl_10_t1 = TR_22 ;
	7'h74 :
		RG_rl_10_t1 = TR_22 ;
	7'h75 :
		RG_rl_10_t1 = TR_22 ;
	7'h76 :
		RG_rl_10_t1 = TR_22 ;
	7'h77 :
		RG_rl_10_t1 = TR_22 ;
	7'h78 :
		RG_rl_10_t1 = TR_22 ;
	7'h79 :
		RG_rl_10_t1 = TR_22 ;
	7'h7a :
		RG_rl_10_t1 = TR_22 ;
	7'h7b :
		RG_rl_10_t1 = TR_22 ;
	7'h7c :
		RG_rl_10_t1 = TR_22 ;
	7'h7d :
		RG_rl_10_t1 = TR_22 ;
	7'h7e :
		RG_rl_10_t1 = TR_22 ;
	7'h7f :
		RG_rl_10_t1 = TR_22 ;
	default :
		RG_rl_10_t1 = 9'hx ;
	endcase
always @ ( RG_rl_10_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_193 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_10_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h0a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_10_t = ( ( { 9{ U_570 } } & RG_rl_193 )
		| ( { 9{ U_569 } } & RG_rl_10_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_10_en = ( U_570 | RG_rl_10_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_10_en )
		RG_rl_10 <= RG_rl_10_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_23 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_11_t1 = TR_23 ;
	7'h01 :
		RG_rl_11_t1 = TR_23 ;
	7'h02 :
		RG_rl_11_t1 = TR_23 ;
	7'h03 :
		RG_rl_11_t1 = TR_23 ;
	7'h04 :
		RG_rl_11_t1 = TR_23 ;
	7'h05 :
		RG_rl_11_t1 = TR_23 ;
	7'h06 :
		RG_rl_11_t1 = TR_23 ;
	7'h07 :
		RG_rl_11_t1 = TR_23 ;
	7'h08 :
		RG_rl_11_t1 = TR_23 ;
	7'h09 :
		RG_rl_11_t1 = TR_23 ;
	7'h0a :
		RG_rl_11_t1 = TR_23 ;
	7'h0b :
		RG_rl_11_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0c :
		RG_rl_11_t1 = TR_23 ;
	7'h0d :
		RG_rl_11_t1 = TR_23 ;
	7'h0e :
		RG_rl_11_t1 = TR_23 ;
	7'h0f :
		RG_rl_11_t1 = TR_23 ;
	7'h10 :
		RG_rl_11_t1 = TR_23 ;
	7'h11 :
		RG_rl_11_t1 = TR_23 ;
	7'h12 :
		RG_rl_11_t1 = TR_23 ;
	7'h13 :
		RG_rl_11_t1 = TR_23 ;
	7'h14 :
		RG_rl_11_t1 = TR_23 ;
	7'h15 :
		RG_rl_11_t1 = TR_23 ;
	7'h16 :
		RG_rl_11_t1 = TR_23 ;
	7'h17 :
		RG_rl_11_t1 = TR_23 ;
	7'h18 :
		RG_rl_11_t1 = TR_23 ;
	7'h19 :
		RG_rl_11_t1 = TR_23 ;
	7'h1a :
		RG_rl_11_t1 = TR_23 ;
	7'h1b :
		RG_rl_11_t1 = TR_23 ;
	7'h1c :
		RG_rl_11_t1 = TR_23 ;
	7'h1d :
		RG_rl_11_t1 = TR_23 ;
	7'h1e :
		RG_rl_11_t1 = TR_23 ;
	7'h1f :
		RG_rl_11_t1 = TR_23 ;
	7'h20 :
		RG_rl_11_t1 = TR_23 ;
	7'h21 :
		RG_rl_11_t1 = TR_23 ;
	7'h22 :
		RG_rl_11_t1 = TR_23 ;
	7'h23 :
		RG_rl_11_t1 = TR_23 ;
	7'h24 :
		RG_rl_11_t1 = TR_23 ;
	7'h25 :
		RG_rl_11_t1 = TR_23 ;
	7'h26 :
		RG_rl_11_t1 = TR_23 ;
	7'h27 :
		RG_rl_11_t1 = TR_23 ;
	7'h28 :
		RG_rl_11_t1 = TR_23 ;
	7'h29 :
		RG_rl_11_t1 = TR_23 ;
	7'h2a :
		RG_rl_11_t1 = TR_23 ;
	7'h2b :
		RG_rl_11_t1 = TR_23 ;
	7'h2c :
		RG_rl_11_t1 = TR_23 ;
	7'h2d :
		RG_rl_11_t1 = TR_23 ;
	7'h2e :
		RG_rl_11_t1 = TR_23 ;
	7'h2f :
		RG_rl_11_t1 = TR_23 ;
	7'h30 :
		RG_rl_11_t1 = TR_23 ;
	7'h31 :
		RG_rl_11_t1 = TR_23 ;
	7'h32 :
		RG_rl_11_t1 = TR_23 ;
	7'h33 :
		RG_rl_11_t1 = TR_23 ;
	7'h34 :
		RG_rl_11_t1 = TR_23 ;
	7'h35 :
		RG_rl_11_t1 = TR_23 ;
	7'h36 :
		RG_rl_11_t1 = TR_23 ;
	7'h37 :
		RG_rl_11_t1 = TR_23 ;
	7'h38 :
		RG_rl_11_t1 = TR_23 ;
	7'h39 :
		RG_rl_11_t1 = TR_23 ;
	7'h3a :
		RG_rl_11_t1 = TR_23 ;
	7'h3b :
		RG_rl_11_t1 = TR_23 ;
	7'h3c :
		RG_rl_11_t1 = TR_23 ;
	7'h3d :
		RG_rl_11_t1 = TR_23 ;
	7'h3e :
		RG_rl_11_t1 = TR_23 ;
	7'h3f :
		RG_rl_11_t1 = TR_23 ;
	7'h40 :
		RG_rl_11_t1 = TR_23 ;
	7'h41 :
		RG_rl_11_t1 = TR_23 ;
	7'h42 :
		RG_rl_11_t1 = TR_23 ;
	7'h43 :
		RG_rl_11_t1 = TR_23 ;
	7'h44 :
		RG_rl_11_t1 = TR_23 ;
	7'h45 :
		RG_rl_11_t1 = TR_23 ;
	7'h46 :
		RG_rl_11_t1 = TR_23 ;
	7'h47 :
		RG_rl_11_t1 = TR_23 ;
	7'h48 :
		RG_rl_11_t1 = TR_23 ;
	7'h49 :
		RG_rl_11_t1 = TR_23 ;
	7'h4a :
		RG_rl_11_t1 = TR_23 ;
	7'h4b :
		RG_rl_11_t1 = TR_23 ;
	7'h4c :
		RG_rl_11_t1 = TR_23 ;
	7'h4d :
		RG_rl_11_t1 = TR_23 ;
	7'h4e :
		RG_rl_11_t1 = TR_23 ;
	7'h4f :
		RG_rl_11_t1 = TR_23 ;
	7'h50 :
		RG_rl_11_t1 = TR_23 ;
	7'h51 :
		RG_rl_11_t1 = TR_23 ;
	7'h52 :
		RG_rl_11_t1 = TR_23 ;
	7'h53 :
		RG_rl_11_t1 = TR_23 ;
	7'h54 :
		RG_rl_11_t1 = TR_23 ;
	7'h55 :
		RG_rl_11_t1 = TR_23 ;
	7'h56 :
		RG_rl_11_t1 = TR_23 ;
	7'h57 :
		RG_rl_11_t1 = TR_23 ;
	7'h58 :
		RG_rl_11_t1 = TR_23 ;
	7'h59 :
		RG_rl_11_t1 = TR_23 ;
	7'h5a :
		RG_rl_11_t1 = TR_23 ;
	7'h5b :
		RG_rl_11_t1 = TR_23 ;
	7'h5c :
		RG_rl_11_t1 = TR_23 ;
	7'h5d :
		RG_rl_11_t1 = TR_23 ;
	7'h5e :
		RG_rl_11_t1 = TR_23 ;
	7'h5f :
		RG_rl_11_t1 = TR_23 ;
	7'h60 :
		RG_rl_11_t1 = TR_23 ;
	7'h61 :
		RG_rl_11_t1 = TR_23 ;
	7'h62 :
		RG_rl_11_t1 = TR_23 ;
	7'h63 :
		RG_rl_11_t1 = TR_23 ;
	7'h64 :
		RG_rl_11_t1 = TR_23 ;
	7'h65 :
		RG_rl_11_t1 = TR_23 ;
	7'h66 :
		RG_rl_11_t1 = TR_23 ;
	7'h67 :
		RG_rl_11_t1 = TR_23 ;
	7'h68 :
		RG_rl_11_t1 = TR_23 ;
	7'h69 :
		RG_rl_11_t1 = TR_23 ;
	7'h6a :
		RG_rl_11_t1 = TR_23 ;
	7'h6b :
		RG_rl_11_t1 = TR_23 ;
	7'h6c :
		RG_rl_11_t1 = TR_23 ;
	7'h6d :
		RG_rl_11_t1 = TR_23 ;
	7'h6e :
		RG_rl_11_t1 = TR_23 ;
	7'h6f :
		RG_rl_11_t1 = TR_23 ;
	7'h70 :
		RG_rl_11_t1 = TR_23 ;
	7'h71 :
		RG_rl_11_t1 = TR_23 ;
	7'h72 :
		RG_rl_11_t1 = TR_23 ;
	7'h73 :
		RG_rl_11_t1 = TR_23 ;
	7'h74 :
		RG_rl_11_t1 = TR_23 ;
	7'h75 :
		RG_rl_11_t1 = TR_23 ;
	7'h76 :
		RG_rl_11_t1 = TR_23 ;
	7'h77 :
		RG_rl_11_t1 = TR_23 ;
	7'h78 :
		RG_rl_11_t1 = TR_23 ;
	7'h79 :
		RG_rl_11_t1 = TR_23 ;
	7'h7a :
		RG_rl_11_t1 = TR_23 ;
	7'h7b :
		RG_rl_11_t1 = TR_23 ;
	7'h7c :
		RG_rl_11_t1 = TR_23 ;
	7'h7d :
		RG_rl_11_t1 = TR_23 ;
	7'h7e :
		RG_rl_11_t1 = TR_23 ;
	7'h7f :
		RG_rl_11_t1 = TR_23 ;
	default :
		RG_rl_11_t1 = 9'hx ;
	endcase
always @ ( RG_rl_11_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_194 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_11_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h0b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_11_t = ( ( { 9{ U_570 } } & RG_rl_194 )
		| ( { 9{ U_569 } } & RG_rl_11_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_11_en = ( U_570 | RG_rl_11_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_11_en )
		RG_rl_11 <= RG_rl_11_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_24 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_12_t1 = TR_24 ;
	7'h01 :
		RG_rl_12_t1 = TR_24 ;
	7'h02 :
		RG_rl_12_t1 = TR_24 ;
	7'h03 :
		RG_rl_12_t1 = TR_24 ;
	7'h04 :
		RG_rl_12_t1 = TR_24 ;
	7'h05 :
		RG_rl_12_t1 = TR_24 ;
	7'h06 :
		RG_rl_12_t1 = TR_24 ;
	7'h07 :
		RG_rl_12_t1 = TR_24 ;
	7'h08 :
		RG_rl_12_t1 = TR_24 ;
	7'h09 :
		RG_rl_12_t1 = TR_24 ;
	7'h0a :
		RG_rl_12_t1 = TR_24 ;
	7'h0b :
		RG_rl_12_t1 = TR_24 ;
	7'h0c :
		RG_rl_12_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0d :
		RG_rl_12_t1 = TR_24 ;
	7'h0e :
		RG_rl_12_t1 = TR_24 ;
	7'h0f :
		RG_rl_12_t1 = TR_24 ;
	7'h10 :
		RG_rl_12_t1 = TR_24 ;
	7'h11 :
		RG_rl_12_t1 = TR_24 ;
	7'h12 :
		RG_rl_12_t1 = TR_24 ;
	7'h13 :
		RG_rl_12_t1 = TR_24 ;
	7'h14 :
		RG_rl_12_t1 = TR_24 ;
	7'h15 :
		RG_rl_12_t1 = TR_24 ;
	7'h16 :
		RG_rl_12_t1 = TR_24 ;
	7'h17 :
		RG_rl_12_t1 = TR_24 ;
	7'h18 :
		RG_rl_12_t1 = TR_24 ;
	7'h19 :
		RG_rl_12_t1 = TR_24 ;
	7'h1a :
		RG_rl_12_t1 = TR_24 ;
	7'h1b :
		RG_rl_12_t1 = TR_24 ;
	7'h1c :
		RG_rl_12_t1 = TR_24 ;
	7'h1d :
		RG_rl_12_t1 = TR_24 ;
	7'h1e :
		RG_rl_12_t1 = TR_24 ;
	7'h1f :
		RG_rl_12_t1 = TR_24 ;
	7'h20 :
		RG_rl_12_t1 = TR_24 ;
	7'h21 :
		RG_rl_12_t1 = TR_24 ;
	7'h22 :
		RG_rl_12_t1 = TR_24 ;
	7'h23 :
		RG_rl_12_t1 = TR_24 ;
	7'h24 :
		RG_rl_12_t1 = TR_24 ;
	7'h25 :
		RG_rl_12_t1 = TR_24 ;
	7'h26 :
		RG_rl_12_t1 = TR_24 ;
	7'h27 :
		RG_rl_12_t1 = TR_24 ;
	7'h28 :
		RG_rl_12_t1 = TR_24 ;
	7'h29 :
		RG_rl_12_t1 = TR_24 ;
	7'h2a :
		RG_rl_12_t1 = TR_24 ;
	7'h2b :
		RG_rl_12_t1 = TR_24 ;
	7'h2c :
		RG_rl_12_t1 = TR_24 ;
	7'h2d :
		RG_rl_12_t1 = TR_24 ;
	7'h2e :
		RG_rl_12_t1 = TR_24 ;
	7'h2f :
		RG_rl_12_t1 = TR_24 ;
	7'h30 :
		RG_rl_12_t1 = TR_24 ;
	7'h31 :
		RG_rl_12_t1 = TR_24 ;
	7'h32 :
		RG_rl_12_t1 = TR_24 ;
	7'h33 :
		RG_rl_12_t1 = TR_24 ;
	7'h34 :
		RG_rl_12_t1 = TR_24 ;
	7'h35 :
		RG_rl_12_t1 = TR_24 ;
	7'h36 :
		RG_rl_12_t1 = TR_24 ;
	7'h37 :
		RG_rl_12_t1 = TR_24 ;
	7'h38 :
		RG_rl_12_t1 = TR_24 ;
	7'h39 :
		RG_rl_12_t1 = TR_24 ;
	7'h3a :
		RG_rl_12_t1 = TR_24 ;
	7'h3b :
		RG_rl_12_t1 = TR_24 ;
	7'h3c :
		RG_rl_12_t1 = TR_24 ;
	7'h3d :
		RG_rl_12_t1 = TR_24 ;
	7'h3e :
		RG_rl_12_t1 = TR_24 ;
	7'h3f :
		RG_rl_12_t1 = TR_24 ;
	7'h40 :
		RG_rl_12_t1 = TR_24 ;
	7'h41 :
		RG_rl_12_t1 = TR_24 ;
	7'h42 :
		RG_rl_12_t1 = TR_24 ;
	7'h43 :
		RG_rl_12_t1 = TR_24 ;
	7'h44 :
		RG_rl_12_t1 = TR_24 ;
	7'h45 :
		RG_rl_12_t1 = TR_24 ;
	7'h46 :
		RG_rl_12_t1 = TR_24 ;
	7'h47 :
		RG_rl_12_t1 = TR_24 ;
	7'h48 :
		RG_rl_12_t1 = TR_24 ;
	7'h49 :
		RG_rl_12_t1 = TR_24 ;
	7'h4a :
		RG_rl_12_t1 = TR_24 ;
	7'h4b :
		RG_rl_12_t1 = TR_24 ;
	7'h4c :
		RG_rl_12_t1 = TR_24 ;
	7'h4d :
		RG_rl_12_t1 = TR_24 ;
	7'h4e :
		RG_rl_12_t1 = TR_24 ;
	7'h4f :
		RG_rl_12_t1 = TR_24 ;
	7'h50 :
		RG_rl_12_t1 = TR_24 ;
	7'h51 :
		RG_rl_12_t1 = TR_24 ;
	7'h52 :
		RG_rl_12_t1 = TR_24 ;
	7'h53 :
		RG_rl_12_t1 = TR_24 ;
	7'h54 :
		RG_rl_12_t1 = TR_24 ;
	7'h55 :
		RG_rl_12_t1 = TR_24 ;
	7'h56 :
		RG_rl_12_t1 = TR_24 ;
	7'h57 :
		RG_rl_12_t1 = TR_24 ;
	7'h58 :
		RG_rl_12_t1 = TR_24 ;
	7'h59 :
		RG_rl_12_t1 = TR_24 ;
	7'h5a :
		RG_rl_12_t1 = TR_24 ;
	7'h5b :
		RG_rl_12_t1 = TR_24 ;
	7'h5c :
		RG_rl_12_t1 = TR_24 ;
	7'h5d :
		RG_rl_12_t1 = TR_24 ;
	7'h5e :
		RG_rl_12_t1 = TR_24 ;
	7'h5f :
		RG_rl_12_t1 = TR_24 ;
	7'h60 :
		RG_rl_12_t1 = TR_24 ;
	7'h61 :
		RG_rl_12_t1 = TR_24 ;
	7'h62 :
		RG_rl_12_t1 = TR_24 ;
	7'h63 :
		RG_rl_12_t1 = TR_24 ;
	7'h64 :
		RG_rl_12_t1 = TR_24 ;
	7'h65 :
		RG_rl_12_t1 = TR_24 ;
	7'h66 :
		RG_rl_12_t1 = TR_24 ;
	7'h67 :
		RG_rl_12_t1 = TR_24 ;
	7'h68 :
		RG_rl_12_t1 = TR_24 ;
	7'h69 :
		RG_rl_12_t1 = TR_24 ;
	7'h6a :
		RG_rl_12_t1 = TR_24 ;
	7'h6b :
		RG_rl_12_t1 = TR_24 ;
	7'h6c :
		RG_rl_12_t1 = TR_24 ;
	7'h6d :
		RG_rl_12_t1 = TR_24 ;
	7'h6e :
		RG_rl_12_t1 = TR_24 ;
	7'h6f :
		RG_rl_12_t1 = TR_24 ;
	7'h70 :
		RG_rl_12_t1 = TR_24 ;
	7'h71 :
		RG_rl_12_t1 = TR_24 ;
	7'h72 :
		RG_rl_12_t1 = TR_24 ;
	7'h73 :
		RG_rl_12_t1 = TR_24 ;
	7'h74 :
		RG_rl_12_t1 = TR_24 ;
	7'h75 :
		RG_rl_12_t1 = TR_24 ;
	7'h76 :
		RG_rl_12_t1 = TR_24 ;
	7'h77 :
		RG_rl_12_t1 = TR_24 ;
	7'h78 :
		RG_rl_12_t1 = TR_24 ;
	7'h79 :
		RG_rl_12_t1 = TR_24 ;
	7'h7a :
		RG_rl_12_t1 = TR_24 ;
	7'h7b :
		RG_rl_12_t1 = TR_24 ;
	7'h7c :
		RG_rl_12_t1 = TR_24 ;
	7'h7d :
		RG_rl_12_t1 = TR_24 ;
	7'h7e :
		RG_rl_12_t1 = TR_24 ;
	7'h7f :
		RG_rl_12_t1 = TR_24 ;
	default :
		RG_rl_12_t1 = 9'hx ;
	endcase
always @ ( RG_rl_12_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_195 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_12_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h0c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_12_t = ( ( { 9{ U_570 } } & RG_rl_195 )
		| ( { 9{ U_569 } } & RG_rl_12_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_12_en = ( U_570 | RG_rl_12_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_12_en )
		RG_rl_12 <= RG_rl_12_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_25 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_13_t1 = TR_25 ;
	7'h01 :
		RG_rl_13_t1 = TR_25 ;
	7'h02 :
		RG_rl_13_t1 = TR_25 ;
	7'h03 :
		RG_rl_13_t1 = TR_25 ;
	7'h04 :
		RG_rl_13_t1 = TR_25 ;
	7'h05 :
		RG_rl_13_t1 = TR_25 ;
	7'h06 :
		RG_rl_13_t1 = TR_25 ;
	7'h07 :
		RG_rl_13_t1 = TR_25 ;
	7'h08 :
		RG_rl_13_t1 = TR_25 ;
	7'h09 :
		RG_rl_13_t1 = TR_25 ;
	7'h0a :
		RG_rl_13_t1 = TR_25 ;
	7'h0b :
		RG_rl_13_t1 = TR_25 ;
	7'h0c :
		RG_rl_13_t1 = TR_25 ;
	7'h0d :
		RG_rl_13_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0e :
		RG_rl_13_t1 = TR_25 ;
	7'h0f :
		RG_rl_13_t1 = TR_25 ;
	7'h10 :
		RG_rl_13_t1 = TR_25 ;
	7'h11 :
		RG_rl_13_t1 = TR_25 ;
	7'h12 :
		RG_rl_13_t1 = TR_25 ;
	7'h13 :
		RG_rl_13_t1 = TR_25 ;
	7'h14 :
		RG_rl_13_t1 = TR_25 ;
	7'h15 :
		RG_rl_13_t1 = TR_25 ;
	7'h16 :
		RG_rl_13_t1 = TR_25 ;
	7'h17 :
		RG_rl_13_t1 = TR_25 ;
	7'h18 :
		RG_rl_13_t1 = TR_25 ;
	7'h19 :
		RG_rl_13_t1 = TR_25 ;
	7'h1a :
		RG_rl_13_t1 = TR_25 ;
	7'h1b :
		RG_rl_13_t1 = TR_25 ;
	7'h1c :
		RG_rl_13_t1 = TR_25 ;
	7'h1d :
		RG_rl_13_t1 = TR_25 ;
	7'h1e :
		RG_rl_13_t1 = TR_25 ;
	7'h1f :
		RG_rl_13_t1 = TR_25 ;
	7'h20 :
		RG_rl_13_t1 = TR_25 ;
	7'h21 :
		RG_rl_13_t1 = TR_25 ;
	7'h22 :
		RG_rl_13_t1 = TR_25 ;
	7'h23 :
		RG_rl_13_t1 = TR_25 ;
	7'h24 :
		RG_rl_13_t1 = TR_25 ;
	7'h25 :
		RG_rl_13_t1 = TR_25 ;
	7'h26 :
		RG_rl_13_t1 = TR_25 ;
	7'h27 :
		RG_rl_13_t1 = TR_25 ;
	7'h28 :
		RG_rl_13_t1 = TR_25 ;
	7'h29 :
		RG_rl_13_t1 = TR_25 ;
	7'h2a :
		RG_rl_13_t1 = TR_25 ;
	7'h2b :
		RG_rl_13_t1 = TR_25 ;
	7'h2c :
		RG_rl_13_t1 = TR_25 ;
	7'h2d :
		RG_rl_13_t1 = TR_25 ;
	7'h2e :
		RG_rl_13_t1 = TR_25 ;
	7'h2f :
		RG_rl_13_t1 = TR_25 ;
	7'h30 :
		RG_rl_13_t1 = TR_25 ;
	7'h31 :
		RG_rl_13_t1 = TR_25 ;
	7'h32 :
		RG_rl_13_t1 = TR_25 ;
	7'h33 :
		RG_rl_13_t1 = TR_25 ;
	7'h34 :
		RG_rl_13_t1 = TR_25 ;
	7'h35 :
		RG_rl_13_t1 = TR_25 ;
	7'h36 :
		RG_rl_13_t1 = TR_25 ;
	7'h37 :
		RG_rl_13_t1 = TR_25 ;
	7'h38 :
		RG_rl_13_t1 = TR_25 ;
	7'h39 :
		RG_rl_13_t1 = TR_25 ;
	7'h3a :
		RG_rl_13_t1 = TR_25 ;
	7'h3b :
		RG_rl_13_t1 = TR_25 ;
	7'h3c :
		RG_rl_13_t1 = TR_25 ;
	7'h3d :
		RG_rl_13_t1 = TR_25 ;
	7'h3e :
		RG_rl_13_t1 = TR_25 ;
	7'h3f :
		RG_rl_13_t1 = TR_25 ;
	7'h40 :
		RG_rl_13_t1 = TR_25 ;
	7'h41 :
		RG_rl_13_t1 = TR_25 ;
	7'h42 :
		RG_rl_13_t1 = TR_25 ;
	7'h43 :
		RG_rl_13_t1 = TR_25 ;
	7'h44 :
		RG_rl_13_t1 = TR_25 ;
	7'h45 :
		RG_rl_13_t1 = TR_25 ;
	7'h46 :
		RG_rl_13_t1 = TR_25 ;
	7'h47 :
		RG_rl_13_t1 = TR_25 ;
	7'h48 :
		RG_rl_13_t1 = TR_25 ;
	7'h49 :
		RG_rl_13_t1 = TR_25 ;
	7'h4a :
		RG_rl_13_t1 = TR_25 ;
	7'h4b :
		RG_rl_13_t1 = TR_25 ;
	7'h4c :
		RG_rl_13_t1 = TR_25 ;
	7'h4d :
		RG_rl_13_t1 = TR_25 ;
	7'h4e :
		RG_rl_13_t1 = TR_25 ;
	7'h4f :
		RG_rl_13_t1 = TR_25 ;
	7'h50 :
		RG_rl_13_t1 = TR_25 ;
	7'h51 :
		RG_rl_13_t1 = TR_25 ;
	7'h52 :
		RG_rl_13_t1 = TR_25 ;
	7'h53 :
		RG_rl_13_t1 = TR_25 ;
	7'h54 :
		RG_rl_13_t1 = TR_25 ;
	7'h55 :
		RG_rl_13_t1 = TR_25 ;
	7'h56 :
		RG_rl_13_t1 = TR_25 ;
	7'h57 :
		RG_rl_13_t1 = TR_25 ;
	7'h58 :
		RG_rl_13_t1 = TR_25 ;
	7'h59 :
		RG_rl_13_t1 = TR_25 ;
	7'h5a :
		RG_rl_13_t1 = TR_25 ;
	7'h5b :
		RG_rl_13_t1 = TR_25 ;
	7'h5c :
		RG_rl_13_t1 = TR_25 ;
	7'h5d :
		RG_rl_13_t1 = TR_25 ;
	7'h5e :
		RG_rl_13_t1 = TR_25 ;
	7'h5f :
		RG_rl_13_t1 = TR_25 ;
	7'h60 :
		RG_rl_13_t1 = TR_25 ;
	7'h61 :
		RG_rl_13_t1 = TR_25 ;
	7'h62 :
		RG_rl_13_t1 = TR_25 ;
	7'h63 :
		RG_rl_13_t1 = TR_25 ;
	7'h64 :
		RG_rl_13_t1 = TR_25 ;
	7'h65 :
		RG_rl_13_t1 = TR_25 ;
	7'h66 :
		RG_rl_13_t1 = TR_25 ;
	7'h67 :
		RG_rl_13_t1 = TR_25 ;
	7'h68 :
		RG_rl_13_t1 = TR_25 ;
	7'h69 :
		RG_rl_13_t1 = TR_25 ;
	7'h6a :
		RG_rl_13_t1 = TR_25 ;
	7'h6b :
		RG_rl_13_t1 = TR_25 ;
	7'h6c :
		RG_rl_13_t1 = TR_25 ;
	7'h6d :
		RG_rl_13_t1 = TR_25 ;
	7'h6e :
		RG_rl_13_t1 = TR_25 ;
	7'h6f :
		RG_rl_13_t1 = TR_25 ;
	7'h70 :
		RG_rl_13_t1 = TR_25 ;
	7'h71 :
		RG_rl_13_t1 = TR_25 ;
	7'h72 :
		RG_rl_13_t1 = TR_25 ;
	7'h73 :
		RG_rl_13_t1 = TR_25 ;
	7'h74 :
		RG_rl_13_t1 = TR_25 ;
	7'h75 :
		RG_rl_13_t1 = TR_25 ;
	7'h76 :
		RG_rl_13_t1 = TR_25 ;
	7'h77 :
		RG_rl_13_t1 = TR_25 ;
	7'h78 :
		RG_rl_13_t1 = TR_25 ;
	7'h79 :
		RG_rl_13_t1 = TR_25 ;
	7'h7a :
		RG_rl_13_t1 = TR_25 ;
	7'h7b :
		RG_rl_13_t1 = TR_25 ;
	7'h7c :
		RG_rl_13_t1 = TR_25 ;
	7'h7d :
		RG_rl_13_t1 = TR_25 ;
	7'h7e :
		RG_rl_13_t1 = TR_25 ;
	7'h7f :
		RG_rl_13_t1 = TR_25 ;
	default :
		RG_rl_13_t1 = 9'hx ;
	endcase
always @ ( RG_rl_13_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_196 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_13_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h0d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_13_t = ( ( { 9{ U_570 } } & RG_rl_196 )
		| ( { 9{ U_569 } } & RG_rl_13_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_13_en = ( U_570 | RG_rl_13_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_13_en )
		RG_rl_13 <= RG_rl_13_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_26 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_14_t1 = TR_26 ;
	7'h01 :
		RG_rl_14_t1 = TR_26 ;
	7'h02 :
		RG_rl_14_t1 = TR_26 ;
	7'h03 :
		RG_rl_14_t1 = TR_26 ;
	7'h04 :
		RG_rl_14_t1 = TR_26 ;
	7'h05 :
		RG_rl_14_t1 = TR_26 ;
	7'h06 :
		RG_rl_14_t1 = TR_26 ;
	7'h07 :
		RG_rl_14_t1 = TR_26 ;
	7'h08 :
		RG_rl_14_t1 = TR_26 ;
	7'h09 :
		RG_rl_14_t1 = TR_26 ;
	7'h0a :
		RG_rl_14_t1 = TR_26 ;
	7'h0b :
		RG_rl_14_t1 = TR_26 ;
	7'h0c :
		RG_rl_14_t1 = TR_26 ;
	7'h0d :
		RG_rl_14_t1 = TR_26 ;
	7'h0e :
		RG_rl_14_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h0f :
		RG_rl_14_t1 = TR_26 ;
	7'h10 :
		RG_rl_14_t1 = TR_26 ;
	7'h11 :
		RG_rl_14_t1 = TR_26 ;
	7'h12 :
		RG_rl_14_t1 = TR_26 ;
	7'h13 :
		RG_rl_14_t1 = TR_26 ;
	7'h14 :
		RG_rl_14_t1 = TR_26 ;
	7'h15 :
		RG_rl_14_t1 = TR_26 ;
	7'h16 :
		RG_rl_14_t1 = TR_26 ;
	7'h17 :
		RG_rl_14_t1 = TR_26 ;
	7'h18 :
		RG_rl_14_t1 = TR_26 ;
	7'h19 :
		RG_rl_14_t1 = TR_26 ;
	7'h1a :
		RG_rl_14_t1 = TR_26 ;
	7'h1b :
		RG_rl_14_t1 = TR_26 ;
	7'h1c :
		RG_rl_14_t1 = TR_26 ;
	7'h1d :
		RG_rl_14_t1 = TR_26 ;
	7'h1e :
		RG_rl_14_t1 = TR_26 ;
	7'h1f :
		RG_rl_14_t1 = TR_26 ;
	7'h20 :
		RG_rl_14_t1 = TR_26 ;
	7'h21 :
		RG_rl_14_t1 = TR_26 ;
	7'h22 :
		RG_rl_14_t1 = TR_26 ;
	7'h23 :
		RG_rl_14_t1 = TR_26 ;
	7'h24 :
		RG_rl_14_t1 = TR_26 ;
	7'h25 :
		RG_rl_14_t1 = TR_26 ;
	7'h26 :
		RG_rl_14_t1 = TR_26 ;
	7'h27 :
		RG_rl_14_t1 = TR_26 ;
	7'h28 :
		RG_rl_14_t1 = TR_26 ;
	7'h29 :
		RG_rl_14_t1 = TR_26 ;
	7'h2a :
		RG_rl_14_t1 = TR_26 ;
	7'h2b :
		RG_rl_14_t1 = TR_26 ;
	7'h2c :
		RG_rl_14_t1 = TR_26 ;
	7'h2d :
		RG_rl_14_t1 = TR_26 ;
	7'h2e :
		RG_rl_14_t1 = TR_26 ;
	7'h2f :
		RG_rl_14_t1 = TR_26 ;
	7'h30 :
		RG_rl_14_t1 = TR_26 ;
	7'h31 :
		RG_rl_14_t1 = TR_26 ;
	7'h32 :
		RG_rl_14_t1 = TR_26 ;
	7'h33 :
		RG_rl_14_t1 = TR_26 ;
	7'h34 :
		RG_rl_14_t1 = TR_26 ;
	7'h35 :
		RG_rl_14_t1 = TR_26 ;
	7'h36 :
		RG_rl_14_t1 = TR_26 ;
	7'h37 :
		RG_rl_14_t1 = TR_26 ;
	7'h38 :
		RG_rl_14_t1 = TR_26 ;
	7'h39 :
		RG_rl_14_t1 = TR_26 ;
	7'h3a :
		RG_rl_14_t1 = TR_26 ;
	7'h3b :
		RG_rl_14_t1 = TR_26 ;
	7'h3c :
		RG_rl_14_t1 = TR_26 ;
	7'h3d :
		RG_rl_14_t1 = TR_26 ;
	7'h3e :
		RG_rl_14_t1 = TR_26 ;
	7'h3f :
		RG_rl_14_t1 = TR_26 ;
	7'h40 :
		RG_rl_14_t1 = TR_26 ;
	7'h41 :
		RG_rl_14_t1 = TR_26 ;
	7'h42 :
		RG_rl_14_t1 = TR_26 ;
	7'h43 :
		RG_rl_14_t1 = TR_26 ;
	7'h44 :
		RG_rl_14_t1 = TR_26 ;
	7'h45 :
		RG_rl_14_t1 = TR_26 ;
	7'h46 :
		RG_rl_14_t1 = TR_26 ;
	7'h47 :
		RG_rl_14_t1 = TR_26 ;
	7'h48 :
		RG_rl_14_t1 = TR_26 ;
	7'h49 :
		RG_rl_14_t1 = TR_26 ;
	7'h4a :
		RG_rl_14_t1 = TR_26 ;
	7'h4b :
		RG_rl_14_t1 = TR_26 ;
	7'h4c :
		RG_rl_14_t1 = TR_26 ;
	7'h4d :
		RG_rl_14_t1 = TR_26 ;
	7'h4e :
		RG_rl_14_t1 = TR_26 ;
	7'h4f :
		RG_rl_14_t1 = TR_26 ;
	7'h50 :
		RG_rl_14_t1 = TR_26 ;
	7'h51 :
		RG_rl_14_t1 = TR_26 ;
	7'h52 :
		RG_rl_14_t1 = TR_26 ;
	7'h53 :
		RG_rl_14_t1 = TR_26 ;
	7'h54 :
		RG_rl_14_t1 = TR_26 ;
	7'h55 :
		RG_rl_14_t1 = TR_26 ;
	7'h56 :
		RG_rl_14_t1 = TR_26 ;
	7'h57 :
		RG_rl_14_t1 = TR_26 ;
	7'h58 :
		RG_rl_14_t1 = TR_26 ;
	7'h59 :
		RG_rl_14_t1 = TR_26 ;
	7'h5a :
		RG_rl_14_t1 = TR_26 ;
	7'h5b :
		RG_rl_14_t1 = TR_26 ;
	7'h5c :
		RG_rl_14_t1 = TR_26 ;
	7'h5d :
		RG_rl_14_t1 = TR_26 ;
	7'h5e :
		RG_rl_14_t1 = TR_26 ;
	7'h5f :
		RG_rl_14_t1 = TR_26 ;
	7'h60 :
		RG_rl_14_t1 = TR_26 ;
	7'h61 :
		RG_rl_14_t1 = TR_26 ;
	7'h62 :
		RG_rl_14_t1 = TR_26 ;
	7'h63 :
		RG_rl_14_t1 = TR_26 ;
	7'h64 :
		RG_rl_14_t1 = TR_26 ;
	7'h65 :
		RG_rl_14_t1 = TR_26 ;
	7'h66 :
		RG_rl_14_t1 = TR_26 ;
	7'h67 :
		RG_rl_14_t1 = TR_26 ;
	7'h68 :
		RG_rl_14_t1 = TR_26 ;
	7'h69 :
		RG_rl_14_t1 = TR_26 ;
	7'h6a :
		RG_rl_14_t1 = TR_26 ;
	7'h6b :
		RG_rl_14_t1 = TR_26 ;
	7'h6c :
		RG_rl_14_t1 = TR_26 ;
	7'h6d :
		RG_rl_14_t1 = TR_26 ;
	7'h6e :
		RG_rl_14_t1 = TR_26 ;
	7'h6f :
		RG_rl_14_t1 = TR_26 ;
	7'h70 :
		RG_rl_14_t1 = TR_26 ;
	7'h71 :
		RG_rl_14_t1 = TR_26 ;
	7'h72 :
		RG_rl_14_t1 = TR_26 ;
	7'h73 :
		RG_rl_14_t1 = TR_26 ;
	7'h74 :
		RG_rl_14_t1 = TR_26 ;
	7'h75 :
		RG_rl_14_t1 = TR_26 ;
	7'h76 :
		RG_rl_14_t1 = TR_26 ;
	7'h77 :
		RG_rl_14_t1 = TR_26 ;
	7'h78 :
		RG_rl_14_t1 = TR_26 ;
	7'h79 :
		RG_rl_14_t1 = TR_26 ;
	7'h7a :
		RG_rl_14_t1 = TR_26 ;
	7'h7b :
		RG_rl_14_t1 = TR_26 ;
	7'h7c :
		RG_rl_14_t1 = TR_26 ;
	7'h7d :
		RG_rl_14_t1 = TR_26 ;
	7'h7e :
		RG_rl_14_t1 = TR_26 ;
	7'h7f :
		RG_rl_14_t1 = TR_26 ;
	default :
		RG_rl_14_t1 = 9'hx ;
	endcase
always @ ( RG_rl_14_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_197 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_14_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h0e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_14_t = ( ( { 9{ U_570 } } & RG_rl_197 )
		| ( { 9{ U_569 } } & RG_rl_14_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_14_en = ( U_570 | RG_rl_14_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_14_en )
		RG_rl_14 <= RG_rl_14_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_27 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_15_t1 = TR_27 ;
	7'h01 :
		RG_rl_15_t1 = TR_27 ;
	7'h02 :
		RG_rl_15_t1 = TR_27 ;
	7'h03 :
		RG_rl_15_t1 = TR_27 ;
	7'h04 :
		RG_rl_15_t1 = TR_27 ;
	7'h05 :
		RG_rl_15_t1 = TR_27 ;
	7'h06 :
		RG_rl_15_t1 = TR_27 ;
	7'h07 :
		RG_rl_15_t1 = TR_27 ;
	7'h08 :
		RG_rl_15_t1 = TR_27 ;
	7'h09 :
		RG_rl_15_t1 = TR_27 ;
	7'h0a :
		RG_rl_15_t1 = TR_27 ;
	7'h0b :
		RG_rl_15_t1 = TR_27 ;
	7'h0c :
		RG_rl_15_t1 = TR_27 ;
	7'h0d :
		RG_rl_15_t1 = TR_27 ;
	7'h0e :
		RG_rl_15_t1 = TR_27 ;
	7'h0f :
		RG_rl_15_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h10 :
		RG_rl_15_t1 = TR_27 ;
	7'h11 :
		RG_rl_15_t1 = TR_27 ;
	7'h12 :
		RG_rl_15_t1 = TR_27 ;
	7'h13 :
		RG_rl_15_t1 = TR_27 ;
	7'h14 :
		RG_rl_15_t1 = TR_27 ;
	7'h15 :
		RG_rl_15_t1 = TR_27 ;
	7'h16 :
		RG_rl_15_t1 = TR_27 ;
	7'h17 :
		RG_rl_15_t1 = TR_27 ;
	7'h18 :
		RG_rl_15_t1 = TR_27 ;
	7'h19 :
		RG_rl_15_t1 = TR_27 ;
	7'h1a :
		RG_rl_15_t1 = TR_27 ;
	7'h1b :
		RG_rl_15_t1 = TR_27 ;
	7'h1c :
		RG_rl_15_t1 = TR_27 ;
	7'h1d :
		RG_rl_15_t1 = TR_27 ;
	7'h1e :
		RG_rl_15_t1 = TR_27 ;
	7'h1f :
		RG_rl_15_t1 = TR_27 ;
	7'h20 :
		RG_rl_15_t1 = TR_27 ;
	7'h21 :
		RG_rl_15_t1 = TR_27 ;
	7'h22 :
		RG_rl_15_t1 = TR_27 ;
	7'h23 :
		RG_rl_15_t1 = TR_27 ;
	7'h24 :
		RG_rl_15_t1 = TR_27 ;
	7'h25 :
		RG_rl_15_t1 = TR_27 ;
	7'h26 :
		RG_rl_15_t1 = TR_27 ;
	7'h27 :
		RG_rl_15_t1 = TR_27 ;
	7'h28 :
		RG_rl_15_t1 = TR_27 ;
	7'h29 :
		RG_rl_15_t1 = TR_27 ;
	7'h2a :
		RG_rl_15_t1 = TR_27 ;
	7'h2b :
		RG_rl_15_t1 = TR_27 ;
	7'h2c :
		RG_rl_15_t1 = TR_27 ;
	7'h2d :
		RG_rl_15_t1 = TR_27 ;
	7'h2e :
		RG_rl_15_t1 = TR_27 ;
	7'h2f :
		RG_rl_15_t1 = TR_27 ;
	7'h30 :
		RG_rl_15_t1 = TR_27 ;
	7'h31 :
		RG_rl_15_t1 = TR_27 ;
	7'h32 :
		RG_rl_15_t1 = TR_27 ;
	7'h33 :
		RG_rl_15_t1 = TR_27 ;
	7'h34 :
		RG_rl_15_t1 = TR_27 ;
	7'h35 :
		RG_rl_15_t1 = TR_27 ;
	7'h36 :
		RG_rl_15_t1 = TR_27 ;
	7'h37 :
		RG_rl_15_t1 = TR_27 ;
	7'h38 :
		RG_rl_15_t1 = TR_27 ;
	7'h39 :
		RG_rl_15_t1 = TR_27 ;
	7'h3a :
		RG_rl_15_t1 = TR_27 ;
	7'h3b :
		RG_rl_15_t1 = TR_27 ;
	7'h3c :
		RG_rl_15_t1 = TR_27 ;
	7'h3d :
		RG_rl_15_t1 = TR_27 ;
	7'h3e :
		RG_rl_15_t1 = TR_27 ;
	7'h3f :
		RG_rl_15_t1 = TR_27 ;
	7'h40 :
		RG_rl_15_t1 = TR_27 ;
	7'h41 :
		RG_rl_15_t1 = TR_27 ;
	7'h42 :
		RG_rl_15_t1 = TR_27 ;
	7'h43 :
		RG_rl_15_t1 = TR_27 ;
	7'h44 :
		RG_rl_15_t1 = TR_27 ;
	7'h45 :
		RG_rl_15_t1 = TR_27 ;
	7'h46 :
		RG_rl_15_t1 = TR_27 ;
	7'h47 :
		RG_rl_15_t1 = TR_27 ;
	7'h48 :
		RG_rl_15_t1 = TR_27 ;
	7'h49 :
		RG_rl_15_t1 = TR_27 ;
	7'h4a :
		RG_rl_15_t1 = TR_27 ;
	7'h4b :
		RG_rl_15_t1 = TR_27 ;
	7'h4c :
		RG_rl_15_t1 = TR_27 ;
	7'h4d :
		RG_rl_15_t1 = TR_27 ;
	7'h4e :
		RG_rl_15_t1 = TR_27 ;
	7'h4f :
		RG_rl_15_t1 = TR_27 ;
	7'h50 :
		RG_rl_15_t1 = TR_27 ;
	7'h51 :
		RG_rl_15_t1 = TR_27 ;
	7'h52 :
		RG_rl_15_t1 = TR_27 ;
	7'h53 :
		RG_rl_15_t1 = TR_27 ;
	7'h54 :
		RG_rl_15_t1 = TR_27 ;
	7'h55 :
		RG_rl_15_t1 = TR_27 ;
	7'h56 :
		RG_rl_15_t1 = TR_27 ;
	7'h57 :
		RG_rl_15_t1 = TR_27 ;
	7'h58 :
		RG_rl_15_t1 = TR_27 ;
	7'h59 :
		RG_rl_15_t1 = TR_27 ;
	7'h5a :
		RG_rl_15_t1 = TR_27 ;
	7'h5b :
		RG_rl_15_t1 = TR_27 ;
	7'h5c :
		RG_rl_15_t1 = TR_27 ;
	7'h5d :
		RG_rl_15_t1 = TR_27 ;
	7'h5e :
		RG_rl_15_t1 = TR_27 ;
	7'h5f :
		RG_rl_15_t1 = TR_27 ;
	7'h60 :
		RG_rl_15_t1 = TR_27 ;
	7'h61 :
		RG_rl_15_t1 = TR_27 ;
	7'h62 :
		RG_rl_15_t1 = TR_27 ;
	7'h63 :
		RG_rl_15_t1 = TR_27 ;
	7'h64 :
		RG_rl_15_t1 = TR_27 ;
	7'h65 :
		RG_rl_15_t1 = TR_27 ;
	7'h66 :
		RG_rl_15_t1 = TR_27 ;
	7'h67 :
		RG_rl_15_t1 = TR_27 ;
	7'h68 :
		RG_rl_15_t1 = TR_27 ;
	7'h69 :
		RG_rl_15_t1 = TR_27 ;
	7'h6a :
		RG_rl_15_t1 = TR_27 ;
	7'h6b :
		RG_rl_15_t1 = TR_27 ;
	7'h6c :
		RG_rl_15_t1 = TR_27 ;
	7'h6d :
		RG_rl_15_t1 = TR_27 ;
	7'h6e :
		RG_rl_15_t1 = TR_27 ;
	7'h6f :
		RG_rl_15_t1 = TR_27 ;
	7'h70 :
		RG_rl_15_t1 = TR_27 ;
	7'h71 :
		RG_rl_15_t1 = TR_27 ;
	7'h72 :
		RG_rl_15_t1 = TR_27 ;
	7'h73 :
		RG_rl_15_t1 = TR_27 ;
	7'h74 :
		RG_rl_15_t1 = TR_27 ;
	7'h75 :
		RG_rl_15_t1 = TR_27 ;
	7'h76 :
		RG_rl_15_t1 = TR_27 ;
	7'h77 :
		RG_rl_15_t1 = TR_27 ;
	7'h78 :
		RG_rl_15_t1 = TR_27 ;
	7'h79 :
		RG_rl_15_t1 = TR_27 ;
	7'h7a :
		RG_rl_15_t1 = TR_27 ;
	7'h7b :
		RG_rl_15_t1 = TR_27 ;
	7'h7c :
		RG_rl_15_t1 = TR_27 ;
	7'h7d :
		RG_rl_15_t1 = TR_27 ;
	7'h7e :
		RG_rl_15_t1 = TR_27 ;
	7'h7f :
		RG_rl_15_t1 = TR_27 ;
	default :
		RG_rl_15_t1 = 9'hx ;
	endcase
always @ ( RG_rl_15_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_198 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_15_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h0f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_15_t = ( ( { 9{ U_570 } } & RG_rl_198 )
		| ( { 9{ U_569 } } & RG_rl_15_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_15_en = ( U_570 | RG_rl_15_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_15_en )
		RG_rl_15 <= RG_rl_15_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_28 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_16_t1 = TR_28 ;
	7'h01 :
		RG_rl_16_t1 = TR_28 ;
	7'h02 :
		RG_rl_16_t1 = TR_28 ;
	7'h03 :
		RG_rl_16_t1 = TR_28 ;
	7'h04 :
		RG_rl_16_t1 = TR_28 ;
	7'h05 :
		RG_rl_16_t1 = TR_28 ;
	7'h06 :
		RG_rl_16_t1 = TR_28 ;
	7'h07 :
		RG_rl_16_t1 = TR_28 ;
	7'h08 :
		RG_rl_16_t1 = TR_28 ;
	7'h09 :
		RG_rl_16_t1 = TR_28 ;
	7'h0a :
		RG_rl_16_t1 = TR_28 ;
	7'h0b :
		RG_rl_16_t1 = TR_28 ;
	7'h0c :
		RG_rl_16_t1 = TR_28 ;
	7'h0d :
		RG_rl_16_t1 = TR_28 ;
	7'h0e :
		RG_rl_16_t1 = TR_28 ;
	7'h0f :
		RG_rl_16_t1 = TR_28 ;
	7'h10 :
		RG_rl_16_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h11 :
		RG_rl_16_t1 = TR_28 ;
	7'h12 :
		RG_rl_16_t1 = TR_28 ;
	7'h13 :
		RG_rl_16_t1 = TR_28 ;
	7'h14 :
		RG_rl_16_t1 = TR_28 ;
	7'h15 :
		RG_rl_16_t1 = TR_28 ;
	7'h16 :
		RG_rl_16_t1 = TR_28 ;
	7'h17 :
		RG_rl_16_t1 = TR_28 ;
	7'h18 :
		RG_rl_16_t1 = TR_28 ;
	7'h19 :
		RG_rl_16_t1 = TR_28 ;
	7'h1a :
		RG_rl_16_t1 = TR_28 ;
	7'h1b :
		RG_rl_16_t1 = TR_28 ;
	7'h1c :
		RG_rl_16_t1 = TR_28 ;
	7'h1d :
		RG_rl_16_t1 = TR_28 ;
	7'h1e :
		RG_rl_16_t1 = TR_28 ;
	7'h1f :
		RG_rl_16_t1 = TR_28 ;
	7'h20 :
		RG_rl_16_t1 = TR_28 ;
	7'h21 :
		RG_rl_16_t1 = TR_28 ;
	7'h22 :
		RG_rl_16_t1 = TR_28 ;
	7'h23 :
		RG_rl_16_t1 = TR_28 ;
	7'h24 :
		RG_rl_16_t1 = TR_28 ;
	7'h25 :
		RG_rl_16_t1 = TR_28 ;
	7'h26 :
		RG_rl_16_t1 = TR_28 ;
	7'h27 :
		RG_rl_16_t1 = TR_28 ;
	7'h28 :
		RG_rl_16_t1 = TR_28 ;
	7'h29 :
		RG_rl_16_t1 = TR_28 ;
	7'h2a :
		RG_rl_16_t1 = TR_28 ;
	7'h2b :
		RG_rl_16_t1 = TR_28 ;
	7'h2c :
		RG_rl_16_t1 = TR_28 ;
	7'h2d :
		RG_rl_16_t1 = TR_28 ;
	7'h2e :
		RG_rl_16_t1 = TR_28 ;
	7'h2f :
		RG_rl_16_t1 = TR_28 ;
	7'h30 :
		RG_rl_16_t1 = TR_28 ;
	7'h31 :
		RG_rl_16_t1 = TR_28 ;
	7'h32 :
		RG_rl_16_t1 = TR_28 ;
	7'h33 :
		RG_rl_16_t1 = TR_28 ;
	7'h34 :
		RG_rl_16_t1 = TR_28 ;
	7'h35 :
		RG_rl_16_t1 = TR_28 ;
	7'h36 :
		RG_rl_16_t1 = TR_28 ;
	7'h37 :
		RG_rl_16_t1 = TR_28 ;
	7'h38 :
		RG_rl_16_t1 = TR_28 ;
	7'h39 :
		RG_rl_16_t1 = TR_28 ;
	7'h3a :
		RG_rl_16_t1 = TR_28 ;
	7'h3b :
		RG_rl_16_t1 = TR_28 ;
	7'h3c :
		RG_rl_16_t1 = TR_28 ;
	7'h3d :
		RG_rl_16_t1 = TR_28 ;
	7'h3e :
		RG_rl_16_t1 = TR_28 ;
	7'h3f :
		RG_rl_16_t1 = TR_28 ;
	7'h40 :
		RG_rl_16_t1 = TR_28 ;
	7'h41 :
		RG_rl_16_t1 = TR_28 ;
	7'h42 :
		RG_rl_16_t1 = TR_28 ;
	7'h43 :
		RG_rl_16_t1 = TR_28 ;
	7'h44 :
		RG_rl_16_t1 = TR_28 ;
	7'h45 :
		RG_rl_16_t1 = TR_28 ;
	7'h46 :
		RG_rl_16_t1 = TR_28 ;
	7'h47 :
		RG_rl_16_t1 = TR_28 ;
	7'h48 :
		RG_rl_16_t1 = TR_28 ;
	7'h49 :
		RG_rl_16_t1 = TR_28 ;
	7'h4a :
		RG_rl_16_t1 = TR_28 ;
	7'h4b :
		RG_rl_16_t1 = TR_28 ;
	7'h4c :
		RG_rl_16_t1 = TR_28 ;
	7'h4d :
		RG_rl_16_t1 = TR_28 ;
	7'h4e :
		RG_rl_16_t1 = TR_28 ;
	7'h4f :
		RG_rl_16_t1 = TR_28 ;
	7'h50 :
		RG_rl_16_t1 = TR_28 ;
	7'h51 :
		RG_rl_16_t1 = TR_28 ;
	7'h52 :
		RG_rl_16_t1 = TR_28 ;
	7'h53 :
		RG_rl_16_t1 = TR_28 ;
	7'h54 :
		RG_rl_16_t1 = TR_28 ;
	7'h55 :
		RG_rl_16_t1 = TR_28 ;
	7'h56 :
		RG_rl_16_t1 = TR_28 ;
	7'h57 :
		RG_rl_16_t1 = TR_28 ;
	7'h58 :
		RG_rl_16_t1 = TR_28 ;
	7'h59 :
		RG_rl_16_t1 = TR_28 ;
	7'h5a :
		RG_rl_16_t1 = TR_28 ;
	7'h5b :
		RG_rl_16_t1 = TR_28 ;
	7'h5c :
		RG_rl_16_t1 = TR_28 ;
	7'h5d :
		RG_rl_16_t1 = TR_28 ;
	7'h5e :
		RG_rl_16_t1 = TR_28 ;
	7'h5f :
		RG_rl_16_t1 = TR_28 ;
	7'h60 :
		RG_rl_16_t1 = TR_28 ;
	7'h61 :
		RG_rl_16_t1 = TR_28 ;
	7'h62 :
		RG_rl_16_t1 = TR_28 ;
	7'h63 :
		RG_rl_16_t1 = TR_28 ;
	7'h64 :
		RG_rl_16_t1 = TR_28 ;
	7'h65 :
		RG_rl_16_t1 = TR_28 ;
	7'h66 :
		RG_rl_16_t1 = TR_28 ;
	7'h67 :
		RG_rl_16_t1 = TR_28 ;
	7'h68 :
		RG_rl_16_t1 = TR_28 ;
	7'h69 :
		RG_rl_16_t1 = TR_28 ;
	7'h6a :
		RG_rl_16_t1 = TR_28 ;
	7'h6b :
		RG_rl_16_t1 = TR_28 ;
	7'h6c :
		RG_rl_16_t1 = TR_28 ;
	7'h6d :
		RG_rl_16_t1 = TR_28 ;
	7'h6e :
		RG_rl_16_t1 = TR_28 ;
	7'h6f :
		RG_rl_16_t1 = TR_28 ;
	7'h70 :
		RG_rl_16_t1 = TR_28 ;
	7'h71 :
		RG_rl_16_t1 = TR_28 ;
	7'h72 :
		RG_rl_16_t1 = TR_28 ;
	7'h73 :
		RG_rl_16_t1 = TR_28 ;
	7'h74 :
		RG_rl_16_t1 = TR_28 ;
	7'h75 :
		RG_rl_16_t1 = TR_28 ;
	7'h76 :
		RG_rl_16_t1 = TR_28 ;
	7'h77 :
		RG_rl_16_t1 = TR_28 ;
	7'h78 :
		RG_rl_16_t1 = TR_28 ;
	7'h79 :
		RG_rl_16_t1 = TR_28 ;
	7'h7a :
		RG_rl_16_t1 = TR_28 ;
	7'h7b :
		RG_rl_16_t1 = TR_28 ;
	7'h7c :
		RG_rl_16_t1 = TR_28 ;
	7'h7d :
		RG_rl_16_t1 = TR_28 ;
	7'h7e :
		RG_rl_16_t1 = TR_28 ;
	7'h7f :
		RG_rl_16_t1 = TR_28 ;
	default :
		RG_rl_16_t1 = 9'hx ;
	endcase
always @ ( RG_rl_16_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_199 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_16_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h10 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_16_t = ( ( { 9{ U_570 } } & RG_rl_199 )
		| ( { 9{ U_569 } } & RG_rl_16_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_16_en = ( U_570 | RG_rl_16_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_16_en )
		RG_rl_16 <= RG_rl_16_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_29 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_17_t1 = TR_29 ;
	7'h01 :
		RG_rl_17_t1 = TR_29 ;
	7'h02 :
		RG_rl_17_t1 = TR_29 ;
	7'h03 :
		RG_rl_17_t1 = TR_29 ;
	7'h04 :
		RG_rl_17_t1 = TR_29 ;
	7'h05 :
		RG_rl_17_t1 = TR_29 ;
	7'h06 :
		RG_rl_17_t1 = TR_29 ;
	7'h07 :
		RG_rl_17_t1 = TR_29 ;
	7'h08 :
		RG_rl_17_t1 = TR_29 ;
	7'h09 :
		RG_rl_17_t1 = TR_29 ;
	7'h0a :
		RG_rl_17_t1 = TR_29 ;
	7'h0b :
		RG_rl_17_t1 = TR_29 ;
	7'h0c :
		RG_rl_17_t1 = TR_29 ;
	7'h0d :
		RG_rl_17_t1 = TR_29 ;
	7'h0e :
		RG_rl_17_t1 = TR_29 ;
	7'h0f :
		RG_rl_17_t1 = TR_29 ;
	7'h10 :
		RG_rl_17_t1 = TR_29 ;
	7'h11 :
		RG_rl_17_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h12 :
		RG_rl_17_t1 = TR_29 ;
	7'h13 :
		RG_rl_17_t1 = TR_29 ;
	7'h14 :
		RG_rl_17_t1 = TR_29 ;
	7'h15 :
		RG_rl_17_t1 = TR_29 ;
	7'h16 :
		RG_rl_17_t1 = TR_29 ;
	7'h17 :
		RG_rl_17_t1 = TR_29 ;
	7'h18 :
		RG_rl_17_t1 = TR_29 ;
	7'h19 :
		RG_rl_17_t1 = TR_29 ;
	7'h1a :
		RG_rl_17_t1 = TR_29 ;
	7'h1b :
		RG_rl_17_t1 = TR_29 ;
	7'h1c :
		RG_rl_17_t1 = TR_29 ;
	7'h1d :
		RG_rl_17_t1 = TR_29 ;
	7'h1e :
		RG_rl_17_t1 = TR_29 ;
	7'h1f :
		RG_rl_17_t1 = TR_29 ;
	7'h20 :
		RG_rl_17_t1 = TR_29 ;
	7'h21 :
		RG_rl_17_t1 = TR_29 ;
	7'h22 :
		RG_rl_17_t1 = TR_29 ;
	7'h23 :
		RG_rl_17_t1 = TR_29 ;
	7'h24 :
		RG_rl_17_t1 = TR_29 ;
	7'h25 :
		RG_rl_17_t1 = TR_29 ;
	7'h26 :
		RG_rl_17_t1 = TR_29 ;
	7'h27 :
		RG_rl_17_t1 = TR_29 ;
	7'h28 :
		RG_rl_17_t1 = TR_29 ;
	7'h29 :
		RG_rl_17_t1 = TR_29 ;
	7'h2a :
		RG_rl_17_t1 = TR_29 ;
	7'h2b :
		RG_rl_17_t1 = TR_29 ;
	7'h2c :
		RG_rl_17_t1 = TR_29 ;
	7'h2d :
		RG_rl_17_t1 = TR_29 ;
	7'h2e :
		RG_rl_17_t1 = TR_29 ;
	7'h2f :
		RG_rl_17_t1 = TR_29 ;
	7'h30 :
		RG_rl_17_t1 = TR_29 ;
	7'h31 :
		RG_rl_17_t1 = TR_29 ;
	7'h32 :
		RG_rl_17_t1 = TR_29 ;
	7'h33 :
		RG_rl_17_t1 = TR_29 ;
	7'h34 :
		RG_rl_17_t1 = TR_29 ;
	7'h35 :
		RG_rl_17_t1 = TR_29 ;
	7'h36 :
		RG_rl_17_t1 = TR_29 ;
	7'h37 :
		RG_rl_17_t1 = TR_29 ;
	7'h38 :
		RG_rl_17_t1 = TR_29 ;
	7'h39 :
		RG_rl_17_t1 = TR_29 ;
	7'h3a :
		RG_rl_17_t1 = TR_29 ;
	7'h3b :
		RG_rl_17_t1 = TR_29 ;
	7'h3c :
		RG_rl_17_t1 = TR_29 ;
	7'h3d :
		RG_rl_17_t1 = TR_29 ;
	7'h3e :
		RG_rl_17_t1 = TR_29 ;
	7'h3f :
		RG_rl_17_t1 = TR_29 ;
	7'h40 :
		RG_rl_17_t1 = TR_29 ;
	7'h41 :
		RG_rl_17_t1 = TR_29 ;
	7'h42 :
		RG_rl_17_t1 = TR_29 ;
	7'h43 :
		RG_rl_17_t1 = TR_29 ;
	7'h44 :
		RG_rl_17_t1 = TR_29 ;
	7'h45 :
		RG_rl_17_t1 = TR_29 ;
	7'h46 :
		RG_rl_17_t1 = TR_29 ;
	7'h47 :
		RG_rl_17_t1 = TR_29 ;
	7'h48 :
		RG_rl_17_t1 = TR_29 ;
	7'h49 :
		RG_rl_17_t1 = TR_29 ;
	7'h4a :
		RG_rl_17_t1 = TR_29 ;
	7'h4b :
		RG_rl_17_t1 = TR_29 ;
	7'h4c :
		RG_rl_17_t1 = TR_29 ;
	7'h4d :
		RG_rl_17_t1 = TR_29 ;
	7'h4e :
		RG_rl_17_t1 = TR_29 ;
	7'h4f :
		RG_rl_17_t1 = TR_29 ;
	7'h50 :
		RG_rl_17_t1 = TR_29 ;
	7'h51 :
		RG_rl_17_t1 = TR_29 ;
	7'h52 :
		RG_rl_17_t1 = TR_29 ;
	7'h53 :
		RG_rl_17_t1 = TR_29 ;
	7'h54 :
		RG_rl_17_t1 = TR_29 ;
	7'h55 :
		RG_rl_17_t1 = TR_29 ;
	7'h56 :
		RG_rl_17_t1 = TR_29 ;
	7'h57 :
		RG_rl_17_t1 = TR_29 ;
	7'h58 :
		RG_rl_17_t1 = TR_29 ;
	7'h59 :
		RG_rl_17_t1 = TR_29 ;
	7'h5a :
		RG_rl_17_t1 = TR_29 ;
	7'h5b :
		RG_rl_17_t1 = TR_29 ;
	7'h5c :
		RG_rl_17_t1 = TR_29 ;
	7'h5d :
		RG_rl_17_t1 = TR_29 ;
	7'h5e :
		RG_rl_17_t1 = TR_29 ;
	7'h5f :
		RG_rl_17_t1 = TR_29 ;
	7'h60 :
		RG_rl_17_t1 = TR_29 ;
	7'h61 :
		RG_rl_17_t1 = TR_29 ;
	7'h62 :
		RG_rl_17_t1 = TR_29 ;
	7'h63 :
		RG_rl_17_t1 = TR_29 ;
	7'h64 :
		RG_rl_17_t1 = TR_29 ;
	7'h65 :
		RG_rl_17_t1 = TR_29 ;
	7'h66 :
		RG_rl_17_t1 = TR_29 ;
	7'h67 :
		RG_rl_17_t1 = TR_29 ;
	7'h68 :
		RG_rl_17_t1 = TR_29 ;
	7'h69 :
		RG_rl_17_t1 = TR_29 ;
	7'h6a :
		RG_rl_17_t1 = TR_29 ;
	7'h6b :
		RG_rl_17_t1 = TR_29 ;
	7'h6c :
		RG_rl_17_t1 = TR_29 ;
	7'h6d :
		RG_rl_17_t1 = TR_29 ;
	7'h6e :
		RG_rl_17_t1 = TR_29 ;
	7'h6f :
		RG_rl_17_t1 = TR_29 ;
	7'h70 :
		RG_rl_17_t1 = TR_29 ;
	7'h71 :
		RG_rl_17_t1 = TR_29 ;
	7'h72 :
		RG_rl_17_t1 = TR_29 ;
	7'h73 :
		RG_rl_17_t1 = TR_29 ;
	7'h74 :
		RG_rl_17_t1 = TR_29 ;
	7'h75 :
		RG_rl_17_t1 = TR_29 ;
	7'h76 :
		RG_rl_17_t1 = TR_29 ;
	7'h77 :
		RG_rl_17_t1 = TR_29 ;
	7'h78 :
		RG_rl_17_t1 = TR_29 ;
	7'h79 :
		RG_rl_17_t1 = TR_29 ;
	7'h7a :
		RG_rl_17_t1 = TR_29 ;
	7'h7b :
		RG_rl_17_t1 = TR_29 ;
	7'h7c :
		RG_rl_17_t1 = TR_29 ;
	7'h7d :
		RG_rl_17_t1 = TR_29 ;
	7'h7e :
		RG_rl_17_t1 = TR_29 ;
	7'h7f :
		RG_rl_17_t1 = TR_29 ;
	default :
		RG_rl_17_t1 = 9'hx ;
	endcase
always @ ( RG_rl_17_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_200 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_17_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h11 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_17_t = ( ( { 9{ U_570 } } & RG_rl_200 )
		| ( { 9{ U_569 } } & RG_rl_17_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_17_en = ( U_570 | RG_rl_17_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_17_en )
		RG_rl_17 <= RG_rl_17_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_30 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_18_t1 = TR_30 ;
	7'h01 :
		RG_rl_18_t1 = TR_30 ;
	7'h02 :
		RG_rl_18_t1 = TR_30 ;
	7'h03 :
		RG_rl_18_t1 = TR_30 ;
	7'h04 :
		RG_rl_18_t1 = TR_30 ;
	7'h05 :
		RG_rl_18_t1 = TR_30 ;
	7'h06 :
		RG_rl_18_t1 = TR_30 ;
	7'h07 :
		RG_rl_18_t1 = TR_30 ;
	7'h08 :
		RG_rl_18_t1 = TR_30 ;
	7'h09 :
		RG_rl_18_t1 = TR_30 ;
	7'h0a :
		RG_rl_18_t1 = TR_30 ;
	7'h0b :
		RG_rl_18_t1 = TR_30 ;
	7'h0c :
		RG_rl_18_t1 = TR_30 ;
	7'h0d :
		RG_rl_18_t1 = TR_30 ;
	7'h0e :
		RG_rl_18_t1 = TR_30 ;
	7'h0f :
		RG_rl_18_t1 = TR_30 ;
	7'h10 :
		RG_rl_18_t1 = TR_30 ;
	7'h11 :
		RG_rl_18_t1 = TR_30 ;
	7'h12 :
		RG_rl_18_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h13 :
		RG_rl_18_t1 = TR_30 ;
	7'h14 :
		RG_rl_18_t1 = TR_30 ;
	7'h15 :
		RG_rl_18_t1 = TR_30 ;
	7'h16 :
		RG_rl_18_t1 = TR_30 ;
	7'h17 :
		RG_rl_18_t1 = TR_30 ;
	7'h18 :
		RG_rl_18_t1 = TR_30 ;
	7'h19 :
		RG_rl_18_t1 = TR_30 ;
	7'h1a :
		RG_rl_18_t1 = TR_30 ;
	7'h1b :
		RG_rl_18_t1 = TR_30 ;
	7'h1c :
		RG_rl_18_t1 = TR_30 ;
	7'h1d :
		RG_rl_18_t1 = TR_30 ;
	7'h1e :
		RG_rl_18_t1 = TR_30 ;
	7'h1f :
		RG_rl_18_t1 = TR_30 ;
	7'h20 :
		RG_rl_18_t1 = TR_30 ;
	7'h21 :
		RG_rl_18_t1 = TR_30 ;
	7'h22 :
		RG_rl_18_t1 = TR_30 ;
	7'h23 :
		RG_rl_18_t1 = TR_30 ;
	7'h24 :
		RG_rl_18_t1 = TR_30 ;
	7'h25 :
		RG_rl_18_t1 = TR_30 ;
	7'h26 :
		RG_rl_18_t1 = TR_30 ;
	7'h27 :
		RG_rl_18_t1 = TR_30 ;
	7'h28 :
		RG_rl_18_t1 = TR_30 ;
	7'h29 :
		RG_rl_18_t1 = TR_30 ;
	7'h2a :
		RG_rl_18_t1 = TR_30 ;
	7'h2b :
		RG_rl_18_t1 = TR_30 ;
	7'h2c :
		RG_rl_18_t1 = TR_30 ;
	7'h2d :
		RG_rl_18_t1 = TR_30 ;
	7'h2e :
		RG_rl_18_t1 = TR_30 ;
	7'h2f :
		RG_rl_18_t1 = TR_30 ;
	7'h30 :
		RG_rl_18_t1 = TR_30 ;
	7'h31 :
		RG_rl_18_t1 = TR_30 ;
	7'h32 :
		RG_rl_18_t1 = TR_30 ;
	7'h33 :
		RG_rl_18_t1 = TR_30 ;
	7'h34 :
		RG_rl_18_t1 = TR_30 ;
	7'h35 :
		RG_rl_18_t1 = TR_30 ;
	7'h36 :
		RG_rl_18_t1 = TR_30 ;
	7'h37 :
		RG_rl_18_t1 = TR_30 ;
	7'h38 :
		RG_rl_18_t1 = TR_30 ;
	7'h39 :
		RG_rl_18_t1 = TR_30 ;
	7'h3a :
		RG_rl_18_t1 = TR_30 ;
	7'h3b :
		RG_rl_18_t1 = TR_30 ;
	7'h3c :
		RG_rl_18_t1 = TR_30 ;
	7'h3d :
		RG_rl_18_t1 = TR_30 ;
	7'h3e :
		RG_rl_18_t1 = TR_30 ;
	7'h3f :
		RG_rl_18_t1 = TR_30 ;
	7'h40 :
		RG_rl_18_t1 = TR_30 ;
	7'h41 :
		RG_rl_18_t1 = TR_30 ;
	7'h42 :
		RG_rl_18_t1 = TR_30 ;
	7'h43 :
		RG_rl_18_t1 = TR_30 ;
	7'h44 :
		RG_rl_18_t1 = TR_30 ;
	7'h45 :
		RG_rl_18_t1 = TR_30 ;
	7'h46 :
		RG_rl_18_t1 = TR_30 ;
	7'h47 :
		RG_rl_18_t1 = TR_30 ;
	7'h48 :
		RG_rl_18_t1 = TR_30 ;
	7'h49 :
		RG_rl_18_t1 = TR_30 ;
	7'h4a :
		RG_rl_18_t1 = TR_30 ;
	7'h4b :
		RG_rl_18_t1 = TR_30 ;
	7'h4c :
		RG_rl_18_t1 = TR_30 ;
	7'h4d :
		RG_rl_18_t1 = TR_30 ;
	7'h4e :
		RG_rl_18_t1 = TR_30 ;
	7'h4f :
		RG_rl_18_t1 = TR_30 ;
	7'h50 :
		RG_rl_18_t1 = TR_30 ;
	7'h51 :
		RG_rl_18_t1 = TR_30 ;
	7'h52 :
		RG_rl_18_t1 = TR_30 ;
	7'h53 :
		RG_rl_18_t1 = TR_30 ;
	7'h54 :
		RG_rl_18_t1 = TR_30 ;
	7'h55 :
		RG_rl_18_t1 = TR_30 ;
	7'h56 :
		RG_rl_18_t1 = TR_30 ;
	7'h57 :
		RG_rl_18_t1 = TR_30 ;
	7'h58 :
		RG_rl_18_t1 = TR_30 ;
	7'h59 :
		RG_rl_18_t1 = TR_30 ;
	7'h5a :
		RG_rl_18_t1 = TR_30 ;
	7'h5b :
		RG_rl_18_t1 = TR_30 ;
	7'h5c :
		RG_rl_18_t1 = TR_30 ;
	7'h5d :
		RG_rl_18_t1 = TR_30 ;
	7'h5e :
		RG_rl_18_t1 = TR_30 ;
	7'h5f :
		RG_rl_18_t1 = TR_30 ;
	7'h60 :
		RG_rl_18_t1 = TR_30 ;
	7'h61 :
		RG_rl_18_t1 = TR_30 ;
	7'h62 :
		RG_rl_18_t1 = TR_30 ;
	7'h63 :
		RG_rl_18_t1 = TR_30 ;
	7'h64 :
		RG_rl_18_t1 = TR_30 ;
	7'h65 :
		RG_rl_18_t1 = TR_30 ;
	7'h66 :
		RG_rl_18_t1 = TR_30 ;
	7'h67 :
		RG_rl_18_t1 = TR_30 ;
	7'h68 :
		RG_rl_18_t1 = TR_30 ;
	7'h69 :
		RG_rl_18_t1 = TR_30 ;
	7'h6a :
		RG_rl_18_t1 = TR_30 ;
	7'h6b :
		RG_rl_18_t1 = TR_30 ;
	7'h6c :
		RG_rl_18_t1 = TR_30 ;
	7'h6d :
		RG_rl_18_t1 = TR_30 ;
	7'h6e :
		RG_rl_18_t1 = TR_30 ;
	7'h6f :
		RG_rl_18_t1 = TR_30 ;
	7'h70 :
		RG_rl_18_t1 = TR_30 ;
	7'h71 :
		RG_rl_18_t1 = TR_30 ;
	7'h72 :
		RG_rl_18_t1 = TR_30 ;
	7'h73 :
		RG_rl_18_t1 = TR_30 ;
	7'h74 :
		RG_rl_18_t1 = TR_30 ;
	7'h75 :
		RG_rl_18_t1 = TR_30 ;
	7'h76 :
		RG_rl_18_t1 = TR_30 ;
	7'h77 :
		RG_rl_18_t1 = TR_30 ;
	7'h78 :
		RG_rl_18_t1 = TR_30 ;
	7'h79 :
		RG_rl_18_t1 = TR_30 ;
	7'h7a :
		RG_rl_18_t1 = TR_30 ;
	7'h7b :
		RG_rl_18_t1 = TR_30 ;
	7'h7c :
		RG_rl_18_t1 = TR_30 ;
	7'h7d :
		RG_rl_18_t1 = TR_30 ;
	7'h7e :
		RG_rl_18_t1 = TR_30 ;
	7'h7f :
		RG_rl_18_t1 = TR_30 ;
	default :
		RG_rl_18_t1 = 9'hx ;
	endcase
always @ ( RG_rl_18_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_201 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_18_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h12 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_18_t = ( ( { 9{ U_570 } } & RG_rl_201 )
		| ( { 9{ U_569 } } & RG_rl_18_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_18_en = ( U_570 | RG_rl_18_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_18_en )
		RG_rl_18 <= RG_rl_18_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_31 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_19_t1 = TR_31 ;
	7'h01 :
		RG_rl_19_t1 = TR_31 ;
	7'h02 :
		RG_rl_19_t1 = TR_31 ;
	7'h03 :
		RG_rl_19_t1 = TR_31 ;
	7'h04 :
		RG_rl_19_t1 = TR_31 ;
	7'h05 :
		RG_rl_19_t1 = TR_31 ;
	7'h06 :
		RG_rl_19_t1 = TR_31 ;
	7'h07 :
		RG_rl_19_t1 = TR_31 ;
	7'h08 :
		RG_rl_19_t1 = TR_31 ;
	7'h09 :
		RG_rl_19_t1 = TR_31 ;
	7'h0a :
		RG_rl_19_t1 = TR_31 ;
	7'h0b :
		RG_rl_19_t1 = TR_31 ;
	7'h0c :
		RG_rl_19_t1 = TR_31 ;
	7'h0d :
		RG_rl_19_t1 = TR_31 ;
	7'h0e :
		RG_rl_19_t1 = TR_31 ;
	7'h0f :
		RG_rl_19_t1 = TR_31 ;
	7'h10 :
		RG_rl_19_t1 = TR_31 ;
	7'h11 :
		RG_rl_19_t1 = TR_31 ;
	7'h12 :
		RG_rl_19_t1 = TR_31 ;
	7'h13 :
		RG_rl_19_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h14 :
		RG_rl_19_t1 = TR_31 ;
	7'h15 :
		RG_rl_19_t1 = TR_31 ;
	7'h16 :
		RG_rl_19_t1 = TR_31 ;
	7'h17 :
		RG_rl_19_t1 = TR_31 ;
	7'h18 :
		RG_rl_19_t1 = TR_31 ;
	7'h19 :
		RG_rl_19_t1 = TR_31 ;
	7'h1a :
		RG_rl_19_t1 = TR_31 ;
	7'h1b :
		RG_rl_19_t1 = TR_31 ;
	7'h1c :
		RG_rl_19_t1 = TR_31 ;
	7'h1d :
		RG_rl_19_t1 = TR_31 ;
	7'h1e :
		RG_rl_19_t1 = TR_31 ;
	7'h1f :
		RG_rl_19_t1 = TR_31 ;
	7'h20 :
		RG_rl_19_t1 = TR_31 ;
	7'h21 :
		RG_rl_19_t1 = TR_31 ;
	7'h22 :
		RG_rl_19_t1 = TR_31 ;
	7'h23 :
		RG_rl_19_t1 = TR_31 ;
	7'h24 :
		RG_rl_19_t1 = TR_31 ;
	7'h25 :
		RG_rl_19_t1 = TR_31 ;
	7'h26 :
		RG_rl_19_t1 = TR_31 ;
	7'h27 :
		RG_rl_19_t1 = TR_31 ;
	7'h28 :
		RG_rl_19_t1 = TR_31 ;
	7'h29 :
		RG_rl_19_t1 = TR_31 ;
	7'h2a :
		RG_rl_19_t1 = TR_31 ;
	7'h2b :
		RG_rl_19_t1 = TR_31 ;
	7'h2c :
		RG_rl_19_t1 = TR_31 ;
	7'h2d :
		RG_rl_19_t1 = TR_31 ;
	7'h2e :
		RG_rl_19_t1 = TR_31 ;
	7'h2f :
		RG_rl_19_t1 = TR_31 ;
	7'h30 :
		RG_rl_19_t1 = TR_31 ;
	7'h31 :
		RG_rl_19_t1 = TR_31 ;
	7'h32 :
		RG_rl_19_t1 = TR_31 ;
	7'h33 :
		RG_rl_19_t1 = TR_31 ;
	7'h34 :
		RG_rl_19_t1 = TR_31 ;
	7'h35 :
		RG_rl_19_t1 = TR_31 ;
	7'h36 :
		RG_rl_19_t1 = TR_31 ;
	7'h37 :
		RG_rl_19_t1 = TR_31 ;
	7'h38 :
		RG_rl_19_t1 = TR_31 ;
	7'h39 :
		RG_rl_19_t1 = TR_31 ;
	7'h3a :
		RG_rl_19_t1 = TR_31 ;
	7'h3b :
		RG_rl_19_t1 = TR_31 ;
	7'h3c :
		RG_rl_19_t1 = TR_31 ;
	7'h3d :
		RG_rl_19_t1 = TR_31 ;
	7'h3e :
		RG_rl_19_t1 = TR_31 ;
	7'h3f :
		RG_rl_19_t1 = TR_31 ;
	7'h40 :
		RG_rl_19_t1 = TR_31 ;
	7'h41 :
		RG_rl_19_t1 = TR_31 ;
	7'h42 :
		RG_rl_19_t1 = TR_31 ;
	7'h43 :
		RG_rl_19_t1 = TR_31 ;
	7'h44 :
		RG_rl_19_t1 = TR_31 ;
	7'h45 :
		RG_rl_19_t1 = TR_31 ;
	7'h46 :
		RG_rl_19_t1 = TR_31 ;
	7'h47 :
		RG_rl_19_t1 = TR_31 ;
	7'h48 :
		RG_rl_19_t1 = TR_31 ;
	7'h49 :
		RG_rl_19_t1 = TR_31 ;
	7'h4a :
		RG_rl_19_t1 = TR_31 ;
	7'h4b :
		RG_rl_19_t1 = TR_31 ;
	7'h4c :
		RG_rl_19_t1 = TR_31 ;
	7'h4d :
		RG_rl_19_t1 = TR_31 ;
	7'h4e :
		RG_rl_19_t1 = TR_31 ;
	7'h4f :
		RG_rl_19_t1 = TR_31 ;
	7'h50 :
		RG_rl_19_t1 = TR_31 ;
	7'h51 :
		RG_rl_19_t1 = TR_31 ;
	7'h52 :
		RG_rl_19_t1 = TR_31 ;
	7'h53 :
		RG_rl_19_t1 = TR_31 ;
	7'h54 :
		RG_rl_19_t1 = TR_31 ;
	7'h55 :
		RG_rl_19_t1 = TR_31 ;
	7'h56 :
		RG_rl_19_t1 = TR_31 ;
	7'h57 :
		RG_rl_19_t1 = TR_31 ;
	7'h58 :
		RG_rl_19_t1 = TR_31 ;
	7'h59 :
		RG_rl_19_t1 = TR_31 ;
	7'h5a :
		RG_rl_19_t1 = TR_31 ;
	7'h5b :
		RG_rl_19_t1 = TR_31 ;
	7'h5c :
		RG_rl_19_t1 = TR_31 ;
	7'h5d :
		RG_rl_19_t1 = TR_31 ;
	7'h5e :
		RG_rl_19_t1 = TR_31 ;
	7'h5f :
		RG_rl_19_t1 = TR_31 ;
	7'h60 :
		RG_rl_19_t1 = TR_31 ;
	7'h61 :
		RG_rl_19_t1 = TR_31 ;
	7'h62 :
		RG_rl_19_t1 = TR_31 ;
	7'h63 :
		RG_rl_19_t1 = TR_31 ;
	7'h64 :
		RG_rl_19_t1 = TR_31 ;
	7'h65 :
		RG_rl_19_t1 = TR_31 ;
	7'h66 :
		RG_rl_19_t1 = TR_31 ;
	7'h67 :
		RG_rl_19_t1 = TR_31 ;
	7'h68 :
		RG_rl_19_t1 = TR_31 ;
	7'h69 :
		RG_rl_19_t1 = TR_31 ;
	7'h6a :
		RG_rl_19_t1 = TR_31 ;
	7'h6b :
		RG_rl_19_t1 = TR_31 ;
	7'h6c :
		RG_rl_19_t1 = TR_31 ;
	7'h6d :
		RG_rl_19_t1 = TR_31 ;
	7'h6e :
		RG_rl_19_t1 = TR_31 ;
	7'h6f :
		RG_rl_19_t1 = TR_31 ;
	7'h70 :
		RG_rl_19_t1 = TR_31 ;
	7'h71 :
		RG_rl_19_t1 = TR_31 ;
	7'h72 :
		RG_rl_19_t1 = TR_31 ;
	7'h73 :
		RG_rl_19_t1 = TR_31 ;
	7'h74 :
		RG_rl_19_t1 = TR_31 ;
	7'h75 :
		RG_rl_19_t1 = TR_31 ;
	7'h76 :
		RG_rl_19_t1 = TR_31 ;
	7'h77 :
		RG_rl_19_t1 = TR_31 ;
	7'h78 :
		RG_rl_19_t1 = TR_31 ;
	7'h79 :
		RG_rl_19_t1 = TR_31 ;
	7'h7a :
		RG_rl_19_t1 = TR_31 ;
	7'h7b :
		RG_rl_19_t1 = TR_31 ;
	7'h7c :
		RG_rl_19_t1 = TR_31 ;
	7'h7d :
		RG_rl_19_t1 = TR_31 ;
	7'h7e :
		RG_rl_19_t1 = TR_31 ;
	7'h7f :
		RG_rl_19_t1 = TR_31 ;
	default :
		RG_rl_19_t1 = 9'hx ;
	endcase
always @ ( RG_rl_19_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_202 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_19_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h13 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_19_t = ( ( { 9{ U_570 } } & RG_rl_202 )
		| ( { 9{ U_569 } } & RG_rl_19_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_19_en = ( U_570 | RG_rl_19_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_19_en )
		RG_rl_19 <= RG_rl_19_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_32 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_20_t1 = TR_32 ;
	7'h01 :
		RG_rl_20_t1 = TR_32 ;
	7'h02 :
		RG_rl_20_t1 = TR_32 ;
	7'h03 :
		RG_rl_20_t1 = TR_32 ;
	7'h04 :
		RG_rl_20_t1 = TR_32 ;
	7'h05 :
		RG_rl_20_t1 = TR_32 ;
	7'h06 :
		RG_rl_20_t1 = TR_32 ;
	7'h07 :
		RG_rl_20_t1 = TR_32 ;
	7'h08 :
		RG_rl_20_t1 = TR_32 ;
	7'h09 :
		RG_rl_20_t1 = TR_32 ;
	7'h0a :
		RG_rl_20_t1 = TR_32 ;
	7'h0b :
		RG_rl_20_t1 = TR_32 ;
	7'h0c :
		RG_rl_20_t1 = TR_32 ;
	7'h0d :
		RG_rl_20_t1 = TR_32 ;
	7'h0e :
		RG_rl_20_t1 = TR_32 ;
	7'h0f :
		RG_rl_20_t1 = TR_32 ;
	7'h10 :
		RG_rl_20_t1 = TR_32 ;
	7'h11 :
		RG_rl_20_t1 = TR_32 ;
	7'h12 :
		RG_rl_20_t1 = TR_32 ;
	7'h13 :
		RG_rl_20_t1 = TR_32 ;
	7'h14 :
		RG_rl_20_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h15 :
		RG_rl_20_t1 = TR_32 ;
	7'h16 :
		RG_rl_20_t1 = TR_32 ;
	7'h17 :
		RG_rl_20_t1 = TR_32 ;
	7'h18 :
		RG_rl_20_t1 = TR_32 ;
	7'h19 :
		RG_rl_20_t1 = TR_32 ;
	7'h1a :
		RG_rl_20_t1 = TR_32 ;
	7'h1b :
		RG_rl_20_t1 = TR_32 ;
	7'h1c :
		RG_rl_20_t1 = TR_32 ;
	7'h1d :
		RG_rl_20_t1 = TR_32 ;
	7'h1e :
		RG_rl_20_t1 = TR_32 ;
	7'h1f :
		RG_rl_20_t1 = TR_32 ;
	7'h20 :
		RG_rl_20_t1 = TR_32 ;
	7'h21 :
		RG_rl_20_t1 = TR_32 ;
	7'h22 :
		RG_rl_20_t1 = TR_32 ;
	7'h23 :
		RG_rl_20_t1 = TR_32 ;
	7'h24 :
		RG_rl_20_t1 = TR_32 ;
	7'h25 :
		RG_rl_20_t1 = TR_32 ;
	7'h26 :
		RG_rl_20_t1 = TR_32 ;
	7'h27 :
		RG_rl_20_t1 = TR_32 ;
	7'h28 :
		RG_rl_20_t1 = TR_32 ;
	7'h29 :
		RG_rl_20_t1 = TR_32 ;
	7'h2a :
		RG_rl_20_t1 = TR_32 ;
	7'h2b :
		RG_rl_20_t1 = TR_32 ;
	7'h2c :
		RG_rl_20_t1 = TR_32 ;
	7'h2d :
		RG_rl_20_t1 = TR_32 ;
	7'h2e :
		RG_rl_20_t1 = TR_32 ;
	7'h2f :
		RG_rl_20_t1 = TR_32 ;
	7'h30 :
		RG_rl_20_t1 = TR_32 ;
	7'h31 :
		RG_rl_20_t1 = TR_32 ;
	7'h32 :
		RG_rl_20_t1 = TR_32 ;
	7'h33 :
		RG_rl_20_t1 = TR_32 ;
	7'h34 :
		RG_rl_20_t1 = TR_32 ;
	7'h35 :
		RG_rl_20_t1 = TR_32 ;
	7'h36 :
		RG_rl_20_t1 = TR_32 ;
	7'h37 :
		RG_rl_20_t1 = TR_32 ;
	7'h38 :
		RG_rl_20_t1 = TR_32 ;
	7'h39 :
		RG_rl_20_t1 = TR_32 ;
	7'h3a :
		RG_rl_20_t1 = TR_32 ;
	7'h3b :
		RG_rl_20_t1 = TR_32 ;
	7'h3c :
		RG_rl_20_t1 = TR_32 ;
	7'h3d :
		RG_rl_20_t1 = TR_32 ;
	7'h3e :
		RG_rl_20_t1 = TR_32 ;
	7'h3f :
		RG_rl_20_t1 = TR_32 ;
	7'h40 :
		RG_rl_20_t1 = TR_32 ;
	7'h41 :
		RG_rl_20_t1 = TR_32 ;
	7'h42 :
		RG_rl_20_t1 = TR_32 ;
	7'h43 :
		RG_rl_20_t1 = TR_32 ;
	7'h44 :
		RG_rl_20_t1 = TR_32 ;
	7'h45 :
		RG_rl_20_t1 = TR_32 ;
	7'h46 :
		RG_rl_20_t1 = TR_32 ;
	7'h47 :
		RG_rl_20_t1 = TR_32 ;
	7'h48 :
		RG_rl_20_t1 = TR_32 ;
	7'h49 :
		RG_rl_20_t1 = TR_32 ;
	7'h4a :
		RG_rl_20_t1 = TR_32 ;
	7'h4b :
		RG_rl_20_t1 = TR_32 ;
	7'h4c :
		RG_rl_20_t1 = TR_32 ;
	7'h4d :
		RG_rl_20_t1 = TR_32 ;
	7'h4e :
		RG_rl_20_t1 = TR_32 ;
	7'h4f :
		RG_rl_20_t1 = TR_32 ;
	7'h50 :
		RG_rl_20_t1 = TR_32 ;
	7'h51 :
		RG_rl_20_t1 = TR_32 ;
	7'h52 :
		RG_rl_20_t1 = TR_32 ;
	7'h53 :
		RG_rl_20_t1 = TR_32 ;
	7'h54 :
		RG_rl_20_t1 = TR_32 ;
	7'h55 :
		RG_rl_20_t1 = TR_32 ;
	7'h56 :
		RG_rl_20_t1 = TR_32 ;
	7'h57 :
		RG_rl_20_t1 = TR_32 ;
	7'h58 :
		RG_rl_20_t1 = TR_32 ;
	7'h59 :
		RG_rl_20_t1 = TR_32 ;
	7'h5a :
		RG_rl_20_t1 = TR_32 ;
	7'h5b :
		RG_rl_20_t1 = TR_32 ;
	7'h5c :
		RG_rl_20_t1 = TR_32 ;
	7'h5d :
		RG_rl_20_t1 = TR_32 ;
	7'h5e :
		RG_rl_20_t1 = TR_32 ;
	7'h5f :
		RG_rl_20_t1 = TR_32 ;
	7'h60 :
		RG_rl_20_t1 = TR_32 ;
	7'h61 :
		RG_rl_20_t1 = TR_32 ;
	7'h62 :
		RG_rl_20_t1 = TR_32 ;
	7'h63 :
		RG_rl_20_t1 = TR_32 ;
	7'h64 :
		RG_rl_20_t1 = TR_32 ;
	7'h65 :
		RG_rl_20_t1 = TR_32 ;
	7'h66 :
		RG_rl_20_t1 = TR_32 ;
	7'h67 :
		RG_rl_20_t1 = TR_32 ;
	7'h68 :
		RG_rl_20_t1 = TR_32 ;
	7'h69 :
		RG_rl_20_t1 = TR_32 ;
	7'h6a :
		RG_rl_20_t1 = TR_32 ;
	7'h6b :
		RG_rl_20_t1 = TR_32 ;
	7'h6c :
		RG_rl_20_t1 = TR_32 ;
	7'h6d :
		RG_rl_20_t1 = TR_32 ;
	7'h6e :
		RG_rl_20_t1 = TR_32 ;
	7'h6f :
		RG_rl_20_t1 = TR_32 ;
	7'h70 :
		RG_rl_20_t1 = TR_32 ;
	7'h71 :
		RG_rl_20_t1 = TR_32 ;
	7'h72 :
		RG_rl_20_t1 = TR_32 ;
	7'h73 :
		RG_rl_20_t1 = TR_32 ;
	7'h74 :
		RG_rl_20_t1 = TR_32 ;
	7'h75 :
		RG_rl_20_t1 = TR_32 ;
	7'h76 :
		RG_rl_20_t1 = TR_32 ;
	7'h77 :
		RG_rl_20_t1 = TR_32 ;
	7'h78 :
		RG_rl_20_t1 = TR_32 ;
	7'h79 :
		RG_rl_20_t1 = TR_32 ;
	7'h7a :
		RG_rl_20_t1 = TR_32 ;
	7'h7b :
		RG_rl_20_t1 = TR_32 ;
	7'h7c :
		RG_rl_20_t1 = TR_32 ;
	7'h7d :
		RG_rl_20_t1 = TR_32 ;
	7'h7e :
		RG_rl_20_t1 = TR_32 ;
	7'h7f :
		RG_rl_20_t1 = TR_32 ;
	default :
		RG_rl_20_t1 = 9'hx ;
	endcase
always @ ( RG_rl_20_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_203 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_20_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h14 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_20_t = ( ( { 9{ U_570 } } & RG_rl_203 )
		| ( { 9{ U_569 } } & RG_rl_20_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_20_en = ( U_570 | RG_rl_20_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_20_en )
		RG_rl_20 <= RG_rl_20_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_33 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_21_t1 = TR_33 ;
	7'h01 :
		RG_rl_21_t1 = TR_33 ;
	7'h02 :
		RG_rl_21_t1 = TR_33 ;
	7'h03 :
		RG_rl_21_t1 = TR_33 ;
	7'h04 :
		RG_rl_21_t1 = TR_33 ;
	7'h05 :
		RG_rl_21_t1 = TR_33 ;
	7'h06 :
		RG_rl_21_t1 = TR_33 ;
	7'h07 :
		RG_rl_21_t1 = TR_33 ;
	7'h08 :
		RG_rl_21_t1 = TR_33 ;
	7'h09 :
		RG_rl_21_t1 = TR_33 ;
	7'h0a :
		RG_rl_21_t1 = TR_33 ;
	7'h0b :
		RG_rl_21_t1 = TR_33 ;
	7'h0c :
		RG_rl_21_t1 = TR_33 ;
	7'h0d :
		RG_rl_21_t1 = TR_33 ;
	7'h0e :
		RG_rl_21_t1 = TR_33 ;
	7'h0f :
		RG_rl_21_t1 = TR_33 ;
	7'h10 :
		RG_rl_21_t1 = TR_33 ;
	7'h11 :
		RG_rl_21_t1 = TR_33 ;
	7'h12 :
		RG_rl_21_t1 = TR_33 ;
	7'h13 :
		RG_rl_21_t1 = TR_33 ;
	7'h14 :
		RG_rl_21_t1 = TR_33 ;
	7'h15 :
		RG_rl_21_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h16 :
		RG_rl_21_t1 = TR_33 ;
	7'h17 :
		RG_rl_21_t1 = TR_33 ;
	7'h18 :
		RG_rl_21_t1 = TR_33 ;
	7'h19 :
		RG_rl_21_t1 = TR_33 ;
	7'h1a :
		RG_rl_21_t1 = TR_33 ;
	7'h1b :
		RG_rl_21_t1 = TR_33 ;
	7'h1c :
		RG_rl_21_t1 = TR_33 ;
	7'h1d :
		RG_rl_21_t1 = TR_33 ;
	7'h1e :
		RG_rl_21_t1 = TR_33 ;
	7'h1f :
		RG_rl_21_t1 = TR_33 ;
	7'h20 :
		RG_rl_21_t1 = TR_33 ;
	7'h21 :
		RG_rl_21_t1 = TR_33 ;
	7'h22 :
		RG_rl_21_t1 = TR_33 ;
	7'h23 :
		RG_rl_21_t1 = TR_33 ;
	7'h24 :
		RG_rl_21_t1 = TR_33 ;
	7'h25 :
		RG_rl_21_t1 = TR_33 ;
	7'h26 :
		RG_rl_21_t1 = TR_33 ;
	7'h27 :
		RG_rl_21_t1 = TR_33 ;
	7'h28 :
		RG_rl_21_t1 = TR_33 ;
	7'h29 :
		RG_rl_21_t1 = TR_33 ;
	7'h2a :
		RG_rl_21_t1 = TR_33 ;
	7'h2b :
		RG_rl_21_t1 = TR_33 ;
	7'h2c :
		RG_rl_21_t1 = TR_33 ;
	7'h2d :
		RG_rl_21_t1 = TR_33 ;
	7'h2e :
		RG_rl_21_t1 = TR_33 ;
	7'h2f :
		RG_rl_21_t1 = TR_33 ;
	7'h30 :
		RG_rl_21_t1 = TR_33 ;
	7'h31 :
		RG_rl_21_t1 = TR_33 ;
	7'h32 :
		RG_rl_21_t1 = TR_33 ;
	7'h33 :
		RG_rl_21_t1 = TR_33 ;
	7'h34 :
		RG_rl_21_t1 = TR_33 ;
	7'h35 :
		RG_rl_21_t1 = TR_33 ;
	7'h36 :
		RG_rl_21_t1 = TR_33 ;
	7'h37 :
		RG_rl_21_t1 = TR_33 ;
	7'h38 :
		RG_rl_21_t1 = TR_33 ;
	7'h39 :
		RG_rl_21_t1 = TR_33 ;
	7'h3a :
		RG_rl_21_t1 = TR_33 ;
	7'h3b :
		RG_rl_21_t1 = TR_33 ;
	7'h3c :
		RG_rl_21_t1 = TR_33 ;
	7'h3d :
		RG_rl_21_t1 = TR_33 ;
	7'h3e :
		RG_rl_21_t1 = TR_33 ;
	7'h3f :
		RG_rl_21_t1 = TR_33 ;
	7'h40 :
		RG_rl_21_t1 = TR_33 ;
	7'h41 :
		RG_rl_21_t1 = TR_33 ;
	7'h42 :
		RG_rl_21_t1 = TR_33 ;
	7'h43 :
		RG_rl_21_t1 = TR_33 ;
	7'h44 :
		RG_rl_21_t1 = TR_33 ;
	7'h45 :
		RG_rl_21_t1 = TR_33 ;
	7'h46 :
		RG_rl_21_t1 = TR_33 ;
	7'h47 :
		RG_rl_21_t1 = TR_33 ;
	7'h48 :
		RG_rl_21_t1 = TR_33 ;
	7'h49 :
		RG_rl_21_t1 = TR_33 ;
	7'h4a :
		RG_rl_21_t1 = TR_33 ;
	7'h4b :
		RG_rl_21_t1 = TR_33 ;
	7'h4c :
		RG_rl_21_t1 = TR_33 ;
	7'h4d :
		RG_rl_21_t1 = TR_33 ;
	7'h4e :
		RG_rl_21_t1 = TR_33 ;
	7'h4f :
		RG_rl_21_t1 = TR_33 ;
	7'h50 :
		RG_rl_21_t1 = TR_33 ;
	7'h51 :
		RG_rl_21_t1 = TR_33 ;
	7'h52 :
		RG_rl_21_t1 = TR_33 ;
	7'h53 :
		RG_rl_21_t1 = TR_33 ;
	7'h54 :
		RG_rl_21_t1 = TR_33 ;
	7'h55 :
		RG_rl_21_t1 = TR_33 ;
	7'h56 :
		RG_rl_21_t1 = TR_33 ;
	7'h57 :
		RG_rl_21_t1 = TR_33 ;
	7'h58 :
		RG_rl_21_t1 = TR_33 ;
	7'h59 :
		RG_rl_21_t1 = TR_33 ;
	7'h5a :
		RG_rl_21_t1 = TR_33 ;
	7'h5b :
		RG_rl_21_t1 = TR_33 ;
	7'h5c :
		RG_rl_21_t1 = TR_33 ;
	7'h5d :
		RG_rl_21_t1 = TR_33 ;
	7'h5e :
		RG_rl_21_t1 = TR_33 ;
	7'h5f :
		RG_rl_21_t1 = TR_33 ;
	7'h60 :
		RG_rl_21_t1 = TR_33 ;
	7'h61 :
		RG_rl_21_t1 = TR_33 ;
	7'h62 :
		RG_rl_21_t1 = TR_33 ;
	7'h63 :
		RG_rl_21_t1 = TR_33 ;
	7'h64 :
		RG_rl_21_t1 = TR_33 ;
	7'h65 :
		RG_rl_21_t1 = TR_33 ;
	7'h66 :
		RG_rl_21_t1 = TR_33 ;
	7'h67 :
		RG_rl_21_t1 = TR_33 ;
	7'h68 :
		RG_rl_21_t1 = TR_33 ;
	7'h69 :
		RG_rl_21_t1 = TR_33 ;
	7'h6a :
		RG_rl_21_t1 = TR_33 ;
	7'h6b :
		RG_rl_21_t1 = TR_33 ;
	7'h6c :
		RG_rl_21_t1 = TR_33 ;
	7'h6d :
		RG_rl_21_t1 = TR_33 ;
	7'h6e :
		RG_rl_21_t1 = TR_33 ;
	7'h6f :
		RG_rl_21_t1 = TR_33 ;
	7'h70 :
		RG_rl_21_t1 = TR_33 ;
	7'h71 :
		RG_rl_21_t1 = TR_33 ;
	7'h72 :
		RG_rl_21_t1 = TR_33 ;
	7'h73 :
		RG_rl_21_t1 = TR_33 ;
	7'h74 :
		RG_rl_21_t1 = TR_33 ;
	7'h75 :
		RG_rl_21_t1 = TR_33 ;
	7'h76 :
		RG_rl_21_t1 = TR_33 ;
	7'h77 :
		RG_rl_21_t1 = TR_33 ;
	7'h78 :
		RG_rl_21_t1 = TR_33 ;
	7'h79 :
		RG_rl_21_t1 = TR_33 ;
	7'h7a :
		RG_rl_21_t1 = TR_33 ;
	7'h7b :
		RG_rl_21_t1 = TR_33 ;
	7'h7c :
		RG_rl_21_t1 = TR_33 ;
	7'h7d :
		RG_rl_21_t1 = TR_33 ;
	7'h7e :
		RG_rl_21_t1 = TR_33 ;
	7'h7f :
		RG_rl_21_t1 = TR_33 ;
	default :
		RG_rl_21_t1 = 9'hx ;
	endcase
always @ ( RG_rl_21_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_204 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_21_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h15 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_21_t = ( ( { 9{ U_570 } } & RG_rl_204 )
		| ( { 9{ U_569 } } & RG_rl_21_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_21_en = ( U_570 | RG_rl_21_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_21_en )
		RG_rl_21 <= RG_rl_21_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_34 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_22_t1 = TR_34 ;
	7'h01 :
		RG_rl_22_t1 = TR_34 ;
	7'h02 :
		RG_rl_22_t1 = TR_34 ;
	7'h03 :
		RG_rl_22_t1 = TR_34 ;
	7'h04 :
		RG_rl_22_t1 = TR_34 ;
	7'h05 :
		RG_rl_22_t1 = TR_34 ;
	7'h06 :
		RG_rl_22_t1 = TR_34 ;
	7'h07 :
		RG_rl_22_t1 = TR_34 ;
	7'h08 :
		RG_rl_22_t1 = TR_34 ;
	7'h09 :
		RG_rl_22_t1 = TR_34 ;
	7'h0a :
		RG_rl_22_t1 = TR_34 ;
	7'h0b :
		RG_rl_22_t1 = TR_34 ;
	7'h0c :
		RG_rl_22_t1 = TR_34 ;
	7'h0d :
		RG_rl_22_t1 = TR_34 ;
	7'h0e :
		RG_rl_22_t1 = TR_34 ;
	7'h0f :
		RG_rl_22_t1 = TR_34 ;
	7'h10 :
		RG_rl_22_t1 = TR_34 ;
	7'h11 :
		RG_rl_22_t1 = TR_34 ;
	7'h12 :
		RG_rl_22_t1 = TR_34 ;
	7'h13 :
		RG_rl_22_t1 = TR_34 ;
	7'h14 :
		RG_rl_22_t1 = TR_34 ;
	7'h15 :
		RG_rl_22_t1 = TR_34 ;
	7'h16 :
		RG_rl_22_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h17 :
		RG_rl_22_t1 = TR_34 ;
	7'h18 :
		RG_rl_22_t1 = TR_34 ;
	7'h19 :
		RG_rl_22_t1 = TR_34 ;
	7'h1a :
		RG_rl_22_t1 = TR_34 ;
	7'h1b :
		RG_rl_22_t1 = TR_34 ;
	7'h1c :
		RG_rl_22_t1 = TR_34 ;
	7'h1d :
		RG_rl_22_t1 = TR_34 ;
	7'h1e :
		RG_rl_22_t1 = TR_34 ;
	7'h1f :
		RG_rl_22_t1 = TR_34 ;
	7'h20 :
		RG_rl_22_t1 = TR_34 ;
	7'h21 :
		RG_rl_22_t1 = TR_34 ;
	7'h22 :
		RG_rl_22_t1 = TR_34 ;
	7'h23 :
		RG_rl_22_t1 = TR_34 ;
	7'h24 :
		RG_rl_22_t1 = TR_34 ;
	7'h25 :
		RG_rl_22_t1 = TR_34 ;
	7'h26 :
		RG_rl_22_t1 = TR_34 ;
	7'h27 :
		RG_rl_22_t1 = TR_34 ;
	7'h28 :
		RG_rl_22_t1 = TR_34 ;
	7'h29 :
		RG_rl_22_t1 = TR_34 ;
	7'h2a :
		RG_rl_22_t1 = TR_34 ;
	7'h2b :
		RG_rl_22_t1 = TR_34 ;
	7'h2c :
		RG_rl_22_t1 = TR_34 ;
	7'h2d :
		RG_rl_22_t1 = TR_34 ;
	7'h2e :
		RG_rl_22_t1 = TR_34 ;
	7'h2f :
		RG_rl_22_t1 = TR_34 ;
	7'h30 :
		RG_rl_22_t1 = TR_34 ;
	7'h31 :
		RG_rl_22_t1 = TR_34 ;
	7'h32 :
		RG_rl_22_t1 = TR_34 ;
	7'h33 :
		RG_rl_22_t1 = TR_34 ;
	7'h34 :
		RG_rl_22_t1 = TR_34 ;
	7'h35 :
		RG_rl_22_t1 = TR_34 ;
	7'h36 :
		RG_rl_22_t1 = TR_34 ;
	7'h37 :
		RG_rl_22_t1 = TR_34 ;
	7'h38 :
		RG_rl_22_t1 = TR_34 ;
	7'h39 :
		RG_rl_22_t1 = TR_34 ;
	7'h3a :
		RG_rl_22_t1 = TR_34 ;
	7'h3b :
		RG_rl_22_t1 = TR_34 ;
	7'h3c :
		RG_rl_22_t1 = TR_34 ;
	7'h3d :
		RG_rl_22_t1 = TR_34 ;
	7'h3e :
		RG_rl_22_t1 = TR_34 ;
	7'h3f :
		RG_rl_22_t1 = TR_34 ;
	7'h40 :
		RG_rl_22_t1 = TR_34 ;
	7'h41 :
		RG_rl_22_t1 = TR_34 ;
	7'h42 :
		RG_rl_22_t1 = TR_34 ;
	7'h43 :
		RG_rl_22_t1 = TR_34 ;
	7'h44 :
		RG_rl_22_t1 = TR_34 ;
	7'h45 :
		RG_rl_22_t1 = TR_34 ;
	7'h46 :
		RG_rl_22_t1 = TR_34 ;
	7'h47 :
		RG_rl_22_t1 = TR_34 ;
	7'h48 :
		RG_rl_22_t1 = TR_34 ;
	7'h49 :
		RG_rl_22_t1 = TR_34 ;
	7'h4a :
		RG_rl_22_t1 = TR_34 ;
	7'h4b :
		RG_rl_22_t1 = TR_34 ;
	7'h4c :
		RG_rl_22_t1 = TR_34 ;
	7'h4d :
		RG_rl_22_t1 = TR_34 ;
	7'h4e :
		RG_rl_22_t1 = TR_34 ;
	7'h4f :
		RG_rl_22_t1 = TR_34 ;
	7'h50 :
		RG_rl_22_t1 = TR_34 ;
	7'h51 :
		RG_rl_22_t1 = TR_34 ;
	7'h52 :
		RG_rl_22_t1 = TR_34 ;
	7'h53 :
		RG_rl_22_t1 = TR_34 ;
	7'h54 :
		RG_rl_22_t1 = TR_34 ;
	7'h55 :
		RG_rl_22_t1 = TR_34 ;
	7'h56 :
		RG_rl_22_t1 = TR_34 ;
	7'h57 :
		RG_rl_22_t1 = TR_34 ;
	7'h58 :
		RG_rl_22_t1 = TR_34 ;
	7'h59 :
		RG_rl_22_t1 = TR_34 ;
	7'h5a :
		RG_rl_22_t1 = TR_34 ;
	7'h5b :
		RG_rl_22_t1 = TR_34 ;
	7'h5c :
		RG_rl_22_t1 = TR_34 ;
	7'h5d :
		RG_rl_22_t1 = TR_34 ;
	7'h5e :
		RG_rl_22_t1 = TR_34 ;
	7'h5f :
		RG_rl_22_t1 = TR_34 ;
	7'h60 :
		RG_rl_22_t1 = TR_34 ;
	7'h61 :
		RG_rl_22_t1 = TR_34 ;
	7'h62 :
		RG_rl_22_t1 = TR_34 ;
	7'h63 :
		RG_rl_22_t1 = TR_34 ;
	7'h64 :
		RG_rl_22_t1 = TR_34 ;
	7'h65 :
		RG_rl_22_t1 = TR_34 ;
	7'h66 :
		RG_rl_22_t1 = TR_34 ;
	7'h67 :
		RG_rl_22_t1 = TR_34 ;
	7'h68 :
		RG_rl_22_t1 = TR_34 ;
	7'h69 :
		RG_rl_22_t1 = TR_34 ;
	7'h6a :
		RG_rl_22_t1 = TR_34 ;
	7'h6b :
		RG_rl_22_t1 = TR_34 ;
	7'h6c :
		RG_rl_22_t1 = TR_34 ;
	7'h6d :
		RG_rl_22_t1 = TR_34 ;
	7'h6e :
		RG_rl_22_t1 = TR_34 ;
	7'h6f :
		RG_rl_22_t1 = TR_34 ;
	7'h70 :
		RG_rl_22_t1 = TR_34 ;
	7'h71 :
		RG_rl_22_t1 = TR_34 ;
	7'h72 :
		RG_rl_22_t1 = TR_34 ;
	7'h73 :
		RG_rl_22_t1 = TR_34 ;
	7'h74 :
		RG_rl_22_t1 = TR_34 ;
	7'h75 :
		RG_rl_22_t1 = TR_34 ;
	7'h76 :
		RG_rl_22_t1 = TR_34 ;
	7'h77 :
		RG_rl_22_t1 = TR_34 ;
	7'h78 :
		RG_rl_22_t1 = TR_34 ;
	7'h79 :
		RG_rl_22_t1 = TR_34 ;
	7'h7a :
		RG_rl_22_t1 = TR_34 ;
	7'h7b :
		RG_rl_22_t1 = TR_34 ;
	7'h7c :
		RG_rl_22_t1 = TR_34 ;
	7'h7d :
		RG_rl_22_t1 = TR_34 ;
	7'h7e :
		RG_rl_22_t1 = TR_34 ;
	7'h7f :
		RG_rl_22_t1 = TR_34 ;
	default :
		RG_rl_22_t1 = 9'hx ;
	endcase
always @ ( RG_rl_22_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_205 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_22_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h16 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_22_t = ( ( { 9{ U_570 } } & RG_rl_205 )
		| ( { 9{ U_569 } } & RG_rl_22_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_22_en = ( U_570 | RG_rl_22_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_22_en )
		RG_rl_22 <= RG_rl_22_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_35 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_23_t1 = TR_35 ;
	7'h01 :
		RG_rl_23_t1 = TR_35 ;
	7'h02 :
		RG_rl_23_t1 = TR_35 ;
	7'h03 :
		RG_rl_23_t1 = TR_35 ;
	7'h04 :
		RG_rl_23_t1 = TR_35 ;
	7'h05 :
		RG_rl_23_t1 = TR_35 ;
	7'h06 :
		RG_rl_23_t1 = TR_35 ;
	7'h07 :
		RG_rl_23_t1 = TR_35 ;
	7'h08 :
		RG_rl_23_t1 = TR_35 ;
	7'h09 :
		RG_rl_23_t1 = TR_35 ;
	7'h0a :
		RG_rl_23_t1 = TR_35 ;
	7'h0b :
		RG_rl_23_t1 = TR_35 ;
	7'h0c :
		RG_rl_23_t1 = TR_35 ;
	7'h0d :
		RG_rl_23_t1 = TR_35 ;
	7'h0e :
		RG_rl_23_t1 = TR_35 ;
	7'h0f :
		RG_rl_23_t1 = TR_35 ;
	7'h10 :
		RG_rl_23_t1 = TR_35 ;
	7'h11 :
		RG_rl_23_t1 = TR_35 ;
	7'h12 :
		RG_rl_23_t1 = TR_35 ;
	7'h13 :
		RG_rl_23_t1 = TR_35 ;
	7'h14 :
		RG_rl_23_t1 = TR_35 ;
	7'h15 :
		RG_rl_23_t1 = TR_35 ;
	7'h16 :
		RG_rl_23_t1 = TR_35 ;
	7'h17 :
		RG_rl_23_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h18 :
		RG_rl_23_t1 = TR_35 ;
	7'h19 :
		RG_rl_23_t1 = TR_35 ;
	7'h1a :
		RG_rl_23_t1 = TR_35 ;
	7'h1b :
		RG_rl_23_t1 = TR_35 ;
	7'h1c :
		RG_rl_23_t1 = TR_35 ;
	7'h1d :
		RG_rl_23_t1 = TR_35 ;
	7'h1e :
		RG_rl_23_t1 = TR_35 ;
	7'h1f :
		RG_rl_23_t1 = TR_35 ;
	7'h20 :
		RG_rl_23_t1 = TR_35 ;
	7'h21 :
		RG_rl_23_t1 = TR_35 ;
	7'h22 :
		RG_rl_23_t1 = TR_35 ;
	7'h23 :
		RG_rl_23_t1 = TR_35 ;
	7'h24 :
		RG_rl_23_t1 = TR_35 ;
	7'h25 :
		RG_rl_23_t1 = TR_35 ;
	7'h26 :
		RG_rl_23_t1 = TR_35 ;
	7'h27 :
		RG_rl_23_t1 = TR_35 ;
	7'h28 :
		RG_rl_23_t1 = TR_35 ;
	7'h29 :
		RG_rl_23_t1 = TR_35 ;
	7'h2a :
		RG_rl_23_t1 = TR_35 ;
	7'h2b :
		RG_rl_23_t1 = TR_35 ;
	7'h2c :
		RG_rl_23_t1 = TR_35 ;
	7'h2d :
		RG_rl_23_t1 = TR_35 ;
	7'h2e :
		RG_rl_23_t1 = TR_35 ;
	7'h2f :
		RG_rl_23_t1 = TR_35 ;
	7'h30 :
		RG_rl_23_t1 = TR_35 ;
	7'h31 :
		RG_rl_23_t1 = TR_35 ;
	7'h32 :
		RG_rl_23_t1 = TR_35 ;
	7'h33 :
		RG_rl_23_t1 = TR_35 ;
	7'h34 :
		RG_rl_23_t1 = TR_35 ;
	7'h35 :
		RG_rl_23_t1 = TR_35 ;
	7'h36 :
		RG_rl_23_t1 = TR_35 ;
	7'h37 :
		RG_rl_23_t1 = TR_35 ;
	7'h38 :
		RG_rl_23_t1 = TR_35 ;
	7'h39 :
		RG_rl_23_t1 = TR_35 ;
	7'h3a :
		RG_rl_23_t1 = TR_35 ;
	7'h3b :
		RG_rl_23_t1 = TR_35 ;
	7'h3c :
		RG_rl_23_t1 = TR_35 ;
	7'h3d :
		RG_rl_23_t1 = TR_35 ;
	7'h3e :
		RG_rl_23_t1 = TR_35 ;
	7'h3f :
		RG_rl_23_t1 = TR_35 ;
	7'h40 :
		RG_rl_23_t1 = TR_35 ;
	7'h41 :
		RG_rl_23_t1 = TR_35 ;
	7'h42 :
		RG_rl_23_t1 = TR_35 ;
	7'h43 :
		RG_rl_23_t1 = TR_35 ;
	7'h44 :
		RG_rl_23_t1 = TR_35 ;
	7'h45 :
		RG_rl_23_t1 = TR_35 ;
	7'h46 :
		RG_rl_23_t1 = TR_35 ;
	7'h47 :
		RG_rl_23_t1 = TR_35 ;
	7'h48 :
		RG_rl_23_t1 = TR_35 ;
	7'h49 :
		RG_rl_23_t1 = TR_35 ;
	7'h4a :
		RG_rl_23_t1 = TR_35 ;
	7'h4b :
		RG_rl_23_t1 = TR_35 ;
	7'h4c :
		RG_rl_23_t1 = TR_35 ;
	7'h4d :
		RG_rl_23_t1 = TR_35 ;
	7'h4e :
		RG_rl_23_t1 = TR_35 ;
	7'h4f :
		RG_rl_23_t1 = TR_35 ;
	7'h50 :
		RG_rl_23_t1 = TR_35 ;
	7'h51 :
		RG_rl_23_t1 = TR_35 ;
	7'h52 :
		RG_rl_23_t1 = TR_35 ;
	7'h53 :
		RG_rl_23_t1 = TR_35 ;
	7'h54 :
		RG_rl_23_t1 = TR_35 ;
	7'h55 :
		RG_rl_23_t1 = TR_35 ;
	7'h56 :
		RG_rl_23_t1 = TR_35 ;
	7'h57 :
		RG_rl_23_t1 = TR_35 ;
	7'h58 :
		RG_rl_23_t1 = TR_35 ;
	7'h59 :
		RG_rl_23_t1 = TR_35 ;
	7'h5a :
		RG_rl_23_t1 = TR_35 ;
	7'h5b :
		RG_rl_23_t1 = TR_35 ;
	7'h5c :
		RG_rl_23_t1 = TR_35 ;
	7'h5d :
		RG_rl_23_t1 = TR_35 ;
	7'h5e :
		RG_rl_23_t1 = TR_35 ;
	7'h5f :
		RG_rl_23_t1 = TR_35 ;
	7'h60 :
		RG_rl_23_t1 = TR_35 ;
	7'h61 :
		RG_rl_23_t1 = TR_35 ;
	7'h62 :
		RG_rl_23_t1 = TR_35 ;
	7'h63 :
		RG_rl_23_t1 = TR_35 ;
	7'h64 :
		RG_rl_23_t1 = TR_35 ;
	7'h65 :
		RG_rl_23_t1 = TR_35 ;
	7'h66 :
		RG_rl_23_t1 = TR_35 ;
	7'h67 :
		RG_rl_23_t1 = TR_35 ;
	7'h68 :
		RG_rl_23_t1 = TR_35 ;
	7'h69 :
		RG_rl_23_t1 = TR_35 ;
	7'h6a :
		RG_rl_23_t1 = TR_35 ;
	7'h6b :
		RG_rl_23_t1 = TR_35 ;
	7'h6c :
		RG_rl_23_t1 = TR_35 ;
	7'h6d :
		RG_rl_23_t1 = TR_35 ;
	7'h6e :
		RG_rl_23_t1 = TR_35 ;
	7'h6f :
		RG_rl_23_t1 = TR_35 ;
	7'h70 :
		RG_rl_23_t1 = TR_35 ;
	7'h71 :
		RG_rl_23_t1 = TR_35 ;
	7'h72 :
		RG_rl_23_t1 = TR_35 ;
	7'h73 :
		RG_rl_23_t1 = TR_35 ;
	7'h74 :
		RG_rl_23_t1 = TR_35 ;
	7'h75 :
		RG_rl_23_t1 = TR_35 ;
	7'h76 :
		RG_rl_23_t1 = TR_35 ;
	7'h77 :
		RG_rl_23_t1 = TR_35 ;
	7'h78 :
		RG_rl_23_t1 = TR_35 ;
	7'h79 :
		RG_rl_23_t1 = TR_35 ;
	7'h7a :
		RG_rl_23_t1 = TR_35 ;
	7'h7b :
		RG_rl_23_t1 = TR_35 ;
	7'h7c :
		RG_rl_23_t1 = TR_35 ;
	7'h7d :
		RG_rl_23_t1 = TR_35 ;
	7'h7e :
		RG_rl_23_t1 = TR_35 ;
	7'h7f :
		RG_rl_23_t1 = TR_35 ;
	default :
		RG_rl_23_t1 = 9'hx ;
	endcase
always @ ( RG_rl_23_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_206 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_23_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h17 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_23_t = ( ( { 9{ U_570 } } & RG_rl_206 )
		| ( { 9{ U_569 } } & RG_rl_23_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_23_en = ( U_570 | RG_rl_23_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_23_en )
		RG_rl_23 <= RG_rl_23_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_36 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_24_t1 = TR_36 ;
	7'h01 :
		RG_rl_24_t1 = TR_36 ;
	7'h02 :
		RG_rl_24_t1 = TR_36 ;
	7'h03 :
		RG_rl_24_t1 = TR_36 ;
	7'h04 :
		RG_rl_24_t1 = TR_36 ;
	7'h05 :
		RG_rl_24_t1 = TR_36 ;
	7'h06 :
		RG_rl_24_t1 = TR_36 ;
	7'h07 :
		RG_rl_24_t1 = TR_36 ;
	7'h08 :
		RG_rl_24_t1 = TR_36 ;
	7'h09 :
		RG_rl_24_t1 = TR_36 ;
	7'h0a :
		RG_rl_24_t1 = TR_36 ;
	7'h0b :
		RG_rl_24_t1 = TR_36 ;
	7'h0c :
		RG_rl_24_t1 = TR_36 ;
	7'h0d :
		RG_rl_24_t1 = TR_36 ;
	7'h0e :
		RG_rl_24_t1 = TR_36 ;
	7'h0f :
		RG_rl_24_t1 = TR_36 ;
	7'h10 :
		RG_rl_24_t1 = TR_36 ;
	7'h11 :
		RG_rl_24_t1 = TR_36 ;
	7'h12 :
		RG_rl_24_t1 = TR_36 ;
	7'h13 :
		RG_rl_24_t1 = TR_36 ;
	7'h14 :
		RG_rl_24_t1 = TR_36 ;
	7'h15 :
		RG_rl_24_t1 = TR_36 ;
	7'h16 :
		RG_rl_24_t1 = TR_36 ;
	7'h17 :
		RG_rl_24_t1 = TR_36 ;
	7'h18 :
		RG_rl_24_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h19 :
		RG_rl_24_t1 = TR_36 ;
	7'h1a :
		RG_rl_24_t1 = TR_36 ;
	7'h1b :
		RG_rl_24_t1 = TR_36 ;
	7'h1c :
		RG_rl_24_t1 = TR_36 ;
	7'h1d :
		RG_rl_24_t1 = TR_36 ;
	7'h1e :
		RG_rl_24_t1 = TR_36 ;
	7'h1f :
		RG_rl_24_t1 = TR_36 ;
	7'h20 :
		RG_rl_24_t1 = TR_36 ;
	7'h21 :
		RG_rl_24_t1 = TR_36 ;
	7'h22 :
		RG_rl_24_t1 = TR_36 ;
	7'h23 :
		RG_rl_24_t1 = TR_36 ;
	7'h24 :
		RG_rl_24_t1 = TR_36 ;
	7'h25 :
		RG_rl_24_t1 = TR_36 ;
	7'h26 :
		RG_rl_24_t1 = TR_36 ;
	7'h27 :
		RG_rl_24_t1 = TR_36 ;
	7'h28 :
		RG_rl_24_t1 = TR_36 ;
	7'h29 :
		RG_rl_24_t1 = TR_36 ;
	7'h2a :
		RG_rl_24_t1 = TR_36 ;
	7'h2b :
		RG_rl_24_t1 = TR_36 ;
	7'h2c :
		RG_rl_24_t1 = TR_36 ;
	7'h2d :
		RG_rl_24_t1 = TR_36 ;
	7'h2e :
		RG_rl_24_t1 = TR_36 ;
	7'h2f :
		RG_rl_24_t1 = TR_36 ;
	7'h30 :
		RG_rl_24_t1 = TR_36 ;
	7'h31 :
		RG_rl_24_t1 = TR_36 ;
	7'h32 :
		RG_rl_24_t1 = TR_36 ;
	7'h33 :
		RG_rl_24_t1 = TR_36 ;
	7'h34 :
		RG_rl_24_t1 = TR_36 ;
	7'h35 :
		RG_rl_24_t1 = TR_36 ;
	7'h36 :
		RG_rl_24_t1 = TR_36 ;
	7'h37 :
		RG_rl_24_t1 = TR_36 ;
	7'h38 :
		RG_rl_24_t1 = TR_36 ;
	7'h39 :
		RG_rl_24_t1 = TR_36 ;
	7'h3a :
		RG_rl_24_t1 = TR_36 ;
	7'h3b :
		RG_rl_24_t1 = TR_36 ;
	7'h3c :
		RG_rl_24_t1 = TR_36 ;
	7'h3d :
		RG_rl_24_t1 = TR_36 ;
	7'h3e :
		RG_rl_24_t1 = TR_36 ;
	7'h3f :
		RG_rl_24_t1 = TR_36 ;
	7'h40 :
		RG_rl_24_t1 = TR_36 ;
	7'h41 :
		RG_rl_24_t1 = TR_36 ;
	7'h42 :
		RG_rl_24_t1 = TR_36 ;
	7'h43 :
		RG_rl_24_t1 = TR_36 ;
	7'h44 :
		RG_rl_24_t1 = TR_36 ;
	7'h45 :
		RG_rl_24_t1 = TR_36 ;
	7'h46 :
		RG_rl_24_t1 = TR_36 ;
	7'h47 :
		RG_rl_24_t1 = TR_36 ;
	7'h48 :
		RG_rl_24_t1 = TR_36 ;
	7'h49 :
		RG_rl_24_t1 = TR_36 ;
	7'h4a :
		RG_rl_24_t1 = TR_36 ;
	7'h4b :
		RG_rl_24_t1 = TR_36 ;
	7'h4c :
		RG_rl_24_t1 = TR_36 ;
	7'h4d :
		RG_rl_24_t1 = TR_36 ;
	7'h4e :
		RG_rl_24_t1 = TR_36 ;
	7'h4f :
		RG_rl_24_t1 = TR_36 ;
	7'h50 :
		RG_rl_24_t1 = TR_36 ;
	7'h51 :
		RG_rl_24_t1 = TR_36 ;
	7'h52 :
		RG_rl_24_t1 = TR_36 ;
	7'h53 :
		RG_rl_24_t1 = TR_36 ;
	7'h54 :
		RG_rl_24_t1 = TR_36 ;
	7'h55 :
		RG_rl_24_t1 = TR_36 ;
	7'h56 :
		RG_rl_24_t1 = TR_36 ;
	7'h57 :
		RG_rl_24_t1 = TR_36 ;
	7'h58 :
		RG_rl_24_t1 = TR_36 ;
	7'h59 :
		RG_rl_24_t1 = TR_36 ;
	7'h5a :
		RG_rl_24_t1 = TR_36 ;
	7'h5b :
		RG_rl_24_t1 = TR_36 ;
	7'h5c :
		RG_rl_24_t1 = TR_36 ;
	7'h5d :
		RG_rl_24_t1 = TR_36 ;
	7'h5e :
		RG_rl_24_t1 = TR_36 ;
	7'h5f :
		RG_rl_24_t1 = TR_36 ;
	7'h60 :
		RG_rl_24_t1 = TR_36 ;
	7'h61 :
		RG_rl_24_t1 = TR_36 ;
	7'h62 :
		RG_rl_24_t1 = TR_36 ;
	7'h63 :
		RG_rl_24_t1 = TR_36 ;
	7'h64 :
		RG_rl_24_t1 = TR_36 ;
	7'h65 :
		RG_rl_24_t1 = TR_36 ;
	7'h66 :
		RG_rl_24_t1 = TR_36 ;
	7'h67 :
		RG_rl_24_t1 = TR_36 ;
	7'h68 :
		RG_rl_24_t1 = TR_36 ;
	7'h69 :
		RG_rl_24_t1 = TR_36 ;
	7'h6a :
		RG_rl_24_t1 = TR_36 ;
	7'h6b :
		RG_rl_24_t1 = TR_36 ;
	7'h6c :
		RG_rl_24_t1 = TR_36 ;
	7'h6d :
		RG_rl_24_t1 = TR_36 ;
	7'h6e :
		RG_rl_24_t1 = TR_36 ;
	7'h6f :
		RG_rl_24_t1 = TR_36 ;
	7'h70 :
		RG_rl_24_t1 = TR_36 ;
	7'h71 :
		RG_rl_24_t1 = TR_36 ;
	7'h72 :
		RG_rl_24_t1 = TR_36 ;
	7'h73 :
		RG_rl_24_t1 = TR_36 ;
	7'h74 :
		RG_rl_24_t1 = TR_36 ;
	7'h75 :
		RG_rl_24_t1 = TR_36 ;
	7'h76 :
		RG_rl_24_t1 = TR_36 ;
	7'h77 :
		RG_rl_24_t1 = TR_36 ;
	7'h78 :
		RG_rl_24_t1 = TR_36 ;
	7'h79 :
		RG_rl_24_t1 = TR_36 ;
	7'h7a :
		RG_rl_24_t1 = TR_36 ;
	7'h7b :
		RG_rl_24_t1 = TR_36 ;
	7'h7c :
		RG_rl_24_t1 = TR_36 ;
	7'h7d :
		RG_rl_24_t1 = TR_36 ;
	7'h7e :
		RG_rl_24_t1 = TR_36 ;
	7'h7f :
		RG_rl_24_t1 = TR_36 ;
	default :
		RG_rl_24_t1 = 9'hx ;
	endcase
always @ ( RG_rl_24_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_207 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_24_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h18 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_24_t = ( ( { 9{ U_570 } } & RG_rl_207 )
		| ( { 9{ U_569 } } & RG_rl_24_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_24_en = ( U_570 | RG_rl_24_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_24_en )
		RG_rl_24 <= RG_rl_24_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_37 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_25_t1 = TR_37 ;
	7'h01 :
		RG_rl_25_t1 = TR_37 ;
	7'h02 :
		RG_rl_25_t1 = TR_37 ;
	7'h03 :
		RG_rl_25_t1 = TR_37 ;
	7'h04 :
		RG_rl_25_t1 = TR_37 ;
	7'h05 :
		RG_rl_25_t1 = TR_37 ;
	7'h06 :
		RG_rl_25_t1 = TR_37 ;
	7'h07 :
		RG_rl_25_t1 = TR_37 ;
	7'h08 :
		RG_rl_25_t1 = TR_37 ;
	7'h09 :
		RG_rl_25_t1 = TR_37 ;
	7'h0a :
		RG_rl_25_t1 = TR_37 ;
	7'h0b :
		RG_rl_25_t1 = TR_37 ;
	7'h0c :
		RG_rl_25_t1 = TR_37 ;
	7'h0d :
		RG_rl_25_t1 = TR_37 ;
	7'h0e :
		RG_rl_25_t1 = TR_37 ;
	7'h0f :
		RG_rl_25_t1 = TR_37 ;
	7'h10 :
		RG_rl_25_t1 = TR_37 ;
	7'h11 :
		RG_rl_25_t1 = TR_37 ;
	7'h12 :
		RG_rl_25_t1 = TR_37 ;
	7'h13 :
		RG_rl_25_t1 = TR_37 ;
	7'h14 :
		RG_rl_25_t1 = TR_37 ;
	7'h15 :
		RG_rl_25_t1 = TR_37 ;
	7'h16 :
		RG_rl_25_t1 = TR_37 ;
	7'h17 :
		RG_rl_25_t1 = TR_37 ;
	7'h18 :
		RG_rl_25_t1 = TR_37 ;
	7'h19 :
		RG_rl_25_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1a :
		RG_rl_25_t1 = TR_37 ;
	7'h1b :
		RG_rl_25_t1 = TR_37 ;
	7'h1c :
		RG_rl_25_t1 = TR_37 ;
	7'h1d :
		RG_rl_25_t1 = TR_37 ;
	7'h1e :
		RG_rl_25_t1 = TR_37 ;
	7'h1f :
		RG_rl_25_t1 = TR_37 ;
	7'h20 :
		RG_rl_25_t1 = TR_37 ;
	7'h21 :
		RG_rl_25_t1 = TR_37 ;
	7'h22 :
		RG_rl_25_t1 = TR_37 ;
	7'h23 :
		RG_rl_25_t1 = TR_37 ;
	7'h24 :
		RG_rl_25_t1 = TR_37 ;
	7'h25 :
		RG_rl_25_t1 = TR_37 ;
	7'h26 :
		RG_rl_25_t1 = TR_37 ;
	7'h27 :
		RG_rl_25_t1 = TR_37 ;
	7'h28 :
		RG_rl_25_t1 = TR_37 ;
	7'h29 :
		RG_rl_25_t1 = TR_37 ;
	7'h2a :
		RG_rl_25_t1 = TR_37 ;
	7'h2b :
		RG_rl_25_t1 = TR_37 ;
	7'h2c :
		RG_rl_25_t1 = TR_37 ;
	7'h2d :
		RG_rl_25_t1 = TR_37 ;
	7'h2e :
		RG_rl_25_t1 = TR_37 ;
	7'h2f :
		RG_rl_25_t1 = TR_37 ;
	7'h30 :
		RG_rl_25_t1 = TR_37 ;
	7'h31 :
		RG_rl_25_t1 = TR_37 ;
	7'h32 :
		RG_rl_25_t1 = TR_37 ;
	7'h33 :
		RG_rl_25_t1 = TR_37 ;
	7'h34 :
		RG_rl_25_t1 = TR_37 ;
	7'h35 :
		RG_rl_25_t1 = TR_37 ;
	7'h36 :
		RG_rl_25_t1 = TR_37 ;
	7'h37 :
		RG_rl_25_t1 = TR_37 ;
	7'h38 :
		RG_rl_25_t1 = TR_37 ;
	7'h39 :
		RG_rl_25_t1 = TR_37 ;
	7'h3a :
		RG_rl_25_t1 = TR_37 ;
	7'h3b :
		RG_rl_25_t1 = TR_37 ;
	7'h3c :
		RG_rl_25_t1 = TR_37 ;
	7'h3d :
		RG_rl_25_t1 = TR_37 ;
	7'h3e :
		RG_rl_25_t1 = TR_37 ;
	7'h3f :
		RG_rl_25_t1 = TR_37 ;
	7'h40 :
		RG_rl_25_t1 = TR_37 ;
	7'h41 :
		RG_rl_25_t1 = TR_37 ;
	7'h42 :
		RG_rl_25_t1 = TR_37 ;
	7'h43 :
		RG_rl_25_t1 = TR_37 ;
	7'h44 :
		RG_rl_25_t1 = TR_37 ;
	7'h45 :
		RG_rl_25_t1 = TR_37 ;
	7'h46 :
		RG_rl_25_t1 = TR_37 ;
	7'h47 :
		RG_rl_25_t1 = TR_37 ;
	7'h48 :
		RG_rl_25_t1 = TR_37 ;
	7'h49 :
		RG_rl_25_t1 = TR_37 ;
	7'h4a :
		RG_rl_25_t1 = TR_37 ;
	7'h4b :
		RG_rl_25_t1 = TR_37 ;
	7'h4c :
		RG_rl_25_t1 = TR_37 ;
	7'h4d :
		RG_rl_25_t1 = TR_37 ;
	7'h4e :
		RG_rl_25_t1 = TR_37 ;
	7'h4f :
		RG_rl_25_t1 = TR_37 ;
	7'h50 :
		RG_rl_25_t1 = TR_37 ;
	7'h51 :
		RG_rl_25_t1 = TR_37 ;
	7'h52 :
		RG_rl_25_t1 = TR_37 ;
	7'h53 :
		RG_rl_25_t1 = TR_37 ;
	7'h54 :
		RG_rl_25_t1 = TR_37 ;
	7'h55 :
		RG_rl_25_t1 = TR_37 ;
	7'h56 :
		RG_rl_25_t1 = TR_37 ;
	7'h57 :
		RG_rl_25_t1 = TR_37 ;
	7'h58 :
		RG_rl_25_t1 = TR_37 ;
	7'h59 :
		RG_rl_25_t1 = TR_37 ;
	7'h5a :
		RG_rl_25_t1 = TR_37 ;
	7'h5b :
		RG_rl_25_t1 = TR_37 ;
	7'h5c :
		RG_rl_25_t1 = TR_37 ;
	7'h5d :
		RG_rl_25_t1 = TR_37 ;
	7'h5e :
		RG_rl_25_t1 = TR_37 ;
	7'h5f :
		RG_rl_25_t1 = TR_37 ;
	7'h60 :
		RG_rl_25_t1 = TR_37 ;
	7'h61 :
		RG_rl_25_t1 = TR_37 ;
	7'h62 :
		RG_rl_25_t1 = TR_37 ;
	7'h63 :
		RG_rl_25_t1 = TR_37 ;
	7'h64 :
		RG_rl_25_t1 = TR_37 ;
	7'h65 :
		RG_rl_25_t1 = TR_37 ;
	7'h66 :
		RG_rl_25_t1 = TR_37 ;
	7'h67 :
		RG_rl_25_t1 = TR_37 ;
	7'h68 :
		RG_rl_25_t1 = TR_37 ;
	7'h69 :
		RG_rl_25_t1 = TR_37 ;
	7'h6a :
		RG_rl_25_t1 = TR_37 ;
	7'h6b :
		RG_rl_25_t1 = TR_37 ;
	7'h6c :
		RG_rl_25_t1 = TR_37 ;
	7'h6d :
		RG_rl_25_t1 = TR_37 ;
	7'h6e :
		RG_rl_25_t1 = TR_37 ;
	7'h6f :
		RG_rl_25_t1 = TR_37 ;
	7'h70 :
		RG_rl_25_t1 = TR_37 ;
	7'h71 :
		RG_rl_25_t1 = TR_37 ;
	7'h72 :
		RG_rl_25_t1 = TR_37 ;
	7'h73 :
		RG_rl_25_t1 = TR_37 ;
	7'h74 :
		RG_rl_25_t1 = TR_37 ;
	7'h75 :
		RG_rl_25_t1 = TR_37 ;
	7'h76 :
		RG_rl_25_t1 = TR_37 ;
	7'h77 :
		RG_rl_25_t1 = TR_37 ;
	7'h78 :
		RG_rl_25_t1 = TR_37 ;
	7'h79 :
		RG_rl_25_t1 = TR_37 ;
	7'h7a :
		RG_rl_25_t1 = TR_37 ;
	7'h7b :
		RG_rl_25_t1 = TR_37 ;
	7'h7c :
		RG_rl_25_t1 = TR_37 ;
	7'h7d :
		RG_rl_25_t1 = TR_37 ;
	7'h7e :
		RG_rl_25_t1 = TR_37 ;
	7'h7f :
		RG_rl_25_t1 = TR_37 ;
	default :
		RG_rl_25_t1 = 9'hx ;
	endcase
always @ ( RG_rl_25_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_208 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_25_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h19 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_25_t = ( ( { 9{ U_570 } } & RG_rl_208 )
		| ( { 9{ U_569 } } & RG_rl_25_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_25_en = ( U_570 | RG_rl_25_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_25_en )
		RG_rl_25 <= RG_rl_25_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_38 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_26_t1 = TR_38 ;
	7'h01 :
		RG_rl_26_t1 = TR_38 ;
	7'h02 :
		RG_rl_26_t1 = TR_38 ;
	7'h03 :
		RG_rl_26_t1 = TR_38 ;
	7'h04 :
		RG_rl_26_t1 = TR_38 ;
	7'h05 :
		RG_rl_26_t1 = TR_38 ;
	7'h06 :
		RG_rl_26_t1 = TR_38 ;
	7'h07 :
		RG_rl_26_t1 = TR_38 ;
	7'h08 :
		RG_rl_26_t1 = TR_38 ;
	7'h09 :
		RG_rl_26_t1 = TR_38 ;
	7'h0a :
		RG_rl_26_t1 = TR_38 ;
	7'h0b :
		RG_rl_26_t1 = TR_38 ;
	7'h0c :
		RG_rl_26_t1 = TR_38 ;
	7'h0d :
		RG_rl_26_t1 = TR_38 ;
	7'h0e :
		RG_rl_26_t1 = TR_38 ;
	7'h0f :
		RG_rl_26_t1 = TR_38 ;
	7'h10 :
		RG_rl_26_t1 = TR_38 ;
	7'h11 :
		RG_rl_26_t1 = TR_38 ;
	7'h12 :
		RG_rl_26_t1 = TR_38 ;
	7'h13 :
		RG_rl_26_t1 = TR_38 ;
	7'h14 :
		RG_rl_26_t1 = TR_38 ;
	7'h15 :
		RG_rl_26_t1 = TR_38 ;
	7'h16 :
		RG_rl_26_t1 = TR_38 ;
	7'h17 :
		RG_rl_26_t1 = TR_38 ;
	7'h18 :
		RG_rl_26_t1 = TR_38 ;
	7'h19 :
		RG_rl_26_t1 = TR_38 ;
	7'h1a :
		RG_rl_26_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1b :
		RG_rl_26_t1 = TR_38 ;
	7'h1c :
		RG_rl_26_t1 = TR_38 ;
	7'h1d :
		RG_rl_26_t1 = TR_38 ;
	7'h1e :
		RG_rl_26_t1 = TR_38 ;
	7'h1f :
		RG_rl_26_t1 = TR_38 ;
	7'h20 :
		RG_rl_26_t1 = TR_38 ;
	7'h21 :
		RG_rl_26_t1 = TR_38 ;
	7'h22 :
		RG_rl_26_t1 = TR_38 ;
	7'h23 :
		RG_rl_26_t1 = TR_38 ;
	7'h24 :
		RG_rl_26_t1 = TR_38 ;
	7'h25 :
		RG_rl_26_t1 = TR_38 ;
	7'h26 :
		RG_rl_26_t1 = TR_38 ;
	7'h27 :
		RG_rl_26_t1 = TR_38 ;
	7'h28 :
		RG_rl_26_t1 = TR_38 ;
	7'h29 :
		RG_rl_26_t1 = TR_38 ;
	7'h2a :
		RG_rl_26_t1 = TR_38 ;
	7'h2b :
		RG_rl_26_t1 = TR_38 ;
	7'h2c :
		RG_rl_26_t1 = TR_38 ;
	7'h2d :
		RG_rl_26_t1 = TR_38 ;
	7'h2e :
		RG_rl_26_t1 = TR_38 ;
	7'h2f :
		RG_rl_26_t1 = TR_38 ;
	7'h30 :
		RG_rl_26_t1 = TR_38 ;
	7'h31 :
		RG_rl_26_t1 = TR_38 ;
	7'h32 :
		RG_rl_26_t1 = TR_38 ;
	7'h33 :
		RG_rl_26_t1 = TR_38 ;
	7'h34 :
		RG_rl_26_t1 = TR_38 ;
	7'h35 :
		RG_rl_26_t1 = TR_38 ;
	7'h36 :
		RG_rl_26_t1 = TR_38 ;
	7'h37 :
		RG_rl_26_t1 = TR_38 ;
	7'h38 :
		RG_rl_26_t1 = TR_38 ;
	7'h39 :
		RG_rl_26_t1 = TR_38 ;
	7'h3a :
		RG_rl_26_t1 = TR_38 ;
	7'h3b :
		RG_rl_26_t1 = TR_38 ;
	7'h3c :
		RG_rl_26_t1 = TR_38 ;
	7'h3d :
		RG_rl_26_t1 = TR_38 ;
	7'h3e :
		RG_rl_26_t1 = TR_38 ;
	7'h3f :
		RG_rl_26_t1 = TR_38 ;
	7'h40 :
		RG_rl_26_t1 = TR_38 ;
	7'h41 :
		RG_rl_26_t1 = TR_38 ;
	7'h42 :
		RG_rl_26_t1 = TR_38 ;
	7'h43 :
		RG_rl_26_t1 = TR_38 ;
	7'h44 :
		RG_rl_26_t1 = TR_38 ;
	7'h45 :
		RG_rl_26_t1 = TR_38 ;
	7'h46 :
		RG_rl_26_t1 = TR_38 ;
	7'h47 :
		RG_rl_26_t1 = TR_38 ;
	7'h48 :
		RG_rl_26_t1 = TR_38 ;
	7'h49 :
		RG_rl_26_t1 = TR_38 ;
	7'h4a :
		RG_rl_26_t1 = TR_38 ;
	7'h4b :
		RG_rl_26_t1 = TR_38 ;
	7'h4c :
		RG_rl_26_t1 = TR_38 ;
	7'h4d :
		RG_rl_26_t1 = TR_38 ;
	7'h4e :
		RG_rl_26_t1 = TR_38 ;
	7'h4f :
		RG_rl_26_t1 = TR_38 ;
	7'h50 :
		RG_rl_26_t1 = TR_38 ;
	7'h51 :
		RG_rl_26_t1 = TR_38 ;
	7'h52 :
		RG_rl_26_t1 = TR_38 ;
	7'h53 :
		RG_rl_26_t1 = TR_38 ;
	7'h54 :
		RG_rl_26_t1 = TR_38 ;
	7'h55 :
		RG_rl_26_t1 = TR_38 ;
	7'h56 :
		RG_rl_26_t1 = TR_38 ;
	7'h57 :
		RG_rl_26_t1 = TR_38 ;
	7'h58 :
		RG_rl_26_t1 = TR_38 ;
	7'h59 :
		RG_rl_26_t1 = TR_38 ;
	7'h5a :
		RG_rl_26_t1 = TR_38 ;
	7'h5b :
		RG_rl_26_t1 = TR_38 ;
	7'h5c :
		RG_rl_26_t1 = TR_38 ;
	7'h5d :
		RG_rl_26_t1 = TR_38 ;
	7'h5e :
		RG_rl_26_t1 = TR_38 ;
	7'h5f :
		RG_rl_26_t1 = TR_38 ;
	7'h60 :
		RG_rl_26_t1 = TR_38 ;
	7'h61 :
		RG_rl_26_t1 = TR_38 ;
	7'h62 :
		RG_rl_26_t1 = TR_38 ;
	7'h63 :
		RG_rl_26_t1 = TR_38 ;
	7'h64 :
		RG_rl_26_t1 = TR_38 ;
	7'h65 :
		RG_rl_26_t1 = TR_38 ;
	7'h66 :
		RG_rl_26_t1 = TR_38 ;
	7'h67 :
		RG_rl_26_t1 = TR_38 ;
	7'h68 :
		RG_rl_26_t1 = TR_38 ;
	7'h69 :
		RG_rl_26_t1 = TR_38 ;
	7'h6a :
		RG_rl_26_t1 = TR_38 ;
	7'h6b :
		RG_rl_26_t1 = TR_38 ;
	7'h6c :
		RG_rl_26_t1 = TR_38 ;
	7'h6d :
		RG_rl_26_t1 = TR_38 ;
	7'h6e :
		RG_rl_26_t1 = TR_38 ;
	7'h6f :
		RG_rl_26_t1 = TR_38 ;
	7'h70 :
		RG_rl_26_t1 = TR_38 ;
	7'h71 :
		RG_rl_26_t1 = TR_38 ;
	7'h72 :
		RG_rl_26_t1 = TR_38 ;
	7'h73 :
		RG_rl_26_t1 = TR_38 ;
	7'h74 :
		RG_rl_26_t1 = TR_38 ;
	7'h75 :
		RG_rl_26_t1 = TR_38 ;
	7'h76 :
		RG_rl_26_t1 = TR_38 ;
	7'h77 :
		RG_rl_26_t1 = TR_38 ;
	7'h78 :
		RG_rl_26_t1 = TR_38 ;
	7'h79 :
		RG_rl_26_t1 = TR_38 ;
	7'h7a :
		RG_rl_26_t1 = TR_38 ;
	7'h7b :
		RG_rl_26_t1 = TR_38 ;
	7'h7c :
		RG_rl_26_t1 = TR_38 ;
	7'h7d :
		RG_rl_26_t1 = TR_38 ;
	7'h7e :
		RG_rl_26_t1 = TR_38 ;
	7'h7f :
		RG_rl_26_t1 = TR_38 ;
	default :
		RG_rl_26_t1 = 9'hx ;
	endcase
always @ ( RG_rl_26_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_209 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_26_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h1a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_26_t = ( ( { 9{ U_570 } } & RG_rl_209 )
		| ( { 9{ U_569 } } & RG_rl_26_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_26_en = ( U_570 | RG_rl_26_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_26_en )
		RG_rl_26 <= RG_rl_26_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_39 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_27_t1 = TR_39 ;
	7'h01 :
		RG_rl_27_t1 = TR_39 ;
	7'h02 :
		RG_rl_27_t1 = TR_39 ;
	7'h03 :
		RG_rl_27_t1 = TR_39 ;
	7'h04 :
		RG_rl_27_t1 = TR_39 ;
	7'h05 :
		RG_rl_27_t1 = TR_39 ;
	7'h06 :
		RG_rl_27_t1 = TR_39 ;
	7'h07 :
		RG_rl_27_t1 = TR_39 ;
	7'h08 :
		RG_rl_27_t1 = TR_39 ;
	7'h09 :
		RG_rl_27_t1 = TR_39 ;
	7'h0a :
		RG_rl_27_t1 = TR_39 ;
	7'h0b :
		RG_rl_27_t1 = TR_39 ;
	7'h0c :
		RG_rl_27_t1 = TR_39 ;
	7'h0d :
		RG_rl_27_t1 = TR_39 ;
	7'h0e :
		RG_rl_27_t1 = TR_39 ;
	7'h0f :
		RG_rl_27_t1 = TR_39 ;
	7'h10 :
		RG_rl_27_t1 = TR_39 ;
	7'h11 :
		RG_rl_27_t1 = TR_39 ;
	7'h12 :
		RG_rl_27_t1 = TR_39 ;
	7'h13 :
		RG_rl_27_t1 = TR_39 ;
	7'h14 :
		RG_rl_27_t1 = TR_39 ;
	7'h15 :
		RG_rl_27_t1 = TR_39 ;
	7'h16 :
		RG_rl_27_t1 = TR_39 ;
	7'h17 :
		RG_rl_27_t1 = TR_39 ;
	7'h18 :
		RG_rl_27_t1 = TR_39 ;
	7'h19 :
		RG_rl_27_t1 = TR_39 ;
	7'h1a :
		RG_rl_27_t1 = TR_39 ;
	7'h1b :
		RG_rl_27_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1c :
		RG_rl_27_t1 = TR_39 ;
	7'h1d :
		RG_rl_27_t1 = TR_39 ;
	7'h1e :
		RG_rl_27_t1 = TR_39 ;
	7'h1f :
		RG_rl_27_t1 = TR_39 ;
	7'h20 :
		RG_rl_27_t1 = TR_39 ;
	7'h21 :
		RG_rl_27_t1 = TR_39 ;
	7'h22 :
		RG_rl_27_t1 = TR_39 ;
	7'h23 :
		RG_rl_27_t1 = TR_39 ;
	7'h24 :
		RG_rl_27_t1 = TR_39 ;
	7'h25 :
		RG_rl_27_t1 = TR_39 ;
	7'h26 :
		RG_rl_27_t1 = TR_39 ;
	7'h27 :
		RG_rl_27_t1 = TR_39 ;
	7'h28 :
		RG_rl_27_t1 = TR_39 ;
	7'h29 :
		RG_rl_27_t1 = TR_39 ;
	7'h2a :
		RG_rl_27_t1 = TR_39 ;
	7'h2b :
		RG_rl_27_t1 = TR_39 ;
	7'h2c :
		RG_rl_27_t1 = TR_39 ;
	7'h2d :
		RG_rl_27_t1 = TR_39 ;
	7'h2e :
		RG_rl_27_t1 = TR_39 ;
	7'h2f :
		RG_rl_27_t1 = TR_39 ;
	7'h30 :
		RG_rl_27_t1 = TR_39 ;
	7'h31 :
		RG_rl_27_t1 = TR_39 ;
	7'h32 :
		RG_rl_27_t1 = TR_39 ;
	7'h33 :
		RG_rl_27_t1 = TR_39 ;
	7'h34 :
		RG_rl_27_t1 = TR_39 ;
	7'h35 :
		RG_rl_27_t1 = TR_39 ;
	7'h36 :
		RG_rl_27_t1 = TR_39 ;
	7'h37 :
		RG_rl_27_t1 = TR_39 ;
	7'h38 :
		RG_rl_27_t1 = TR_39 ;
	7'h39 :
		RG_rl_27_t1 = TR_39 ;
	7'h3a :
		RG_rl_27_t1 = TR_39 ;
	7'h3b :
		RG_rl_27_t1 = TR_39 ;
	7'h3c :
		RG_rl_27_t1 = TR_39 ;
	7'h3d :
		RG_rl_27_t1 = TR_39 ;
	7'h3e :
		RG_rl_27_t1 = TR_39 ;
	7'h3f :
		RG_rl_27_t1 = TR_39 ;
	7'h40 :
		RG_rl_27_t1 = TR_39 ;
	7'h41 :
		RG_rl_27_t1 = TR_39 ;
	7'h42 :
		RG_rl_27_t1 = TR_39 ;
	7'h43 :
		RG_rl_27_t1 = TR_39 ;
	7'h44 :
		RG_rl_27_t1 = TR_39 ;
	7'h45 :
		RG_rl_27_t1 = TR_39 ;
	7'h46 :
		RG_rl_27_t1 = TR_39 ;
	7'h47 :
		RG_rl_27_t1 = TR_39 ;
	7'h48 :
		RG_rl_27_t1 = TR_39 ;
	7'h49 :
		RG_rl_27_t1 = TR_39 ;
	7'h4a :
		RG_rl_27_t1 = TR_39 ;
	7'h4b :
		RG_rl_27_t1 = TR_39 ;
	7'h4c :
		RG_rl_27_t1 = TR_39 ;
	7'h4d :
		RG_rl_27_t1 = TR_39 ;
	7'h4e :
		RG_rl_27_t1 = TR_39 ;
	7'h4f :
		RG_rl_27_t1 = TR_39 ;
	7'h50 :
		RG_rl_27_t1 = TR_39 ;
	7'h51 :
		RG_rl_27_t1 = TR_39 ;
	7'h52 :
		RG_rl_27_t1 = TR_39 ;
	7'h53 :
		RG_rl_27_t1 = TR_39 ;
	7'h54 :
		RG_rl_27_t1 = TR_39 ;
	7'h55 :
		RG_rl_27_t1 = TR_39 ;
	7'h56 :
		RG_rl_27_t1 = TR_39 ;
	7'h57 :
		RG_rl_27_t1 = TR_39 ;
	7'h58 :
		RG_rl_27_t1 = TR_39 ;
	7'h59 :
		RG_rl_27_t1 = TR_39 ;
	7'h5a :
		RG_rl_27_t1 = TR_39 ;
	7'h5b :
		RG_rl_27_t1 = TR_39 ;
	7'h5c :
		RG_rl_27_t1 = TR_39 ;
	7'h5d :
		RG_rl_27_t1 = TR_39 ;
	7'h5e :
		RG_rl_27_t1 = TR_39 ;
	7'h5f :
		RG_rl_27_t1 = TR_39 ;
	7'h60 :
		RG_rl_27_t1 = TR_39 ;
	7'h61 :
		RG_rl_27_t1 = TR_39 ;
	7'h62 :
		RG_rl_27_t1 = TR_39 ;
	7'h63 :
		RG_rl_27_t1 = TR_39 ;
	7'h64 :
		RG_rl_27_t1 = TR_39 ;
	7'h65 :
		RG_rl_27_t1 = TR_39 ;
	7'h66 :
		RG_rl_27_t1 = TR_39 ;
	7'h67 :
		RG_rl_27_t1 = TR_39 ;
	7'h68 :
		RG_rl_27_t1 = TR_39 ;
	7'h69 :
		RG_rl_27_t1 = TR_39 ;
	7'h6a :
		RG_rl_27_t1 = TR_39 ;
	7'h6b :
		RG_rl_27_t1 = TR_39 ;
	7'h6c :
		RG_rl_27_t1 = TR_39 ;
	7'h6d :
		RG_rl_27_t1 = TR_39 ;
	7'h6e :
		RG_rl_27_t1 = TR_39 ;
	7'h6f :
		RG_rl_27_t1 = TR_39 ;
	7'h70 :
		RG_rl_27_t1 = TR_39 ;
	7'h71 :
		RG_rl_27_t1 = TR_39 ;
	7'h72 :
		RG_rl_27_t1 = TR_39 ;
	7'h73 :
		RG_rl_27_t1 = TR_39 ;
	7'h74 :
		RG_rl_27_t1 = TR_39 ;
	7'h75 :
		RG_rl_27_t1 = TR_39 ;
	7'h76 :
		RG_rl_27_t1 = TR_39 ;
	7'h77 :
		RG_rl_27_t1 = TR_39 ;
	7'h78 :
		RG_rl_27_t1 = TR_39 ;
	7'h79 :
		RG_rl_27_t1 = TR_39 ;
	7'h7a :
		RG_rl_27_t1 = TR_39 ;
	7'h7b :
		RG_rl_27_t1 = TR_39 ;
	7'h7c :
		RG_rl_27_t1 = TR_39 ;
	7'h7d :
		RG_rl_27_t1 = TR_39 ;
	7'h7e :
		RG_rl_27_t1 = TR_39 ;
	7'h7f :
		RG_rl_27_t1 = TR_39 ;
	default :
		RG_rl_27_t1 = 9'hx ;
	endcase
always @ ( RG_rl_27_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_210 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_27_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h1b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_27_t = ( ( { 9{ U_570 } } & RG_rl_210 )
		| ( { 9{ U_569 } } & RG_rl_27_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_27_en = ( U_570 | RG_rl_27_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_27_en )
		RG_rl_27 <= RG_rl_27_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_40 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_28_t1 = TR_40 ;
	7'h01 :
		RG_rl_28_t1 = TR_40 ;
	7'h02 :
		RG_rl_28_t1 = TR_40 ;
	7'h03 :
		RG_rl_28_t1 = TR_40 ;
	7'h04 :
		RG_rl_28_t1 = TR_40 ;
	7'h05 :
		RG_rl_28_t1 = TR_40 ;
	7'h06 :
		RG_rl_28_t1 = TR_40 ;
	7'h07 :
		RG_rl_28_t1 = TR_40 ;
	7'h08 :
		RG_rl_28_t1 = TR_40 ;
	7'h09 :
		RG_rl_28_t1 = TR_40 ;
	7'h0a :
		RG_rl_28_t1 = TR_40 ;
	7'h0b :
		RG_rl_28_t1 = TR_40 ;
	7'h0c :
		RG_rl_28_t1 = TR_40 ;
	7'h0d :
		RG_rl_28_t1 = TR_40 ;
	7'h0e :
		RG_rl_28_t1 = TR_40 ;
	7'h0f :
		RG_rl_28_t1 = TR_40 ;
	7'h10 :
		RG_rl_28_t1 = TR_40 ;
	7'h11 :
		RG_rl_28_t1 = TR_40 ;
	7'h12 :
		RG_rl_28_t1 = TR_40 ;
	7'h13 :
		RG_rl_28_t1 = TR_40 ;
	7'h14 :
		RG_rl_28_t1 = TR_40 ;
	7'h15 :
		RG_rl_28_t1 = TR_40 ;
	7'h16 :
		RG_rl_28_t1 = TR_40 ;
	7'h17 :
		RG_rl_28_t1 = TR_40 ;
	7'h18 :
		RG_rl_28_t1 = TR_40 ;
	7'h19 :
		RG_rl_28_t1 = TR_40 ;
	7'h1a :
		RG_rl_28_t1 = TR_40 ;
	7'h1b :
		RG_rl_28_t1 = TR_40 ;
	7'h1c :
		RG_rl_28_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1d :
		RG_rl_28_t1 = TR_40 ;
	7'h1e :
		RG_rl_28_t1 = TR_40 ;
	7'h1f :
		RG_rl_28_t1 = TR_40 ;
	7'h20 :
		RG_rl_28_t1 = TR_40 ;
	7'h21 :
		RG_rl_28_t1 = TR_40 ;
	7'h22 :
		RG_rl_28_t1 = TR_40 ;
	7'h23 :
		RG_rl_28_t1 = TR_40 ;
	7'h24 :
		RG_rl_28_t1 = TR_40 ;
	7'h25 :
		RG_rl_28_t1 = TR_40 ;
	7'h26 :
		RG_rl_28_t1 = TR_40 ;
	7'h27 :
		RG_rl_28_t1 = TR_40 ;
	7'h28 :
		RG_rl_28_t1 = TR_40 ;
	7'h29 :
		RG_rl_28_t1 = TR_40 ;
	7'h2a :
		RG_rl_28_t1 = TR_40 ;
	7'h2b :
		RG_rl_28_t1 = TR_40 ;
	7'h2c :
		RG_rl_28_t1 = TR_40 ;
	7'h2d :
		RG_rl_28_t1 = TR_40 ;
	7'h2e :
		RG_rl_28_t1 = TR_40 ;
	7'h2f :
		RG_rl_28_t1 = TR_40 ;
	7'h30 :
		RG_rl_28_t1 = TR_40 ;
	7'h31 :
		RG_rl_28_t1 = TR_40 ;
	7'h32 :
		RG_rl_28_t1 = TR_40 ;
	7'h33 :
		RG_rl_28_t1 = TR_40 ;
	7'h34 :
		RG_rl_28_t1 = TR_40 ;
	7'h35 :
		RG_rl_28_t1 = TR_40 ;
	7'h36 :
		RG_rl_28_t1 = TR_40 ;
	7'h37 :
		RG_rl_28_t1 = TR_40 ;
	7'h38 :
		RG_rl_28_t1 = TR_40 ;
	7'h39 :
		RG_rl_28_t1 = TR_40 ;
	7'h3a :
		RG_rl_28_t1 = TR_40 ;
	7'h3b :
		RG_rl_28_t1 = TR_40 ;
	7'h3c :
		RG_rl_28_t1 = TR_40 ;
	7'h3d :
		RG_rl_28_t1 = TR_40 ;
	7'h3e :
		RG_rl_28_t1 = TR_40 ;
	7'h3f :
		RG_rl_28_t1 = TR_40 ;
	7'h40 :
		RG_rl_28_t1 = TR_40 ;
	7'h41 :
		RG_rl_28_t1 = TR_40 ;
	7'h42 :
		RG_rl_28_t1 = TR_40 ;
	7'h43 :
		RG_rl_28_t1 = TR_40 ;
	7'h44 :
		RG_rl_28_t1 = TR_40 ;
	7'h45 :
		RG_rl_28_t1 = TR_40 ;
	7'h46 :
		RG_rl_28_t1 = TR_40 ;
	7'h47 :
		RG_rl_28_t1 = TR_40 ;
	7'h48 :
		RG_rl_28_t1 = TR_40 ;
	7'h49 :
		RG_rl_28_t1 = TR_40 ;
	7'h4a :
		RG_rl_28_t1 = TR_40 ;
	7'h4b :
		RG_rl_28_t1 = TR_40 ;
	7'h4c :
		RG_rl_28_t1 = TR_40 ;
	7'h4d :
		RG_rl_28_t1 = TR_40 ;
	7'h4e :
		RG_rl_28_t1 = TR_40 ;
	7'h4f :
		RG_rl_28_t1 = TR_40 ;
	7'h50 :
		RG_rl_28_t1 = TR_40 ;
	7'h51 :
		RG_rl_28_t1 = TR_40 ;
	7'h52 :
		RG_rl_28_t1 = TR_40 ;
	7'h53 :
		RG_rl_28_t1 = TR_40 ;
	7'h54 :
		RG_rl_28_t1 = TR_40 ;
	7'h55 :
		RG_rl_28_t1 = TR_40 ;
	7'h56 :
		RG_rl_28_t1 = TR_40 ;
	7'h57 :
		RG_rl_28_t1 = TR_40 ;
	7'h58 :
		RG_rl_28_t1 = TR_40 ;
	7'h59 :
		RG_rl_28_t1 = TR_40 ;
	7'h5a :
		RG_rl_28_t1 = TR_40 ;
	7'h5b :
		RG_rl_28_t1 = TR_40 ;
	7'h5c :
		RG_rl_28_t1 = TR_40 ;
	7'h5d :
		RG_rl_28_t1 = TR_40 ;
	7'h5e :
		RG_rl_28_t1 = TR_40 ;
	7'h5f :
		RG_rl_28_t1 = TR_40 ;
	7'h60 :
		RG_rl_28_t1 = TR_40 ;
	7'h61 :
		RG_rl_28_t1 = TR_40 ;
	7'h62 :
		RG_rl_28_t1 = TR_40 ;
	7'h63 :
		RG_rl_28_t1 = TR_40 ;
	7'h64 :
		RG_rl_28_t1 = TR_40 ;
	7'h65 :
		RG_rl_28_t1 = TR_40 ;
	7'h66 :
		RG_rl_28_t1 = TR_40 ;
	7'h67 :
		RG_rl_28_t1 = TR_40 ;
	7'h68 :
		RG_rl_28_t1 = TR_40 ;
	7'h69 :
		RG_rl_28_t1 = TR_40 ;
	7'h6a :
		RG_rl_28_t1 = TR_40 ;
	7'h6b :
		RG_rl_28_t1 = TR_40 ;
	7'h6c :
		RG_rl_28_t1 = TR_40 ;
	7'h6d :
		RG_rl_28_t1 = TR_40 ;
	7'h6e :
		RG_rl_28_t1 = TR_40 ;
	7'h6f :
		RG_rl_28_t1 = TR_40 ;
	7'h70 :
		RG_rl_28_t1 = TR_40 ;
	7'h71 :
		RG_rl_28_t1 = TR_40 ;
	7'h72 :
		RG_rl_28_t1 = TR_40 ;
	7'h73 :
		RG_rl_28_t1 = TR_40 ;
	7'h74 :
		RG_rl_28_t1 = TR_40 ;
	7'h75 :
		RG_rl_28_t1 = TR_40 ;
	7'h76 :
		RG_rl_28_t1 = TR_40 ;
	7'h77 :
		RG_rl_28_t1 = TR_40 ;
	7'h78 :
		RG_rl_28_t1 = TR_40 ;
	7'h79 :
		RG_rl_28_t1 = TR_40 ;
	7'h7a :
		RG_rl_28_t1 = TR_40 ;
	7'h7b :
		RG_rl_28_t1 = TR_40 ;
	7'h7c :
		RG_rl_28_t1 = TR_40 ;
	7'h7d :
		RG_rl_28_t1 = TR_40 ;
	7'h7e :
		RG_rl_28_t1 = TR_40 ;
	7'h7f :
		RG_rl_28_t1 = TR_40 ;
	default :
		RG_rl_28_t1 = 9'hx ;
	endcase
always @ ( RG_rl_28_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_211 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_28_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h1c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_28_t = ( ( { 9{ U_570 } } & RG_rl_211 )
		| ( { 9{ U_569 } } & RG_rl_28_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_28_en = ( U_570 | RG_rl_28_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_28_en )
		RG_rl_28 <= RG_rl_28_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_41 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_29_t1 = TR_41 ;
	7'h01 :
		RG_rl_29_t1 = TR_41 ;
	7'h02 :
		RG_rl_29_t1 = TR_41 ;
	7'h03 :
		RG_rl_29_t1 = TR_41 ;
	7'h04 :
		RG_rl_29_t1 = TR_41 ;
	7'h05 :
		RG_rl_29_t1 = TR_41 ;
	7'h06 :
		RG_rl_29_t1 = TR_41 ;
	7'h07 :
		RG_rl_29_t1 = TR_41 ;
	7'h08 :
		RG_rl_29_t1 = TR_41 ;
	7'h09 :
		RG_rl_29_t1 = TR_41 ;
	7'h0a :
		RG_rl_29_t1 = TR_41 ;
	7'h0b :
		RG_rl_29_t1 = TR_41 ;
	7'h0c :
		RG_rl_29_t1 = TR_41 ;
	7'h0d :
		RG_rl_29_t1 = TR_41 ;
	7'h0e :
		RG_rl_29_t1 = TR_41 ;
	7'h0f :
		RG_rl_29_t1 = TR_41 ;
	7'h10 :
		RG_rl_29_t1 = TR_41 ;
	7'h11 :
		RG_rl_29_t1 = TR_41 ;
	7'h12 :
		RG_rl_29_t1 = TR_41 ;
	7'h13 :
		RG_rl_29_t1 = TR_41 ;
	7'h14 :
		RG_rl_29_t1 = TR_41 ;
	7'h15 :
		RG_rl_29_t1 = TR_41 ;
	7'h16 :
		RG_rl_29_t1 = TR_41 ;
	7'h17 :
		RG_rl_29_t1 = TR_41 ;
	7'h18 :
		RG_rl_29_t1 = TR_41 ;
	7'h19 :
		RG_rl_29_t1 = TR_41 ;
	7'h1a :
		RG_rl_29_t1 = TR_41 ;
	7'h1b :
		RG_rl_29_t1 = TR_41 ;
	7'h1c :
		RG_rl_29_t1 = TR_41 ;
	7'h1d :
		RG_rl_29_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1e :
		RG_rl_29_t1 = TR_41 ;
	7'h1f :
		RG_rl_29_t1 = TR_41 ;
	7'h20 :
		RG_rl_29_t1 = TR_41 ;
	7'h21 :
		RG_rl_29_t1 = TR_41 ;
	7'h22 :
		RG_rl_29_t1 = TR_41 ;
	7'h23 :
		RG_rl_29_t1 = TR_41 ;
	7'h24 :
		RG_rl_29_t1 = TR_41 ;
	7'h25 :
		RG_rl_29_t1 = TR_41 ;
	7'h26 :
		RG_rl_29_t1 = TR_41 ;
	7'h27 :
		RG_rl_29_t1 = TR_41 ;
	7'h28 :
		RG_rl_29_t1 = TR_41 ;
	7'h29 :
		RG_rl_29_t1 = TR_41 ;
	7'h2a :
		RG_rl_29_t1 = TR_41 ;
	7'h2b :
		RG_rl_29_t1 = TR_41 ;
	7'h2c :
		RG_rl_29_t1 = TR_41 ;
	7'h2d :
		RG_rl_29_t1 = TR_41 ;
	7'h2e :
		RG_rl_29_t1 = TR_41 ;
	7'h2f :
		RG_rl_29_t1 = TR_41 ;
	7'h30 :
		RG_rl_29_t1 = TR_41 ;
	7'h31 :
		RG_rl_29_t1 = TR_41 ;
	7'h32 :
		RG_rl_29_t1 = TR_41 ;
	7'h33 :
		RG_rl_29_t1 = TR_41 ;
	7'h34 :
		RG_rl_29_t1 = TR_41 ;
	7'h35 :
		RG_rl_29_t1 = TR_41 ;
	7'h36 :
		RG_rl_29_t1 = TR_41 ;
	7'h37 :
		RG_rl_29_t1 = TR_41 ;
	7'h38 :
		RG_rl_29_t1 = TR_41 ;
	7'h39 :
		RG_rl_29_t1 = TR_41 ;
	7'h3a :
		RG_rl_29_t1 = TR_41 ;
	7'h3b :
		RG_rl_29_t1 = TR_41 ;
	7'h3c :
		RG_rl_29_t1 = TR_41 ;
	7'h3d :
		RG_rl_29_t1 = TR_41 ;
	7'h3e :
		RG_rl_29_t1 = TR_41 ;
	7'h3f :
		RG_rl_29_t1 = TR_41 ;
	7'h40 :
		RG_rl_29_t1 = TR_41 ;
	7'h41 :
		RG_rl_29_t1 = TR_41 ;
	7'h42 :
		RG_rl_29_t1 = TR_41 ;
	7'h43 :
		RG_rl_29_t1 = TR_41 ;
	7'h44 :
		RG_rl_29_t1 = TR_41 ;
	7'h45 :
		RG_rl_29_t1 = TR_41 ;
	7'h46 :
		RG_rl_29_t1 = TR_41 ;
	7'h47 :
		RG_rl_29_t1 = TR_41 ;
	7'h48 :
		RG_rl_29_t1 = TR_41 ;
	7'h49 :
		RG_rl_29_t1 = TR_41 ;
	7'h4a :
		RG_rl_29_t1 = TR_41 ;
	7'h4b :
		RG_rl_29_t1 = TR_41 ;
	7'h4c :
		RG_rl_29_t1 = TR_41 ;
	7'h4d :
		RG_rl_29_t1 = TR_41 ;
	7'h4e :
		RG_rl_29_t1 = TR_41 ;
	7'h4f :
		RG_rl_29_t1 = TR_41 ;
	7'h50 :
		RG_rl_29_t1 = TR_41 ;
	7'h51 :
		RG_rl_29_t1 = TR_41 ;
	7'h52 :
		RG_rl_29_t1 = TR_41 ;
	7'h53 :
		RG_rl_29_t1 = TR_41 ;
	7'h54 :
		RG_rl_29_t1 = TR_41 ;
	7'h55 :
		RG_rl_29_t1 = TR_41 ;
	7'h56 :
		RG_rl_29_t1 = TR_41 ;
	7'h57 :
		RG_rl_29_t1 = TR_41 ;
	7'h58 :
		RG_rl_29_t1 = TR_41 ;
	7'h59 :
		RG_rl_29_t1 = TR_41 ;
	7'h5a :
		RG_rl_29_t1 = TR_41 ;
	7'h5b :
		RG_rl_29_t1 = TR_41 ;
	7'h5c :
		RG_rl_29_t1 = TR_41 ;
	7'h5d :
		RG_rl_29_t1 = TR_41 ;
	7'h5e :
		RG_rl_29_t1 = TR_41 ;
	7'h5f :
		RG_rl_29_t1 = TR_41 ;
	7'h60 :
		RG_rl_29_t1 = TR_41 ;
	7'h61 :
		RG_rl_29_t1 = TR_41 ;
	7'h62 :
		RG_rl_29_t1 = TR_41 ;
	7'h63 :
		RG_rl_29_t1 = TR_41 ;
	7'h64 :
		RG_rl_29_t1 = TR_41 ;
	7'h65 :
		RG_rl_29_t1 = TR_41 ;
	7'h66 :
		RG_rl_29_t1 = TR_41 ;
	7'h67 :
		RG_rl_29_t1 = TR_41 ;
	7'h68 :
		RG_rl_29_t1 = TR_41 ;
	7'h69 :
		RG_rl_29_t1 = TR_41 ;
	7'h6a :
		RG_rl_29_t1 = TR_41 ;
	7'h6b :
		RG_rl_29_t1 = TR_41 ;
	7'h6c :
		RG_rl_29_t1 = TR_41 ;
	7'h6d :
		RG_rl_29_t1 = TR_41 ;
	7'h6e :
		RG_rl_29_t1 = TR_41 ;
	7'h6f :
		RG_rl_29_t1 = TR_41 ;
	7'h70 :
		RG_rl_29_t1 = TR_41 ;
	7'h71 :
		RG_rl_29_t1 = TR_41 ;
	7'h72 :
		RG_rl_29_t1 = TR_41 ;
	7'h73 :
		RG_rl_29_t1 = TR_41 ;
	7'h74 :
		RG_rl_29_t1 = TR_41 ;
	7'h75 :
		RG_rl_29_t1 = TR_41 ;
	7'h76 :
		RG_rl_29_t1 = TR_41 ;
	7'h77 :
		RG_rl_29_t1 = TR_41 ;
	7'h78 :
		RG_rl_29_t1 = TR_41 ;
	7'h79 :
		RG_rl_29_t1 = TR_41 ;
	7'h7a :
		RG_rl_29_t1 = TR_41 ;
	7'h7b :
		RG_rl_29_t1 = TR_41 ;
	7'h7c :
		RG_rl_29_t1 = TR_41 ;
	7'h7d :
		RG_rl_29_t1 = TR_41 ;
	7'h7e :
		RG_rl_29_t1 = TR_41 ;
	7'h7f :
		RG_rl_29_t1 = TR_41 ;
	default :
		RG_rl_29_t1 = 9'hx ;
	endcase
always @ ( RG_rl_29_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_212 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_29_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h1d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_29_t = ( ( { 9{ U_570 } } & RG_rl_212 )
		| ( { 9{ U_569 } } & RG_rl_29_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_29_en = ( U_570 | RG_rl_29_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_29_en )
		RG_rl_29 <= RG_rl_29_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_42 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_30_t1 = TR_42 ;
	7'h01 :
		RG_rl_30_t1 = TR_42 ;
	7'h02 :
		RG_rl_30_t1 = TR_42 ;
	7'h03 :
		RG_rl_30_t1 = TR_42 ;
	7'h04 :
		RG_rl_30_t1 = TR_42 ;
	7'h05 :
		RG_rl_30_t1 = TR_42 ;
	7'h06 :
		RG_rl_30_t1 = TR_42 ;
	7'h07 :
		RG_rl_30_t1 = TR_42 ;
	7'h08 :
		RG_rl_30_t1 = TR_42 ;
	7'h09 :
		RG_rl_30_t1 = TR_42 ;
	7'h0a :
		RG_rl_30_t1 = TR_42 ;
	7'h0b :
		RG_rl_30_t1 = TR_42 ;
	7'h0c :
		RG_rl_30_t1 = TR_42 ;
	7'h0d :
		RG_rl_30_t1 = TR_42 ;
	7'h0e :
		RG_rl_30_t1 = TR_42 ;
	7'h0f :
		RG_rl_30_t1 = TR_42 ;
	7'h10 :
		RG_rl_30_t1 = TR_42 ;
	7'h11 :
		RG_rl_30_t1 = TR_42 ;
	7'h12 :
		RG_rl_30_t1 = TR_42 ;
	7'h13 :
		RG_rl_30_t1 = TR_42 ;
	7'h14 :
		RG_rl_30_t1 = TR_42 ;
	7'h15 :
		RG_rl_30_t1 = TR_42 ;
	7'h16 :
		RG_rl_30_t1 = TR_42 ;
	7'h17 :
		RG_rl_30_t1 = TR_42 ;
	7'h18 :
		RG_rl_30_t1 = TR_42 ;
	7'h19 :
		RG_rl_30_t1 = TR_42 ;
	7'h1a :
		RG_rl_30_t1 = TR_42 ;
	7'h1b :
		RG_rl_30_t1 = TR_42 ;
	7'h1c :
		RG_rl_30_t1 = TR_42 ;
	7'h1d :
		RG_rl_30_t1 = TR_42 ;
	7'h1e :
		RG_rl_30_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h1f :
		RG_rl_30_t1 = TR_42 ;
	7'h20 :
		RG_rl_30_t1 = TR_42 ;
	7'h21 :
		RG_rl_30_t1 = TR_42 ;
	7'h22 :
		RG_rl_30_t1 = TR_42 ;
	7'h23 :
		RG_rl_30_t1 = TR_42 ;
	7'h24 :
		RG_rl_30_t1 = TR_42 ;
	7'h25 :
		RG_rl_30_t1 = TR_42 ;
	7'h26 :
		RG_rl_30_t1 = TR_42 ;
	7'h27 :
		RG_rl_30_t1 = TR_42 ;
	7'h28 :
		RG_rl_30_t1 = TR_42 ;
	7'h29 :
		RG_rl_30_t1 = TR_42 ;
	7'h2a :
		RG_rl_30_t1 = TR_42 ;
	7'h2b :
		RG_rl_30_t1 = TR_42 ;
	7'h2c :
		RG_rl_30_t1 = TR_42 ;
	7'h2d :
		RG_rl_30_t1 = TR_42 ;
	7'h2e :
		RG_rl_30_t1 = TR_42 ;
	7'h2f :
		RG_rl_30_t1 = TR_42 ;
	7'h30 :
		RG_rl_30_t1 = TR_42 ;
	7'h31 :
		RG_rl_30_t1 = TR_42 ;
	7'h32 :
		RG_rl_30_t1 = TR_42 ;
	7'h33 :
		RG_rl_30_t1 = TR_42 ;
	7'h34 :
		RG_rl_30_t1 = TR_42 ;
	7'h35 :
		RG_rl_30_t1 = TR_42 ;
	7'h36 :
		RG_rl_30_t1 = TR_42 ;
	7'h37 :
		RG_rl_30_t1 = TR_42 ;
	7'h38 :
		RG_rl_30_t1 = TR_42 ;
	7'h39 :
		RG_rl_30_t1 = TR_42 ;
	7'h3a :
		RG_rl_30_t1 = TR_42 ;
	7'h3b :
		RG_rl_30_t1 = TR_42 ;
	7'h3c :
		RG_rl_30_t1 = TR_42 ;
	7'h3d :
		RG_rl_30_t1 = TR_42 ;
	7'h3e :
		RG_rl_30_t1 = TR_42 ;
	7'h3f :
		RG_rl_30_t1 = TR_42 ;
	7'h40 :
		RG_rl_30_t1 = TR_42 ;
	7'h41 :
		RG_rl_30_t1 = TR_42 ;
	7'h42 :
		RG_rl_30_t1 = TR_42 ;
	7'h43 :
		RG_rl_30_t1 = TR_42 ;
	7'h44 :
		RG_rl_30_t1 = TR_42 ;
	7'h45 :
		RG_rl_30_t1 = TR_42 ;
	7'h46 :
		RG_rl_30_t1 = TR_42 ;
	7'h47 :
		RG_rl_30_t1 = TR_42 ;
	7'h48 :
		RG_rl_30_t1 = TR_42 ;
	7'h49 :
		RG_rl_30_t1 = TR_42 ;
	7'h4a :
		RG_rl_30_t1 = TR_42 ;
	7'h4b :
		RG_rl_30_t1 = TR_42 ;
	7'h4c :
		RG_rl_30_t1 = TR_42 ;
	7'h4d :
		RG_rl_30_t1 = TR_42 ;
	7'h4e :
		RG_rl_30_t1 = TR_42 ;
	7'h4f :
		RG_rl_30_t1 = TR_42 ;
	7'h50 :
		RG_rl_30_t1 = TR_42 ;
	7'h51 :
		RG_rl_30_t1 = TR_42 ;
	7'h52 :
		RG_rl_30_t1 = TR_42 ;
	7'h53 :
		RG_rl_30_t1 = TR_42 ;
	7'h54 :
		RG_rl_30_t1 = TR_42 ;
	7'h55 :
		RG_rl_30_t1 = TR_42 ;
	7'h56 :
		RG_rl_30_t1 = TR_42 ;
	7'h57 :
		RG_rl_30_t1 = TR_42 ;
	7'h58 :
		RG_rl_30_t1 = TR_42 ;
	7'h59 :
		RG_rl_30_t1 = TR_42 ;
	7'h5a :
		RG_rl_30_t1 = TR_42 ;
	7'h5b :
		RG_rl_30_t1 = TR_42 ;
	7'h5c :
		RG_rl_30_t1 = TR_42 ;
	7'h5d :
		RG_rl_30_t1 = TR_42 ;
	7'h5e :
		RG_rl_30_t1 = TR_42 ;
	7'h5f :
		RG_rl_30_t1 = TR_42 ;
	7'h60 :
		RG_rl_30_t1 = TR_42 ;
	7'h61 :
		RG_rl_30_t1 = TR_42 ;
	7'h62 :
		RG_rl_30_t1 = TR_42 ;
	7'h63 :
		RG_rl_30_t1 = TR_42 ;
	7'h64 :
		RG_rl_30_t1 = TR_42 ;
	7'h65 :
		RG_rl_30_t1 = TR_42 ;
	7'h66 :
		RG_rl_30_t1 = TR_42 ;
	7'h67 :
		RG_rl_30_t1 = TR_42 ;
	7'h68 :
		RG_rl_30_t1 = TR_42 ;
	7'h69 :
		RG_rl_30_t1 = TR_42 ;
	7'h6a :
		RG_rl_30_t1 = TR_42 ;
	7'h6b :
		RG_rl_30_t1 = TR_42 ;
	7'h6c :
		RG_rl_30_t1 = TR_42 ;
	7'h6d :
		RG_rl_30_t1 = TR_42 ;
	7'h6e :
		RG_rl_30_t1 = TR_42 ;
	7'h6f :
		RG_rl_30_t1 = TR_42 ;
	7'h70 :
		RG_rl_30_t1 = TR_42 ;
	7'h71 :
		RG_rl_30_t1 = TR_42 ;
	7'h72 :
		RG_rl_30_t1 = TR_42 ;
	7'h73 :
		RG_rl_30_t1 = TR_42 ;
	7'h74 :
		RG_rl_30_t1 = TR_42 ;
	7'h75 :
		RG_rl_30_t1 = TR_42 ;
	7'h76 :
		RG_rl_30_t1 = TR_42 ;
	7'h77 :
		RG_rl_30_t1 = TR_42 ;
	7'h78 :
		RG_rl_30_t1 = TR_42 ;
	7'h79 :
		RG_rl_30_t1 = TR_42 ;
	7'h7a :
		RG_rl_30_t1 = TR_42 ;
	7'h7b :
		RG_rl_30_t1 = TR_42 ;
	7'h7c :
		RG_rl_30_t1 = TR_42 ;
	7'h7d :
		RG_rl_30_t1 = TR_42 ;
	7'h7e :
		RG_rl_30_t1 = TR_42 ;
	7'h7f :
		RG_rl_30_t1 = TR_42 ;
	default :
		RG_rl_30_t1 = 9'hx ;
	endcase
always @ ( RG_rl_30_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_213 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_30_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h1e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_30_t = ( ( { 9{ U_570 } } & RG_rl_213 )
		| ( { 9{ U_569 } } & RG_rl_30_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_30_en = ( U_570 | RG_rl_30_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_30_en )
		RG_rl_30 <= RG_rl_30_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_43 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_31_t1 = TR_43 ;
	7'h01 :
		RG_rl_31_t1 = TR_43 ;
	7'h02 :
		RG_rl_31_t1 = TR_43 ;
	7'h03 :
		RG_rl_31_t1 = TR_43 ;
	7'h04 :
		RG_rl_31_t1 = TR_43 ;
	7'h05 :
		RG_rl_31_t1 = TR_43 ;
	7'h06 :
		RG_rl_31_t1 = TR_43 ;
	7'h07 :
		RG_rl_31_t1 = TR_43 ;
	7'h08 :
		RG_rl_31_t1 = TR_43 ;
	7'h09 :
		RG_rl_31_t1 = TR_43 ;
	7'h0a :
		RG_rl_31_t1 = TR_43 ;
	7'h0b :
		RG_rl_31_t1 = TR_43 ;
	7'h0c :
		RG_rl_31_t1 = TR_43 ;
	7'h0d :
		RG_rl_31_t1 = TR_43 ;
	7'h0e :
		RG_rl_31_t1 = TR_43 ;
	7'h0f :
		RG_rl_31_t1 = TR_43 ;
	7'h10 :
		RG_rl_31_t1 = TR_43 ;
	7'h11 :
		RG_rl_31_t1 = TR_43 ;
	7'h12 :
		RG_rl_31_t1 = TR_43 ;
	7'h13 :
		RG_rl_31_t1 = TR_43 ;
	7'h14 :
		RG_rl_31_t1 = TR_43 ;
	7'h15 :
		RG_rl_31_t1 = TR_43 ;
	7'h16 :
		RG_rl_31_t1 = TR_43 ;
	7'h17 :
		RG_rl_31_t1 = TR_43 ;
	7'h18 :
		RG_rl_31_t1 = TR_43 ;
	7'h19 :
		RG_rl_31_t1 = TR_43 ;
	7'h1a :
		RG_rl_31_t1 = TR_43 ;
	7'h1b :
		RG_rl_31_t1 = TR_43 ;
	7'h1c :
		RG_rl_31_t1 = TR_43 ;
	7'h1d :
		RG_rl_31_t1 = TR_43 ;
	7'h1e :
		RG_rl_31_t1 = TR_43 ;
	7'h1f :
		RG_rl_31_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h20 :
		RG_rl_31_t1 = TR_43 ;
	7'h21 :
		RG_rl_31_t1 = TR_43 ;
	7'h22 :
		RG_rl_31_t1 = TR_43 ;
	7'h23 :
		RG_rl_31_t1 = TR_43 ;
	7'h24 :
		RG_rl_31_t1 = TR_43 ;
	7'h25 :
		RG_rl_31_t1 = TR_43 ;
	7'h26 :
		RG_rl_31_t1 = TR_43 ;
	7'h27 :
		RG_rl_31_t1 = TR_43 ;
	7'h28 :
		RG_rl_31_t1 = TR_43 ;
	7'h29 :
		RG_rl_31_t1 = TR_43 ;
	7'h2a :
		RG_rl_31_t1 = TR_43 ;
	7'h2b :
		RG_rl_31_t1 = TR_43 ;
	7'h2c :
		RG_rl_31_t1 = TR_43 ;
	7'h2d :
		RG_rl_31_t1 = TR_43 ;
	7'h2e :
		RG_rl_31_t1 = TR_43 ;
	7'h2f :
		RG_rl_31_t1 = TR_43 ;
	7'h30 :
		RG_rl_31_t1 = TR_43 ;
	7'h31 :
		RG_rl_31_t1 = TR_43 ;
	7'h32 :
		RG_rl_31_t1 = TR_43 ;
	7'h33 :
		RG_rl_31_t1 = TR_43 ;
	7'h34 :
		RG_rl_31_t1 = TR_43 ;
	7'h35 :
		RG_rl_31_t1 = TR_43 ;
	7'h36 :
		RG_rl_31_t1 = TR_43 ;
	7'h37 :
		RG_rl_31_t1 = TR_43 ;
	7'h38 :
		RG_rl_31_t1 = TR_43 ;
	7'h39 :
		RG_rl_31_t1 = TR_43 ;
	7'h3a :
		RG_rl_31_t1 = TR_43 ;
	7'h3b :
		RG_rl_31_t1 = TR_43 ;
	7'h3c :
		RG_rl_31_t1 = TR_43 ;
	7'h3d :
		RG_rl_31_t1 = TR_43 ;
	7'h3e :
		RG_rl_31_t1 = TR_43 ;
	7'h3f :
		RG_rl_31_t1 = TR_43 ;
	7'h40 :
		RG_rl_31_t1 = TR_43 ;
	7'h41 :
		RG_rl_31_t1 = TR_43 ;
	7'h42 :
		RG_rl_31_t1 = TR_43 ;
	7'h43 :
		RG_rl_31_t1 = TR_43 ;
	7'h44 :
		RG_rl_31_t1 = TR_43 ;
	7'h45 :
		RG_rl_31_t1 = TR_43 ;
	7'h46 :
		RG_rl_31_t1 = TR_43 ;
	7'h47 :
		RG_rl_31_t1 = TR_43 ;
	7'h48 :
		RG_rl_31_t1 = TR_43 ;
	7'h49 :
		RG_rl_31_t1 = TR_43 ;
	7'h4a :
		RG_rl_31_t1 = TR_43 ;
	7'h4b :
		RG_rl_31_t1 = TR_43 ;
	7'h4c :
		RG_rl_31_t1 = TR_43 ;
	7'h4d :
		RG_rl_31_t1 = TR_43 ;
	7'h4e :
		RG_rl_31_t1 = TR_43 ;
	7'h4f :
		RG_rl_31_t1 = TR_43 ;
	7'h50 :
		RG_rl_31_t1 = TR_43 ;
	7'h51 :
		RG_rl_31_t1 = TR_43 ;
	7'h52 :
		RG_rl_31_t1 = TR_43 ;
	7'h53 :
		RG_rl_31_t1 = TR_43 ;
	7'h54 :
		RG_rl_31_t1 = TR_43 ;
	7'h55 :
		RG_rl_31_t1 = TR_43 ;
	7'h56 :
		RG_rl_31_t1 = TR_43 ;
	7'h57 :
		RG_rl_31_t1 = TR_43 ;
	7'h58 :
		RG_rl_31_t1 = TR_43 ;
	7'h59 :
		RG_rl_31_t1 = TR_43 ;
	7'h5a :
		RG_rl_31_t1 = TR_43 ;
	7'h5b :
		RG_rl_31_t1 = TR_43 ;
	7'h5c :
		RG_rl_31_t1 = TR_43 ;
	7'h5d :
		RG_rl_31_t1 = TR_43 ;
	7'h5e :
		RG_rl_31_t1 = TR_43 ;
	7'h5f :
		RG_rl_31_t1 = TR_43 ;
	7'h60 :
		RG_rl_31_t1 = TR_43 ;
	7'h61 :
		RG_rl_31_t1 = TR_43 ;
	7'h62 :
		RG_rl_31_t1 = TR_43 ;
	7'h63 :
		RG_rl_31_t1 = TR_43 ;
	7'h64 :
		RG_rl_31_t1 = TR_43 ;
	7'h65 :
		RG_rl_31_t1 = TR_43 ;
	7'h66 :
		RG_rl_31_t1 = TR_43 ;
	7'h67 :
		RG_rl_31_t1 = TR_43 ;
	7'h68 :
		RG_rl_31_t1 = TR_43 ;
	7'h69 :
		RG_rl_31_t1 = TR_43 ;
	7'h6a :
		RG_rl_31_t1 = TR_43 ;
	7'h6b :
		RG_rl_31_t1 = TR_43 ;
	7'h6c :
		RG_rl_31_t1 = TR_43 ;
	7'h6d :
		RG_rl_31_t1 = TR_43 ;
	7'h6e :
		RG_rl_31_t1 = TR_43 ;
	7'h6f :
		RG_rl_31_t1 = TR_43 ;
	7'h70 :
		RG_rl_31_t1 = TR_43 ;
	7'h71 :
		RG_rl_31_t1 = TR_43 ;
	7'h72 :
		RG_rl_31_t1 = TR_43 ;
	7'h73 :
		RG_rl_31_t1 = TR_43 ;
	7'h74 :
		RG_rl_31_t1 = TR_43 ;
	7'h75 :
		RG_rl_31_t1 = TR_43 ;
	7'h76 :
		RG_rl_31_t1 = TR_43 ;
	7'h77 :
		RG_rl_31_t1 = TR_43 ;
	7'h78 :
		RG_rl_31_t1 = TR_43 ;
	7'h79 :
		RG_rl_31_t1 = TR_43 ;
	7'h7a :
		RG_rl_31_t1 = TR_43 ;
	7'h7b :
		RG_rl_31_t1 = TR_43 ;
	7'h7c :
		RG_rl_31_t1 = TR_43 ;
	7'h7d :
		RG_rl_31_t1 = TR_43 ;
	7'h7e :
		RG_rl_31_t1 = TR_43 ;
	7'h7f :
		RG_rl_31_t1 = TR_43 ;
	default :
		RG_rl_31_t1 = 9'hx ;
	endcase
always @ ( RG_rl_31_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_214 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_31_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h1f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_31_t = ( ( { 9{ U_570 } } & RG_rl_214 )
		| ( { 9{ U_569 } } & RG_rl_31_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_31_en = ( U_570 | RG_rl_31_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_31_en )
		RG_rl_31 <= RG_rl_31_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_44 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_32_t1 = TR_44 ;
	7'h01 :
		RG_rl_32_t1 = TR_44 ;
	7'h02 :
		RG_rl_32_t1 = TR_44 ;
	7'h03 :
		RG_rl_32_t1 = TR_44 ;
	7'h04 :
		RG_rl_32_t1 = TR_44 ;
	7'h05 :
		RG_rl_32_t1 = TR_44 ;
	7'h06 :
		RG_rl_32_t1 = TR_44 ;
	7'h07 :
		RG_rl_32_t1 = TR_44 ;
	7'h08 :
		RG_rl_32_t1 = TR_44 ;
	7'h09 :
		RG_rl_32_t1 = TR_44 ;
	7'h0a :
		RG_rl_32_t1 = TR_44 ;
	7'h0b :
		RG_rl_32_t1 = TR_44 ;
	7'h0c :
		RG_rl_32_t1 = TR_44 ;
	7'h0d :
		RG_rl_32_t1 = TR_44 ;
	7'h0e :
		RG_rl_32_t1 = TR_44 ;
	7'h0f :
		RG_rl_32_t1 = TR_44 ;
	7'h10 :
		RG_rl_32_t1 = TR_44 ;
	7'h11 :
		RG_rl_32_t1 = TR_44 ;
	7'h12 :
		RG_rl_32_t1 = TR_44 ;
	7'h13 :
		RG_rl_32_t1 = TR_44 ;
	7'h14 :
		RG_rl_32_t1 = TR_44 ;
	7'h15 :
		RG_rl_32_t1 = TR_44 ;
	7'h16 :
		RG_rl_32_t1 = TR_44 ;
	7'h17 :
		RG_rl_32_t1 = TR_44 ;
	7'h18 :
		RG_rl_32_t1 = TR_44 ;
	7'h19 :
		RG_rl_32_t1 = TR_44 ;
	7'h1a :
		RG_rl_32_t1 = TR_44 ;
	7'h1b :
		RG_rl_32_t1 = TR_44 ;
	7'h1c :
		RG_rl_32_t1 = TR_44 ;
	7'h1d :
		RG_rl_32_t1 = TR_44 ;
	7'h1e :
		RG_rl_32_t1 = TR_44 ;
	7'h1f :
		RG_rl_32_t1 = TR_44 ;
	7'h20 :
		RG_rl_32_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h21 :
		RG_rl_32_t1 = TR_44 ;
	7'h22 :
		RG_rl_32_t1 = TR_44 ;
	7'h23 :
		RG_rl_32_t1 = TR_44 ;
	7'h24 :
		RG_rl_32_t1 = TR_44 ;
	7'h25 :
		RG_rl_32_t1 = TR_44 ;
	7'h26 :
		RG_rl_32_t1 = TR_44 ;
	7'h27 :
		RG_rl_32_t1 = TR_44 ;
	7'h28 :
		RG_rl_32_t1 = TR_44 ;
	7'h29 :
		RG_rl_32_t1 = TR_44 ;
	7'h2a :
		RG_rl_32_t1 = TR_44 ;
	7'h2b :
		RG_rl_32_t1 = TR_44 ;
	7'h2c :
		RG_rl_32_t1 = TR_44 ;
	7'h2d :
		RG_rl_32_t1 = TR_44 ;
	7'h2e :
		RG_rl_32_t1 = TR_44 ;
	7'h2f :
		RG_rl_32_t1 = TR_44 ;
	7'h30 :
		RG_rl_32_t1 = TR_44 ;
	7'h31 :
		RG_rl_32_t1 = TR_44 ;
	7'h32 :
		RG_rl_32_t1 = TR_44 ;
	7'h33 :
		RG_rl_32_t1 = TR_44 ;
	7'h34 :
		RG_rl_32_t1 = TR_44 ;
	7'h35 :
		RG_rl_32_t1 = TR_44 ;
	7'h36 :
		RG_rl_32_t1 = TR_44 ;
	7'h37 :
		RG_rl_32_t1 = TR_44 ;
	7'h38 :
		RG_rl_32_t1 = TR_44 ;
	7'h39 :
		RG_rl_32_t1 = TR_44 ;
	7'h3a :
		RG_rl_32_t1 = TR_44 ;
	7'h3b :
		RG_rl_32_t1 = TR_44 ;
	7'h3c :
		RG_rl_32_t1 = TR_44 ;
	7'h3d :
		RG_rl_32_t1 = TR_44 ;
	7'h3e :
		RG_rl_32_t1 = TR_44 ;
	7'h3f :
		RG_rl_32_t1 = TR_44 ;
	7'h40 :
		RG_rl_32_t1 = TR_44 ;
	7'h41 :
		RG_rl_32_t1 = TR_44 ;
	7'h42 :
		RG_rl_32_t1 = TR_44 ;
	7'h43 :
		RG_rl_32_t1 = TR_44 ;
	7'h44 :
		RG_rl_32_t1 = TR_44 ;
	7'h45 :
		RG_rl_32_t1 = TR_44 ;
	7'h46 :
		RG_rl_32_t1 = TR_44 ;
	7'h47 :
		RG_rl_32_t1 = TR_44 ;
	7'h48 :
		RG_rl_32_t1 = TR_44 ;
	7'h49 :
		RG_rl_32_t1 = TR_44 ;
	7'h4a :
		RG_rl_32_t1 = TR_44 ;
	7'h4b :
		RG_rl_32_t1 = TR_44 ;
	7'h4c :
		RG_rl_32_t1 = TR_44 ;
	7'h4d :
		RG_rl_32_t1 = TR_44 ;
	7'h4e :
		RG_rl_32_t1 = TR_44 ;
	7'h4f :
		RG_rl_32_t1 = TR_44 ;
	7'h50 :
		RG_rl_32_t1 = TR_44 ;
	7'h51 :
		RG_rl_32_t1 = TR_44 ;
	7'h52 :
		RG_rl_32_t1 = TR_44 ;
	7'h53 :
		RG_rl_32_t1 = TR_44 ;
	7'h54 :
		RG_rl_32_t1 = TR_44 ;
	7'h55 :
		RG_rl_32_t1 = TR_44 ;
	7'h56 :
		RG_rl_32_t1 = TR_44 ;
	7'h57 :
		RG_rl_32_t1 = TR_44 ;
	7'h58 :
		RG_rl_32_t1 = TR_44 ;
	7'h59 :
		RG_rl_32_t1 = TR_44 ;
	7'h5a :
		RG_rl_32_t1 = TR_44 ;
	7'h5b :
		RG_rl_32_t1 = TR_44 ;
	7'h5c :
		RG_rl_32_t1 = TR_44 ;
	7'h5d :
		RG_rl_32_t1 = TR_44 ;
	7'h5e :
		RG_rl_32_t1 = TR_44 ;
	7'h5f :
		RG_rl_32_t1 = TR_44 ;
	7'h60 :
		RG_rl_32_t1 = TR_44 ;
	7'h61 :
		RG_rl_32_t1 = TR_44 ;
	7'h62 :
		RG_rl_32_t1 = TR_44 ;
	7'h63 :
		RG_rl_32_t1 = TR_44 ;
	7'h64 :
		RG_rl_32_t1 = TR_44 ;
	7'h65 :
		RG_rl_32_t1 = TR_44 ;
	7'h66 :
		RG_rl_32_t1 = TR_44 ;
	7'h67 :
		RG_rl_32_t1 = TR_44 ;
	7'h68 :
		RG_rl_32_t1 = TR_44 ;
	7'h69 :
		RG_rl_32_t1 = TR_44 ;
	7'h6a :
		RG_rl_32_t1 = TR_44 ;
	7'h6b :
		RG_rl_32_t1 = TR_44 ;
	7'h6c :
		RG_rl_32_t1 = TR_44 ;
	7'h6d :
		RG_rl_32_t1 = TR_44 ;
	7'h6e :
		RG_rl_32_t1 = TR_44 ;
	7'h6f :
		RG_rl_32_t1 = TR_44 ;
	7'h70 :
		RG_rl_32_t1 = TR_44 ;
	7'h71 :
		RG_rl_32_t1 = TR_44 ;
	7'h72 :
		RG_rl_32_t1 = TR_44 ;
	7'h73 :
		RG_rl_32_t1 = TR_44 ;
	7'h74 :
		RG_rl_32_t1 = TR_44 ;
	7'h75 :
		RG_rl_32_t1 = TR_44 ;
	7'h76 :
		RG_rl_32_t1 = TR_44 ;
	7'h77 :
		RG_rl_32_t1 = TR_44 ;
	7'h78 :
		RG_rl_32_t1 = TR_44 ;
	7'h79 :
		RG_rl_32_t1 = TR_44 ;
	7'h7a :
		RG_rl_32_t1 = TR_44 ;
	7'h7b :
		RG_rl_32_t1 = TR_44 ;
	7'h7c :
		RG_rl_32_t1 = TR_44 ;
	7'h7d :
		RG_rl_32_t1 = TR_44 ;
	7'h7e :
		RG_rl_32_t1 = TR_44 ;
	7'h7f :
		RG_rl_32_t1 = TR_44 ;
	default :
		RG_rl_32_t1 = 9'hx ;
	endcase
always @ ( RG_rl_32_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_215 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_32_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h20 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_32_t = ( ( { 9{ U_570 } } & RG_rl_215 )
		| ( { 9{ U_569 } } & RG_rl_32_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_32_en = ( U_570 | RG_rl_32_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_32_en )
		RG_rl_32 <= RG_rl_32_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_45 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_33_t1 = TR_45 ;
	7'h01 :
		RG_rl_33_t1 = TR_45 ;
	7'h02 :
		RG_rl_33_t1 = TR_45 ;
	7'h03 :
		RG_rl_33_t1 = TR_45 ;
	7'h04 :
		RG_rl_33_t1 = TR_45 ;
	7'h05 :
		RG_rl_33_t1 = TR_45 ;
	7'h06 :
		RG_rl_33_t1 = TR_45 ;
	7'h07 :
		RG_rl_33_t1 = TR_45 ;
	7'h08 :
		RG_rl_33_t1 = TR_45 ;
	7'h09 :
		RG_rl_33_t1 = TR_45 ;
	7'h0a :
		RG_rl_33_t1 = TR_45 ;
	7'h0b :
		RG_rl_33_t1 = TR_45 ;
	7'h0c :
		RG_rl_33_t1 = TR_45 ;
	7'h0d :
		RG_rl_33_t1 = TR_45 ;
	7'h0e :
		RG_rl_33_t1 = TR_45 ;
	7'h0f :
		RG_rl_33_t1 = TR_45 ;
	7'h10 :
		RG_rl_33_t1 = TR_45 ;
	7'h11 :
		RG_rl_33_t1 = TR_45 ;
	7'h12 :
		RG_rl_33_t1 = TR_45 ;
	7'h13 :
		RG_rl_33_t1 = TR_45 ;
	7'h14 :
		RG_rl_33_t1 = TR_45 ;
	7'h15 :
		RG_rl_33_t1 = TR_45 ;
	7'h16 :
		RG_rl_33_t1 = TR_45 ;
	7'h17 :
		RG_rl_33_t1 = TR_45 ;
	7'h18 :
		RG_rl_33_t1 = TR_45 ;
	7'h19 :
		RG_rl_33_t1 = TR_45 ;
	7'h1a :
		RG_rl_33_t1 = TR_45 ;
	7'h1b :
		RG_rl_33_t1 = TR_45 ;
	7'h1c :
		RG_rl_33_t1 = TR_45 ;
	7'h1d :
		RG_rl_33_t1 = TR_45 ;
	7'h1e :
		RG_rl_33_t1 = TR_45 ;
	7'h1f :
		RG_rl_33_t1 = TR_45 ;
	7'h20 :
		RG_rl_33_t1 = TR_45 ;
	7'h21 :
		RG_rl_33_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h22 :
		RG_rl_33_t1 = TR_45 ;
	7'h23 :
		RG_rl_33_t1 = TR_45 ;
	7'h24 :
		RG_rl_33_t1 = TR_45 ;
	7'h25 :
		RG_rl_33_t1 = TR_45 ;
	7'h26 :
		RG_rl_33_t1 = TR_45 ;
	7'h27 :
		RG_rl_33_t1 = TR_45 ;
	7'h28 :
		RG_rl_33_t1 = TR_45 ;
	7'h29 :
		RG_rl_33_t1 = TR_45 ;
	7'h2a :
		RG_rl_33_t1 = TR_45 ;
	7'h2b :
		RG_rl_33_t1 = TR_45 ;
	7'h2c :
		RG_rl_33_t1 = TR_45 ;
	7'h2d :
		RG_rl_33_t1 = TR_45 ;
	7'h2e :
		RG_rl_33_t1 = TR_45 ;
	7'h2f :
		RG_rl_33_t1 = TR_45 ;
	7'h30 :
		RG_rl_33_t1 = TR_45 ;
	7'h31 :
		RG_rl_33_t1 = TR_45 ;
	7'h32 :
		RG_rl_33_t1 = TR_45 ;
	7'h33 :
		RG_rl_33_t1 = TR_45 ;
	7'h34 :
		RG_rl_33_t1 = TR_45 ;
	7'h35 :
		RG_rl_33_t1 = TR_45 ;
	7'h36 :
		RG_rl_33_t1 = TR_45 ;
	7'h37 :
		RG_rl_33_t1 = TR_45 ;
	7'h38 :
		RG_rl_33_t1 = TR_45 ;
	7'h39 :
		RG_rl_33_t1 = TR_45 ;
	7'h3a :
		RG_rl_33_t1 = TR_45 ;
	7'h3b :
		RG_rl_33_t1 = TR_45 ;
	7'h3c :
		RG_rl_33_t1 = TR_45 ;
	7'h3d :
		RG_rl_33_t1 = TR_45 ;
	7'h3e :
		RG_rl_33_t1 = TR_45 ;
	7'h3f :
		RG_rl_33_t1 = TR_45 ;
	7'h40 :
		RG_rl_33_t1 = TR_45 ;
	7'h41 :
		RG_rl_33_t1 = TR_45 ;
	7'h42 :
		RG_rl_33_t1 = TR_45 ;
	7'h43 :
		RG_rl_33_t1 = TR_45 ;
	7'h44 :
		RG_rl_33_t1 = TR_45 ;
	7'h45 :
		RG_rl_33_t1 = TR_45 ;
	7'h46 :
		RG_rl_33_t1 = TR_45 ;
	7'h47 :
		RG_rl_33_t1 = TR_45 ;
	7'h48 :
		RG_rl_33_t1 = TR_45 ;
	7'h49 :
		RG_rl_33_t1 = TR_45 ;
	7'h4a :
		RG_rl_33_t1 = TR_45 ;
	7'h4b :
		RG_rl_33_t1 = TR_45 ;
	7'h4c :
		RG_rl_33_t1 = TR_45 ;
	7'h4d :
		RG_rl_33_t1 = TR_45 ;
	7'h4e :
		RG_rl_33_t1 = TR_45 ;
	7'h4f :
		RG_rl_33_t1 = TR_45 ;
	7'h50 :
		RG_rl_33_t1 = TR_45 ;
	7'h51 :
		RG_rl_33_t1 = TR_45 ;
	7'h52 :
		RG_rl_33_t1 = TR_45 ;
	7'h53 :
		RG_rl_33_t1 = TR_45 ;
	7'h54 :
		RG_rl_33_t1 = TR_45 ;
	7'h55 :
		RG_rl_33_t1 = TR_45 ;
	7'h56 :
		RG_rl_33_t1 = TR_45 ;
	7'h57 :
		RG_rl_33_t1 = TR_45 ;
	7'h58 :
		RG_rl_33_t1 = TR_45 ;
	7'h59 :
		RG_rl_33_t1 = TR_45 ;
	7'h5a :
		RG_rl_33_t1 = TR_45 ;
	7'h5b :
		RG_rl_33_t1 = TR_45 ;
	7'h5c :
		RG_rl_33_t1 = TR_45 ;
	7'h5d :
		RG_rl_33_t1 = TR_45 ;
	7'h5e :
		RG_rl_33_t1 = TR_45 ;
	7'h5f :
		RG_rl_33_t1 = TR_45 ;
	7'h60 :
		RG_rl_33_t1 = TR_45 ;
	7'h61 :
		RG_rl_33_t1 = TR_45 ;
	7'h62 :
		RG_rl_33_t1 = TR_45 ;
	7'h63 :
		RG_rl_33_t1 = TR_45 ;
	7'h64 :
		RG_rl_33_t1 = TR_45 ;
	7'h65 :
		RG_rl_33_t1 = TR_45 ;
	7'h66 :
		RG_rl_33_t1 = TR_45 ;
	7'h67 :
		RG_rl_33_t1 = TR_45 ;
	7'h68 :
		RG_rl_33_t1 = TR_45 ;
	7'h69 :
		RG_rl_33_t1 = TR_45 ;
	7'h6a :
		RG_rl_33_t1 = TR_45 ;
	7'h6b :
		RG_rl_33_t1 = TR_45 ;
	7'h6c :
		RG_rl_33_t1 = TR_45 ;
	7'h6d :
		RG_rl_33_t1 = TR_45 ;
	7'h6e :
		RG_rl_33_t1 = TR_45 ;
	7'h6f :
		RG_rl_33_t1 = TR_45 ;
	7'h70 :
		RG_rl_33_t1 = TR_45 ;
	7'h71 :
		RG_rl_33_t1 = TR_45 ;
	7'h72 :
		RG_rl_33_t1 = TR_45 ;
	7'h73 :
		RG_rl_33_t1 = TR_45 ;
	7'h74 :
		RG_rl_33_t1 = TR_45 ;
	7'h75 :
		RG_rl_33_t1 = TR_45 ;
	7'h76 :
		RG_rl_33_t1 = TR_45 ;
	7'h77 :
		RG_rl_33_t1 = TR_45 ;
	7'h78 :
		RG_rl_33_t1 = TR_45 ;
	7'h79 :
		RG_rl_33_t1 = TR_45 ;
	7'h7a :
		RG_rl_33_t1 = TR_45 ;
	7'h7b :
		RG_rl_33_t1 = TR_45 ;
	7'h7c :
		RG_rl_33_t1 = TR_45 ;
	7'h7d :
		RG_rl_33_t1 = TR_45 ;
	7'h7e :
		RG_rl_33_t1 = TR_45 ;
	7'h7f :
		RG_rl_33_t1 = TR_45 ;
	default :
		RG_rl_33_t1 = 9'hx ;
	endcase
always @ ( RG_rl_33_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_216 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_33_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h21 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_33_t = ( ( { 9{ U_570 } } & RG_rl_216 )
		| ( { 9{ U_569 } } & RG_rl_33_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_33_en = ( U_570 | RG_rl_33_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_33_en )
		RG_rl_33 <= RG_rl_33_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_46 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_34_t1 = TR_46 ;
	7'h01 :
		RG_rl_34_t1 = TR_46 ;
	7'h02 :
		RG_rl_34_t1 = TR_46 ;
	7'h03 :
		RG_rl_34_t1 = TR_46 ;
	7'h04 :
		RG_rl_34_t1 = TR_46 ;
	7'h05 :
		RG_rl_34_t1 = TR_46 ;
	7'h06 :
		RG_rl_34_t1 = TR_46 ;
	7'h07 :
		RG_rl_34_t1 = TR_46 ;
	7'h08 :
		RG_rl_34_t1 = TR_46 ;
	7'h09 :
		RG_rl_34_t1 = TR_46 ;
	7'h0a :
		RG_rl_34_t1 = TR_46 ;
	7'h0b :
		RG_rl_34_t1 = TR_46 ;
	7'h0c :
		RG_rl_34_t1 = TR_46 ;
	7'h0d :
		RG_rl_34_t1 = TR_46 ;
	7'h0e :
		RG_rl_34_t1 = TR_46 ;
	7'h0f :
		RG_rl_34_t1 = TR_46 ;
	7'h10 :
		RG_rl_34_t1 = TR_46 ;
	7'h11 :
		RG_rl_34_t1 = TR_46 ;
	7'h12 :
		RG_rl_34_t1 = TR_46 ;
	7'h13 :
		RG_rl_34_t1 = TR_46 ;
	7'h14 :
		RG_rl_34_t1 = TR_46 ;
	7'h15 :
		RG_rl_34_t1 = TR_46 ;
	7'h16 :
		RG_rl_34_t1 = TR_46 ;
	7'h17 :
		RG_rl_34_t1 = TR_46 ;
	7'h18 :
		RG_rl_34_t1 = TR_46 ;
	7'h19 :
		RG_rl_34_t1 = TR_46 ;
	7'h1a :
		RG_rl_34_t1 = TR_46 ;
	7'h1b :
		RG_rl_34_t1 = TR_46 ;
	7'h1c :
		RG_rl_34_t1 = TR_46 ;
	7'h1d :
		RG_rl_34_t1 = TR_46 ;
	7'h1e :
		RG_rl_34_t1 = TR_46 ;
	7'h1f :
		RG_rl_34_t1 = TR_46 ;
	7'h20 :
		RG_rl_34_t1 = TR_46 ;
	7'h21 :
		RG_rl_34_t1 = TR_46 ;
	7'h22 :
		RG_rl_34_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h23 :
		RG_rl_34_t1 = TR_46 ;
	7'h24 :
		RG_rl_34_t1 = TR_46 ;
	7'h25 :
		RG_rl_34_t1 = TR_46 ;
	7'h26 :
		RG_rl_34_t1 = TR_46 ;
	7'h27 :
		RG_rl_34_t1 = TR_46 ;
	7'h28 :
		RG_rl_34_t1 = TR_46 ;
	7'h29 :
		RG_rl_34_t1 = TR_46 ;
	7'h2a :
		RG_rl_34_t1 = TR_46 ;
	7'h2b :
		RG_rl_34_t1 = TR_46 ;
	7'h2c :
		RG_rl_34_t1 = TR_46 ;
	7'h2d :
		RG_rl_34_t1 = TR_46 ;
	7'h2e :
		RG_rl_34_t1 = TR_46 ;
	7'h2f :
		RG_rl_34_t1 = TR_46 ;
	7'h30 :
		RG_rl_34_t1 = TR_46 ;
	7'h31 :
		RG_rl_34_t1 = TR_46 ;
	7'h32 :
		RG_rl_34_t1 = TR_46 ;
	7'h33 :
		RG_rl_34_t1 = TR_46 ;
	7'h34 :
		RG_rl_34_t1 = TR_46 ;
	7'h35 :
		RG_rl_34_t1 = TR_46 ;
	7'h36 :
		RG_rl_34_t1 = TR_46 ;
	7'h37 :
		RG_rl_34_t1 = TR_46 ;
	7'h38 :
		RG_rl_34_t1 = TR_46 ;
	7'h39 :
		RG_rl_34_t1 = TR_46 ;
	7'h3a :
		RG_rl_34_t1 = TR_46 ;
	7'h3b :
		RG_rl_34_t1 = TR_46 ;
	7'h3c :
		RG_rl_34_t1 = TR_46 ;
	7'h3d :
		RG_rl_34_t1 = TR_46 ;
	7'h3e :
		RG_rl_34_t1 = TR_46 ;
	7'h3f :
		RG_rl_34_t1 = TR_46 ;
	7'h40 :
		RG_rl_34_t1 = TR_46 ;
	7'h41 :
		RG_rl_34_t1 = TR_46 ;
	7'h42 :
		RG_rl_34_t1 = TR_46 ;
	7'h43 :
		RG_rl_34_t1 = TR_46 ;
	7'h44 :
		RG_rl_34_t1 = TR_46 ;
	7'h45 :
		RG_rl_34_t1 = TR_46 ;
	7'h46 :
		RG_rl_34_t1 = TR_46 ;
	7'h47 :
		RG_rl_34_t1 = TR_46 ;
	7'h48 :
		RG_rl_34_t1 = TR_46 ;
	7'h49 :
		RG_rl_34_t1 = TR_46 ;
	7'h4a :
		RG_rl_34_t1 = TR_46 ;
	7'h4b :
		RG_rl_34_t1 = TR_46 ;
	7'h4c :
		RG_rl_34_t1 = TR_46 ;
	7'h4d :
		RG_rl_34_t1 = TR_46 ;
	7'h4e :
		RG_rl_34_t1 = TR_46 ;
	7'h4f :
		RG_rl_34_t1 = TR_46 ;
	7'h50 :
		RG_rl_34_t1 = TR_46 ;
	7'h51 :
		RG_rl_34_t1 = TR_46 ;
	7'h52 :
		RG_rl_34_t1 = TR_46 ;
	7'h53 :
		RG_rl_34_t1 = TR_46 ;
	7'h54 :
		RG_rl_34_t1 = TR_46 ;
	7'h55 :
		RG_rl_34_t1 = TR_46 ;
	7'h56 :
		RG_rl_34_t1 = TR_46 ;
	7'h57 :
		RG_rl_34_t1 = TR_46 ;
	7'h58 :
		RG_rl_34_t1 = TR_46 ;
	7'h59 :
		RG_rl_34_t1 = TR_46 ;
	7'h5a :
		RG_rl_34_t1 = TR_46 ;
	7'h5b :
		RG_rl_34_t1 = TR_46 ;
	7'h5c :
		RG_rl_34_t1 = TR_46 ;
	7'h5d :
		RG_rl_34_t1 = TR_46 ;
	7'h5e :
		RG_rl_34_t1 = TR_46 ;
	7'h5f :
		RG_rl_34_t1 = TR_46 ;
	7'h60 :
		RG_rl_34_t1 = TR_46 ;
	7'h61 :
		RG_rl_34_t1 = TR_46 ;
	7'h62 :
		RG_rl_34_t1 = TR_46 ;
	7'h63 :
		RG_rl_34_t1 = TR_46 ;
	7'h64 :
		RG_rl_34_t1 = TR_46 ;
	7'h65 :
		RG_rl_34_t1 = TR_46 ;
	7'h66 :
		RG_rl_34_t1 = TR_46 ;
	7'h67 :
		RG_rl_34_t1 = TR_46 ;
	7'h68 :
		RG_rl_34_t1 = TR_46 ;
	7'h69 :
		RG_rl_34_t1 = TR_46 ;
	7'h6a :
		RG_rl_34_t1 = TR_46 ;
	7'h6b :
		RG_rl_34_t1 = TR_46 ;
	7'h6c :
		RG_rl_34_t1 = TR_46 ;
	7'h6d :
		RG_rl_34_t1 = TR_46 ;
	7'h6e :
		RG_rl_34_t1 = TR_46 ;
	7'h6f :
		RG_rl_34_t1 = TR_46 ;
	7'h70 :
		RG_rl_34_t1 = TR_46 ;
	7'h71 :
		RG_rl_34_t1 = TR_46 ;
	7'h72 :
		RG_rl_34_t1 = TR_46 ;
	7'h73 :
		RG_rl_34_t1 = TR_46 ;
	7'h74 :
		RG_rl_34_t1 = TR_46 ;
	7'h75 :
		RG_rl_34_t1 = TR_46 ;
	7'h76 :
		RG_rl_34_t1 = TR_46 ;
	7'h77 :
		RG_rl_34_t1 = TR_46 ;
	7'h78 :
		RG_rl_34_t1 = TR_46 ;
	7'h79 :
		RG_rl_34_t1 = TR_46 ;
	7'h7a :
		RG_rl_34_t1 = TR_46 ;
	7'h7b :
		RG_rl_34_t1 = TR_46 ;
	7'h7c :
		RG_rl_34_t1 = TR_46 ;
	7'h7d :
		RG_rl_34_t1 = TR_46 ;
	7'h7e :
		RG_rl_34_t1 = TR_46 ;
	7'h7f :
		RG_rl_34_t1 = TR_46 ;
	default :
		RG_rl_34_t1 = 9'hx ;
	endcase
always @ ( RG_rl_34_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_217 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_34_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h22 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_34_t = ( ( { 9{ U_570 } } & RG_rl_217 )
		| ( { 9{ U_569 } } & RG_rl_34_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_34_en = ( U_570 | RG_rl_34_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_34_en )
		RG_rl_34 <= RG_rl_34_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_47 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_35_t1 = TR_47 ;
	7'h01 :
		RG_rl_35_t1 = TR_47 ;
	7'h02 :
		RG_rl_35_t1 = TR_47 ;
	7'h03 :
		RG_rl_35_t1 = TR_47 ;
	7'h04 :
		RG_rl_35_t1 = TR_47 ;
	7'h05 :
		RG_rl_35_t1 = TR_47 ;
	7'h06 :
		RG_rl_35_t1 = TR_47 ;
	7'h07 :
		RG_rl_35_t1 = TR_47 ;
	7'h08 :
		RG_rl_35_t1 = TR_47 ;
	7'h09 :
		RG_rl_35_t1 = TR_47 ;
	7'h0a :
		RG_rl_35_t1 = TR_47 ;
	7'h0b :
		RG_rl_35_t1 = TR_47 ;
	7'h0c :
		RG_rl_35_t1 = TR_47 ;
	7'h0d :
		RG_rl_35_t1 = TR_47 ;
	7'h0e :
		RG_rl_35_t1 = TR_47 ;
	7'h0f :
		RG_rl_35_t1 = TR_47 ;
	7'h10 :
		RG_rl_35_t1 = TR_47 ;
	7'h11 :
		RG_rl_35_t1 = TR_47 ;
	7'h12 :
		RG_rl_35_t1 = TR_47 ;
	7'h13 :
		RG_rl_35_t1 = TR_47 ;
	7'h14 :
		RG_rl_35_t1 = TR_47 ;
	7'h15 :
		RG_rl_35_t1 = TR_47 ;
	7'h16 :
		RG_rl_35_t1 = TR_47 ;
	7'h17 :
		RG_rl_35_t1 = TR_47 ;
	7'h18 :
		RG_rl_35_t1 = TR_47 ;
	7'h19 :
		RG_rl_35_t1 = TR_47 ;
	7'h1a :
		RG_rl_35_t1 = TR_47 ;
	7'h1b :
		RG_rl_35_t1 = TR_47 ;
	7'h1c :
		RG_rl_35_t1 = TR_47 ;
	7'h1d :
		RG_rl_35_t1 = TR_47 ;
	7'h1e :
		RG_rl_35_t1 = TR_47 ;
	7'h1f :
		RG_rl_35_t1 = TR_47 ;
	7'h20 :
		RG_rl_35_t1 = TR_47 ;
	7'h21 :
		RG_rl_35_t1 = TR_47 ;
	7'h22 :
		RG_rl_35_t1 = TR_47 ;
	7'h23 :
		RG_rl_35_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h24 :
		RG_rl_35_t1 = TR_47 ;
	7'h25 :
		RG_rl_35_t1 = TR_47 ;
	7'h26 :
		RG_rl_35_t1 = TR_47 ;
	7'h27 :
		RG_rl_35_t1 = TR_47 ;
	7'h28 :
		RG_rl_35_t1 = TR_47 ;
	7'h29 :
		RG_rl_35_t1 = TR_47 ;
	7'h2a :
		RG_rl_35_t1 = TR_47 ;
	7'h2b :
		RG_rl_35_t1 = TR_47 ;
	7'h2c :
		RG_rl_35_t1 = TR_47 ;
	7'h2d :
		RG_rl_35_t1 = TR_47 ;
	7'h2e :
		RG_rl_35_t1 = TR_47 ;
	7'h2f :
		RG_rl_35_t1 = TR_47 ;
	7'h30 :
		RG_rl_35_t1 = TR_47 ;
	7'h31 :
		RG_rl_35_t1 = TR_47 ;
	7'h32 :
		RG_rl_35_t1 = TR_47 ;
	7'h33 :
		RG_rl_35_t1 = TR_47 ;
	7'h34 :
		RG_rl_35_t1 = TR_47 ;
	7'h35 :
		RG_rl_35_t1 = TR_47 ;
	7'h36 :
		RG_rl_35_t1 = TR_47 ;
	7'h37 :
		RG_rl_35_t1 = TR_47 ;
	7'h38 :
		RG_rl_35_t1 = TR_47 ;
	7'h39 :
		RG_rl_35_t1 = TR_47 ;
	7'h3a :
		RG_rl_35_t1 = TR_47 ;
	7'h3b :
		RG_rl_35_t1 = TR_47 ;
	7'h3c :
		RG_rl_35_t1 = TR_47 ;
	7'h3d :
		RG_rl_35_t1 = TR_47 ;
	7'h3e :
		RG_rl_35_t1 = TR_47 ;
	7'h3f :
		RG_rl_35_t1 = TR_47 ;
	7'h40 :
		RG_rl_35_t1 = TR_47 ;
	7'h41 :
		RG_rl_35_t1 = TR_47 ;
	7'h42 :
		RG_rl_35_t1 = TR_47 ;
	7'h43 :
		RG_rl_35_t1 = TR_47 ;
	7'h44 :
		RG_rl_35_t1 = TR_47 ;
	7'h45 :
		RG_rl_35_t1 = TR_47 ;
	7'h46 :
		RG_rl_35_t1 = TR_47 ;
	7'h47 :
		RG_rl_35_t1 = TR_47 ;
	7'h48 :
		RG_rl_35_t1 = TR_47 ;
	7'h49 :
		RG_rl_35_t1 = TR_47 ;
	7'h4a :
		RG_rl_35_t1 = TR_47 ;
	7'h4b :
		RG_rl_35_t1 = TR_47 ;
	7'h4c :
		RG_rl_35_t1 = TR_47 ;
	7'h4d :
		RG_rl_35_t1 = TR_47 ;
	7'h4e :
		RG_rl_35_t1 = TR_47 ;
	7'h4f :
		RG_rl_35_t1 = TR_47 ;
	7'h50 :
		RG_rl_35_t1 = TR_47 ;
	7'h51 :
		RG_rl_35_t1 = TR_47 ;
	7'h52 :
		RG_rl_35_t1 = TR_47 ;
	7'h53 :
		RG_rl_35_t1 = TR_47 ;
	7'h54 :
		RG_rl_35_t1 = TR_47 ;
	7'h55 :
		RG_rl_35_t1 = TR_47 ;
	7'h56 :
		RG_rl_35_t1 = TR_47 ;
	7'h57 :
		RG_rl_35_t1 = TR_47 ;
	7'h58 :
		RG_rl_35_t1 = TR_47 ;
	7'h59 :
		RG_rl_35_t1 = TR_47 ;
	7'h5a :
		RG_rl_35_t1 = TR_47 ;
	7'h5b :
		RG_rl_35_t1 = TR_47 ;
	7'h5c :
		RG_rl_35_t1 = TR_47 ;
	7'h5d :
		RG_rl_35_t1 = TR_47 ;
	7'h5e :
		RG_rl_35_t1 = TR_47 ;
	7'h5f :
		RG_rl_35_t1 = TR_47 ;
	7'h60 :
		RG_rl_35_t1 = TR_47 ;
	7'h61 :
		RG_rl_35_t1 = TR_47 ;
	7'h62 :
		RG_rl_35_t1 = TR_47 ;
	7'h63 :
		RG_rl_35_t1 = TR_47 ;
	7'h64 :
		RG_rl_35_t1 = TR_47 ;
	7'h65 :
		RG_rl_35_t1 = TR_47 ;
	7'h66 :
		RG_rl_35_t1 = TR_47 ;
	7'h67 :
		RG_rl_35_t1 = TR_47 ;
	7'h68 :
		RG_rl_35_t1 = TR_47 ;
	7'h69 :
		RG_rl_35_t1 = TR_47 ;
	7'h6a :
		RG_rl_35_t1 = TR_47 ;
	7'h6b :
		RG_rl_35_t1 = TR_47 ;
	7'h6c :
		RG_rl_35_t1 = TR_47 ;
	7'h6d :
		RG_rl_35_t1 = TR_47 ;
	7'h6e :
		RG_rl_35_t1 = TR_47 ;
	7'h6f :
		RG_rl_35_t1 = TR_47 ;
	7'h70 :
		RG_rl_35_t1 = TR_47 ;
	7'h71 :
		RG_rl_35_t1 = TR_47 ;
	7'h72 :
		RG_rl_35_t1 = TR_47 ;
	7'h73 :
		RG_rl_35_t1 = TR_47 ;
	7'h74 :
		RG_rl_35_t1 = TR_47 ;
	7'h75 :
		RG_rl_35_t1 = TR_47 ;
	7'h76 :
		RG_rl_35_t1 = TR_47 ;
	7'h77 :
		RG_rl_35_t1 = TR_47 ;
	7'h78 :
		RG_rl_35_t1 = TR_47 ;
	7'h79 :
		RG_rl_35_t1 = TR_47 ;
	7'h7a :
		RG_rl_35_t1 = TR_47 ;
	7'h7b :
		RG_rl_35_t1 = TR_47 ;
	7'h7c :
		RG_rl_35_t1 = TR_47 ;
	7'h7d :
		RG_rl_35_t1 = TR_47 ;
	7'h7e :
		RG_rl_35_t1 = TR_47 ;
	7'h7f :
		RG_rl_35_t1 = TR_47 ;
	default :
		RG_rl_35_t1 = 9'hx ;
	endcase
always @ ( RG_rl_35_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_218 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_35_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h23 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_35_t = ( ( { 9{ U_570 } } & RG_rl_218 )
		| ( { 9{ U_569 } } & RG_rl_35_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_35_en = ( U_570 | RG_rl_35_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_35_en )
		RG_rl_35 <= RG_rl_35_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_48 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_36_t1 = TR_48 ;
	7'h01 :
		RG_rl_36_t1 = TR_48 ;
	7'h02 :
		RG_rl_36_t1 = TR_48 ;
	7'h03 :
		RG_rl_36_t1 = TR_48 ;
	7'h04 :
		RG_rl_36_t1 = TR_48 ;
	7'h05 :
		RG_rl_36_t1 = TR_48 ;
	7'h06 :
		RG_rl_36_t1 = TR_48 ;
	7'h07 :
		RG_rl_36_t1 = TR_48 ;
	7'h08 :
		RG_rl_36_t1 = TR_48 ;
	7'h09 :
		RG_rl_36_t1 = TR_48 ;
	7'h0a :
		RG_rl_36_t1 = TR_48 ;
	7'h0b :
		RG_rl_36_t1 = TR_48 ;
	7'h0c :
		RG_rl_36_t1 = TR_48 ;
	7'h0d :
		RG_rl_36_t1 = TR_48 ;
	7'h0e :
		RG_rl_36_t1 = TR_48 ;
	7'h0f :
		RG_rl_36_t1 = TR_48 ;
	7'h10 :
		RG_rl_36_t1 = TR_48 ;
	7'h11 :
		RG_rl_36_t1 = TR_48 ;
	7'h12 :
		RG_rl_36_t1 = TR_48 ;
	7'h13 :
		RG_rl_36_t1 = TR_48 ;
	7'h14 :
		RG_rl_36_t1 = TR_48 ;
	7'h15 :
		RG_rl_36_t1 = TR_48 ;
	7'h16 :
		RG_rl_36_t1 = TR_48 ;
	7'h17 :
		RG_rl_36_t1 = TR_48 ;
	7'h18 :
		RG_rl_36_t1 = TR_48 ;
	7'h19 :
		RG_rl_36_t1 = TR_48 ;
	7'h1a :
		RG_rl_36_t1 = TR_48 ;
	7'h1b :
		RG_rl_36_t1 = TR_48 ;
	7'h1c :
		RG_rl_36_t1 = TR_48 ;
	7'h1d :
		RG_rl_36_t1 = TR_48 ;
	7'h1e :
		RG_rl_36_t1 = TR_48 ;
	7'h1f :
		RG_rl_36_t1 = TR_48 ;
	7'h20 :
		RG_rl_36_t1 = TR_48 ;
	7'h21 :
		RG_rl_36_t1 = TR_48 ;
	7'h22 :
		RG_rl_36_t1 = TR_48 ;
	7'h23 :
		RG_rl_36_t1 = TR_48 ;
	7'h24 :
		RG_rl_36_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h25 :
		RG_rl_36_t1 = TR_48 ;
	7'h26 :
		RG_rl_36_t1 = TR_48 ;
	7'h27 :
		RG_rl_36_t1 = TR_48 ;
	7'h28 :
		RG_rl_36_t1 = TR_48 ;
	7'h29 :
		RG_rl_36_t1 = TR_48 ;
	7'h2a :
		RG_rl_36_t1 = TR_48 ;
	7'h2b :
		RG_rl_36_t1 = TR_48 ;
	7'h2c :
		RG_rl_36_t1 = TR_48 ;
	7'h2d :
		RG_rl_36_t1 = TR_48 ;
	7'h2e :
		RG_rl_36_t1 = TR_48 ;
	7'h2f :
		RG_rl_36_t1 = TR_48 ;
	7'h30 :
		RG_rl_36_t1 = TR_48 ;
	7'h31 :
		RG_rl_36_t1 = TR_48 ;
	7'h32 :
		RG_rl_36_t1 = TR_48 ;
	7'h33 :
		RG_rl_36_t1 = TR_48 ;
	7'h34 :
		RG_rl_36_t1 = TR_48 ;
	7'h35 :
		RG_rl_36_t1 = TR_48 ;
	7'h36 :
		RG_rl_36_t1 = TR_48 ;
	7'h37 :
		RG_rl_36_t1 = TR_48 ;
	7'h38 :
		RG_rl_36_t1 = TR_48 ;
	7'h39 :
		RG_rl_36_t1 = TR_48 ;
	7'h3a :
		RG_rl_36_t1 = TR_48 ;
	7'h3b :
		RG_rl_36_t1 = TR_48 ;
	7'h3c :
		RG_rl_36_t1 = TR_48 ;
	7'h3d :
		RG_rl_36_t1 = TR_48 ;
	7'h3e :
		RG_rl_36_t1 = TR_48 ;
	7'h3f :
		RG_rl_36_t1 = TR_48 ;
	7'h40 :
		RG_rl_36_t1 = TR_48 ;
	7'h41 :
		RG_rl_36_t1 = TR_48 ;
	7'h42 :
		RG_rl_36_t1 = TR_48 ;
	7'h43 :
		RG_rl_36_t1 = TR_48 ;
	7'h44 :
		RG_rl_36_t1 = TR_48 ;
	7'h45 :
		RG_rl_36_t1 = TR_48 ;
	7'h46 :
		RG_rl_36_t1 = TR_48 ;
	7'h47 :
		RG_rl_36_t1 = TR_48 ;
	7'h48 :
		RG_rl_36_t1 = TR_48 ;
	7'h49 :
		RG_rl_36_t1 = TR_48 ;
	7'h4a :
		RG_rl_36_t1 = TR_48 ;
	7'h4b :
		RG_rl_36_t1 = TR_48 ;
	7'h4c :
		RG_rl_36_t1 = TR_48 ;
	7'h4d :
		RG_rl_36_t1 = TR_48 ;
	7'h4e :
		RG_rl_36_t1 = TR_48 ;
	7'h4f :
		RG_rl_36_t1 = TR_48 ;
	7'h50 :
		RG_rl_36_t1 = TR_48 ;
	7'h51 :
		RG_rl_36_t1 = TR_48 ;
	7'h52 :
		RG_rl_36_t1 = TR_48 ;
	7'h53 :
		RG_rl_36_t1 = TR_48 ;
	7'h54 :
		RG_rl_36_t1 = TR_48 ;
	7'h55 :
		RG_rl_36_t1 = TR_48 ;
	7'h56 :
		RG_rl_36_t1 = TR_48 ;
	7'h57 :
		RG_rl_36_t1 = TR_48 ;
	7'h58 :
		RG_rl_36_t1 = TR_48 ;
	7'h59 :
		RG_rl_36_t1 = TR_48 ;
	7'h5a :
		RG_rl_36_t1 = TR_48 ;
	7'h5b :
		RG_rl_36_t1 = TR_48 ;
	7'h5c :
		RG_rl_36_t1 = TR_48 ;
	7'h5d :
		RG_rl_36_t1 = TR_48 ;
	7'h5e :
		RG_rl_36_t1 = TR_48 ;
	7'h5f :
		RG_rl_36_t1 = TR_48 ;
	7'h60 :
		RG_rl_36_t1 = TR_48 ;
	7'h61 :
		RG_rl_36_t1 = TR_48 ;
	7'h62 :
		RG_rl_36_t1 = TR_48 ;
	7'h63 :
		RG_rl_36_t1 = TR_48 ;
	7'h64 :
		RG_rl_36_t1 = TR_48 ;
	7'h65 :
		RG_rl_36_t1 = TR_48 ;
	7'h66 :
		RG_rl_36_t1 = TR_48 ;
	7'h67 :
		RG_rl_36_t1 = TR_48 ;
	7'h68 :
		RG_rl_36_t1 = TR_48 ;
	7'h69 :
		RG_rl_36_t1 = TR_48 ;
	7'h6a :
		RG_rl_36_t1 = TR_48 ;
	7'h6b :
		RG_rl_36_t1 = TR_48 ;
	7'h6c :
		RG_rl_36_t1 = TR_48 ;
	7'h6d :
		RG_rl_36_t1 = TR_48 ;
	7'h6e :
		RG_rl_36_t1 = TR_48 ;
	7'h6f :
		RG_rl_36_t1 = TR_48 ;
	7'h70 :
		RG_rl_36_t1 = TR_48 ;
	7'h71 :
		RG_rl_36_t1 = TR_48 ;
	7'h72 :
		RG_rl_36_t1 = TR_48 ;
	7'h73 :
		RG_rl_36_t1 = TR_48 ;
	7'h74 :
		RG_rl_36_t1 = TR_48 ;
	7'h75 :
		RG_rl_36_t1 = TR_48 ;
	7'h76 :
		RG_rl_36_t1 = TR_48 ;
	7'h77 :
		RG_rl_36_t1 = TR_48 ;
	7'h78 :
		RG_rl_36_t1 = TR_48 ;
	7'h79 :
		RG_rl_36_t1 = TR_48 ;
	7'h7a :
		RG_rl_36_t1 = TR_48 ;
	7'h7b :
		RG_rl_36_t1 = TR_48 ;
	7'h7c :
		RG_rl_36_t1 = TR_48 ;
	7'h7d :
		RG_rl_36_t1 = TR_48 ;
	7'h7e :
		RG_rl_36_t1 = TR_48 ;
	7'h7f :
		RG_rl_36_t1 = TR_48 ;
	default :
		RG_rl_36_t1 = 9'hx ;
	endcase
always @ ( RG_rl_36_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_219 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_36_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h24 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_36_t = ( ( { 9{ U_570 } } & RG_rl_219 )
		| ( { 9{ U_569 } } & RG_rl_36_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_36_en = ( U_570 | RG_rl_36_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_36_en )
		RG_rl_36 <= RG_rl_36_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_49 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_37_t1 = TR_49 ;
	7'h01 :
		RG_rl_37_t1 = TR_49 ;
	7'h02 :
		RG_rl_37_t1 = TR_49 ;
	7'h03 :
		RG_rl_37_t1 = TR_49 ;
	7'h04 :
		RG_rl_37_t1 = TR_49 ;
	7'h05 :
		RG_rl_37_t1 = TR_49 ;
	7'h06 :
		RG_rl_37_t1 = TR_49 ;
	7'h07 :
		RG_rl_37_t1 = TR_49 ;
	7'h08 :
		RG_rl_37_t1 = TR_49 ;
	7'h09 :
		RG_rl_37_t1 = TR_49 ;
	7'h0a :
		RG_rl_37_t1 = TR_49 ;
	7'h0b :
		RG_rl_37_t1 = TR_49 ;
	7'h0c :
		RG_rl_37_t1 = TR_49 ;
	7'h0d :
		RG_rl_37_t1 = TR_49 ;
	7'h0e :
		RG_rl_37_t1 = TR_49 ;
	7'h0f :
		RG_rl_37_t1 = TR_49 ;
	7'h10 :
		RG_rl_37_t1 = TR_49 ;
	7'h11 :
		RG_rl_37_t1 = TR_49 ;
	7'h12 :
		RG_rl_37_t1 = TR_49 ;
	7'h13 :
		RG_rl_37_t1 = TR_49 ;
	7'h14 :
		RG_rl_37_t1 = TR_49 ;
	7'h15 :
		RG_rl_37_t1 = TR_49 ;
	7'h16 :
		RG_rl_37_t1 = TR_49 ;
	7'h17 :
		RG_rl_37_t1 = TR_49 ;
	7'h18 :
		RG_rl_37_t1 = TR_49 ;
	7'h19 :
		RG_rl_37_t1 = TR_49 ;
	7'h1a :
		RG_rl_37_t1 = TR_49 ;
	7'h1b :
		RG_rl_37_t1 = TR_49 ;
	7'h1c :
		RG_rl_37_t1 = TR_49 ;
	7'h1d :
		RG_rl_37_t1 = TR_49 ;
	7'h1e :
		RG_rl_37_t1 = TR_49 ;
	7'h1f :
		RG_rl_37_t1 = TR_49 ;
	7'h20 :
		RG_rl_37_t1 = TR_49 ;
	7'h21 :
		RG_rl_37_t1 = TR_49 ;
	7'h22 :
		RG_rl_37_t1 = TR_49 ;
	7'h23 :
		RG_rl_37_t1 = TR_49 ;
	7'h24 :
		RG_rl_37_t1 = TR_49 ;
	7'h25 :
		RG_rl_37_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h26 :
		RG_rl_37_t1 = TR_49 ;
	7'h27 :
		RG_rl_37_t1 = TR_49 ;
	7'h28 :
		RG_rl_37_t1 = TR_49 ;
	7'h29 :
		RG_rl_37_t1 = TR_49 ;
	7'h2a :
		RG_rl_37_t1 = TR_49 ;
	7'h2b :
		RG_rl_37_t1 = TR_49 ;
	7'h2c :
		RG_rl_37_t1 = TR_49 ;
	7'h2d :
		RG_rl_37_t1 = TR_49 ;
	7'h2e :
		RG_rl_37_t1 = TR_49 ;
	7'h2f :
		RG_rl_37_t1 = TR_49 ;
	7'h30 :
		RG_rl_37_t1 = TR_49 ;
	7'h31 :
		RG_rl_37_t1 = TR_49 ;
	7'h32 :
		RG_rl_37_t1 = TR_49 ;
	7'h33 :
		RG_rl_37_t1 = TR_49 ;
	7'h34 :
		RG_rl_37_t1 = TR_49 ;
	7'h35 :
		RG_rl_37_t1 = TR_49 ;
	7'h36 :
		RG_rl_37_t1 = TR_49 ;
	7'h37 :
		RG_rl_37_t1 = TR_49 ;
	7'h38 :
		RG_rl_37_t1 = TR_49 ;
	7'h39 :
		RG_rl_37_t1 = TR_49 ;
	7'h3a :
		RG_rl_37_t1 = TR_49 ;
	7'h3b :
		RG_rl_37_t1 = TR_49 ;
	7'h3c :
		RG_rl_37_t1 = TR_49 ;
	7'h3d :
		RG_rl_37_t1 = TR_49 ;
	7'h3e :
		RG_rl_37_t1 = TR_49 ;
	7'h3f :
		RG_rl_37_t1 = TR_49 ;
	7'h40 :
		RG_rl_37_t1 = TR_49 ;
	7'h41 :
		RG_rl_37_t1 = TR_49 ;
	7'h42 :
		RG_rl_37_t1 = TR_49 ;
	7'h43 :
		RG_rl_37_t1 = TR_49 ;
	7'h44 :
		RG_rl_37_t1 = TR_49 ;
	7'h45 :
		RG_rl_37_t1 = TR_49 ;
	7'h46 :
		RG_rl_37_t1 = TR_49 ;
	7'h47 :
		RG_rl_37_t1 = TR_49 ;
	7'h48 :
		RG_rl_37_t1 = TR_49 ;
	7'h49 :
		RG_rl_37_t1 = TR_49 ;
	7'h4a :
		RG_rl_37_t1 = TR_49 ;
	7'h4b :
		RG_rl_37_t1 = TR_49 ;
	7'h4c :
		RG_rl_37_t1 = TR_49 ;
	7'h4d :
		RG_rl_37_t1 = TR_49 ;
	7'h4e :
		RG_rl_37_t1 = TR_49 ;
	7'h4f :
		RG_rl_37_t1 = TR_49 ;
	7'h50 :
		RG_rl_37_t1 = TR_49 ;
	7'h51 :
		RG_rl_37_t1 = TR_49 ;
	7'h52 :
		RG_rl_37_t1 = TR_49 ;
	7'h53 :
		RG_rl_37_t1 = TR_49 ;
	7'h54 :
		RG_rl_37_t1 = TR_49 ;
	7'h55 :
		RG_rl_37_t1 = TR_49 ;
	7'h56 :
		RG_rl_37_t1 = TR_49 ;
	7'h57 :
		RG_rl_37_t1 = TR_49 ;
	7'h58 :
		RG_rl_37_t1 = TR_49 ;
	7'h59 :
		RG_rl_37_t1 = TR_49 ;
	7'h5a :
		RG_rl_37_t1 = TR_49 ;
	7'h5b :
		RG_rl_37_t1 = TR_49 ;
	7'h5c :
		RG_rl_37_t1 = TR_49 ;
	7'h5d :
		RG_rl_37_t1 = TR_49 ;
	7'h5e :
		RG_rl_37_t1 = TR_49 ;
	7'h5f :
		RG_rl_37_t1 = TR_49 ;
	7'h60 :
		RG_rl_37_t1 = TR_49 ;
	7'h61 :
		RG_rl_37_t1 = TR_49 ;
	7'h62 :
		RG_rl_37_t1 = TR_49 ;
	7'h63 :
		RG_rl_37_t1 = TR_49 ;
	7'h64 :
		RG_rl_37_t1 = TR_49 ;
	7'h65 :
		RG_rl_37_t1 = TR_49 ;
	7'h66 :
		RG_rl_37_t1 = TR_49 ;
	7'h67 :
		RG_rl_37_t1 = TR_49 ;
	7'h68 :
		RG_rl_37_t1 = TR_49 ;
	7'h69 :
		RG_rl_37_t1 = TR_49 ;
	7'h6a :
		RG_rl_37_t1 = TR_49 ;
	7'h6b :
		RG_rl_37_t1 = TR_49 ;
	7'h6c :
		RG_rl_37_t1 = TR_49 ;
	7'h6d :
		RG_rl_37_t1 = TR_49 ;
	7'h6e :
		RG_rl_37_t1 = TR_49 ;
	7'h6f :
		RG_rl_37_t1 = TR_49 ;
	7'h70 :
		RG_rl_37_t1 = TR_49 ;
	7'h71 :
		RG_rl_37_t1 = TR_49 ;
	7'h72 :
		RG_rl_37_t1 = TR_49 ;
	7'h73 :
		RG_rl_37_t1 = TR_49 ;
	7'h74 :
		RG_rl_37_t1 = TR_49 ;
	7'h75 :
		RG_rl_37_t1 = TR_49 ;
	7'h76 :
		RG_rl_37_t1 = TR_49 ;
	7'h77 :
		RG_rl_37_t1 = TR_49 ;
	7'h78 :
		RG_rl_37_t1 = TR_49 ;
	7'h79 :
		RG_rl_37_t1 = TR_49 ;
	7'h7a :
		RG_rl_37_t1 = TR_49 ;
	7'h7b :
		RG_rl_37_t1 = TR_49 ;
	7'h7c :
		RG_rl_37_t1 = TR_49 ;
	7'h7d :
		RG_rl_37_t1 = TR_49 ;
	7'h7e :
		RG_rl_37_t1 = TR_49 ;
	7'h7f :
		RG_rl_37_t1 = TR_49 ;
	default :
		RG_rl_37_t1 = 9'hx ;
	endcase
always @ ( RG_rl_37_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_220 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_37_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h25 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_37_t = ( ( { 9{ U_570 } } & RG_rl_220 )
		| ( { 9{ U_569 } } & RG_rl_37_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_37_en = ( U_570 | RG_rl_37_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_37_en )
		RG_rl_37 <= RG_rl_37_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_50 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_38_t1 = TR_50 ;
	7'h01 :
		RG_rl_38_t1 = TR_50 ;
	7'h02 :
		RG_rl_38_t1 = TR_50 ;
	7'h03 :
		RG_rl_38_t1 = TR_50 ;
	7'h04 :
		RG_rl_38_t1 = TR_50 ;
	7'h05 :
		RG_rl_38_t1 = TR_50 ;
	7'h06 :
		RG_rl_38_t1 = TR_50 ;
	7'h07 :
		RG_rl_38_t1 = TR_50 ;
	7'h08 :
		RG_rl_38_t1 = TR_50 ;
	7'h09 :
		RG_rl_38_t1 = TR_50 ;
	7'h0a :
		RG_rl_38_t1 = TR_50 ;
	7'h0b :
		RG_rl_38_t1 = TR_50 ;
	7'h0c :
		RG_rl_38_t1 = TR_50 ;
	7'h0d :
		RG_rl_38_t1 = TR_50 ;
	7'h0e :
		RG_rl_38_t1 = TR_50 ;
	7'h0f :
		RG_rl_38_t1 = TR_50 ;
	7'h10 :
		RG_rl_38_t1 = TR_50 ;
	7'h11 :
		RG_rl_38_t1 = TR_50 ;
	7'h12 :
		RG_rl_38_t1 = TR_50 ;
	7'h13 :
		RG_rl_38_t1 = TR_50 ;
	7'h14 :
		RG_rl_38_t1 = TR_50 ;
	7'h15 :
		RG_rl_38_t1 = TR_50 ;
	7'h16 :
		RG_rl_38_t1 = TR_50 ;
	7'h17 :
		RG_rl_38_t1 = TR_50 ;
	7'h18 :
		RG_rl_38_t1 = TR_50 ;
	7'h19 :
		RG_rl_38_t1 = TR_50 ;
	7'h1a :
		RG_rl_38_t1 = TR_50 ;
	7'h1b :
		RG_rl_38_t1 = TR_50 ;
	7'h1c :
		RG_rl_38_t1 = TR_50 ;
	7'h1d :
		RG_rl_38_t1 = TR_50 ;
	7'h1e :
		RG_rl_38_t1 = TR_50 ;
	7'h1f :
		RG_rl_38_t1 = TR_50 ;
	7'h20 :
		RG_rl_38_t1 = TR_50 ;
	7'h21 :
		RG_rl_38_t1 = TR_50 ;
	7'h22 :
		RG_rl_38_t1 = TR_50 ;
	7'h23 :
		RG_rl_38_t1 = TR_50 ;
	7'h24 :
		RG_rl_38_t1 = TR_50 ;
	7'h25 :
		RG_rl_38_t1 = TR_50 ;
	7'h26 :
		RG_rl_38_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h27 :
		RG_rl_38_t1 = TR_50 ;
	7'h28 :
		RG_rl_38_t1 = TR_50 ;
	7'h29 :
		RG_rl_38_t1 = TR_50 ;
	7'h2a :
		RG_rl_38_t1 = TR_50 ;
	7'h2b :
		RG_rl_38_t1 = TR_50 ;
	7'h2c :
		RG_rl_38_t1 = TR_50 ;
	7'h2d :
		RG_rl_38_t1 = TR_50 ;
	7'h2e :
		RG_rl_38_t1 = TR_50 ;
	7'h2f :
		RG_rl_38_t1 = TR_50 ;
	7'h30 :
		RG_rl_38_t1 = TR_50 ;
	7'h31 :
		RG_rl_38_t1 = TR_50 ;
	7'h32 :
		RG_rl_38_t1 = TR_50 ;
	7'h33 :
		RG_rl_38_t1 = TR_50 ;
	7'h34 :
		RG_rl_38_t1 = TR_50 ;
	7'h35 :
		RG_rl_38_t1 = TR_50 ;
	7'h36 :
		RG_rl_38_t1 = TR_50 ;
	7'h37 :
		RG_rl_38_t1 = TR_50 ;
	7'h38 :
		RG_rl_38_t1 = TR_50 ;
	7'h39 :
		RG_rl_38_t1 = TR_50 ;
	7'h3a :
		RG_rl_38_t1 = TR_50 ;
	7'h3b :
		RG_rl_38_t1 = TR_50 ;
	7'h3c :
		RG_rl_38_t1 = TR_50 ;
	7'h3d :
		RG_rl_38_t1 = TR_50 ;
	7'h3e :
		RG_rl_38_t1 = TR_50 ;
	7'h3f :
		RG_rl_38_t1 = TR_50 ;
	7'h40 :
		RG_rl_38_t1 = TR_50 ;
	7'h41 :
		RG_rl_38_t1 = TR_50 ;
	7'h42 :
		RG_rl_38_t1 = TR_50 ;
	7'h43 :
		RG_rl_38_t1 = TR_50 ;
	7'h44 :
		RG_rl_38_t1 = TR_50 ;
	7'h45 :
		RG_rl_38_t1 = TR_50 ;
	7'h46 :
		RG_rl_38_t1 = TR_50 ;
	7'h47 :
		RG_rl_38_t1 = TR_50 ;
	7'h48 :
		RG_rl_38_t1 = TR_50 ;
	7'h49 :
		RG_rl_38_t1 = TR_50 ;
	7'h4a :
		RG_rl_38_t1 = TR_50 ;
	7'h4b :
		RG_rl_38_t1 = TR_50 ;
	7'h4c :
		RG_rl_38_t1 = TR_50 ;
	7'h4d :
		RG_rl_38_t1 = TR_50 ;
	7'h4e :
		RG_rl_38_t1 = TR_50 ;
	7'h4f :
		RG_rl_38_t1 = TR_50 ;
	7'h50 :
		RG_rl_38_t1 = TR_50 ;
	7'h51 :
		RG_rl_38_t1 = TR_50 ;
	7'h52 :
		RG_rl_38_t1 = TR_50 ;
	7'h53 :
		RG_rl_38_t1 = TR_50 ;
	7'h54 :
		RG_rl_38_t1 = TR_50 ;
	7'h55 :
		RG_rl_38_t1 = TR_50 ;
	7'h56 :
		RG_rl_38_t1 = TR_50 ;
	7'h57 :
		RG_rl_38_t1 = TR_50 ;
	7'h58 :
		RG_rl_38_t1 = TR_50 ;
	7'h59 :
		RG_rl_38_t1 = TR_50 ;
	7'h5a :
		RG_rl_38_t1 = TR_50 ;
	7'h5b :
		RG_rl_38_t1 = TR_50 ;
	7'h5c :
		RG_rl_38_t1 = TR_50 ;
	7'h5d :
		RG_rl_38_t1 = TR_50 ;
	7'h5e :
		RG_rl_38_t1 = TR_50 ;
	7'h5f :
		RG_rl_38_t1 = TR_50 ;
	7'h60 :
		RG_rl_38_t1 = TR_50 ;
	7'h61 :
		RG_rl_38_t1 = TR_50 ;
	7'h62 :
		RG_rl_38_t1 = TR_50 ;
	7'h63 :
		RG_rl_38_t1 = TR_50 ;
	7'h64 :
		RG_rl_38_t1 = TR_50 ;
	7'h65 :
		RG_rl_38_t1 = TR_50 ;
	7'h66 :
		RG_rl_38_t1 = TR_50 ;
	7'h67 :
		RG_rl_38_t1 = TR_50 ;
	7'h68 :
		RG_rl_38_t1 = TR_50 ;
	7'h69 :
		RG_rl_38_t1 = TR_50 ;
	7'h6a :
		RG_rl_38_t1 = TR_50 ;
	7'h6b :
		RG_rl_38_t1 = TR_50 ;
	7'h6c :
		RG_rl_38_t1 = TR_50 ;
	7'h6d :
		RG_rl_38_t1 = TR_50 ;
	7'h6e :
		RG_rl_38_t1 = TR_50 ;
	7'h6f :
		RG_rl_38_t1 = TR_50 ;
	7'h70 :
		RG_rl_38_t1 = TR_50 ;
	7'h71 :
		RG_rl_38_t1 = TR_50 ;
	7'h72 :
		RG_rl_38_t1 = TR_50 ;
	7'h73 :
		RG_rl_38_t1 = TR_50 ;
	7'h74 :
		RG_rl_38_t1 = TR_50 ;
	7'h75 :
		RG_rl_38_t1 = TR_50 ;
	7'h76 :
		RG_rl_38_t1 = TR_50 ;
	7'h77 :
		RG_rl_38_t1 = TR_50 ;
	7'h78 :
		RG_rl_38_t1 = TR_50 ;
	7'h79 :
		RG_rl_38_t1 = TR_50 ;
	7'h7a :
		RG_rl_38_t1 = TR_50 ;
	7'h7b :
		RG_rl_38_t1 = TR_50 ;
	7'h7c :
		RG_rl_38_t1 = TR_50 ;
	7'h7d :
		RG_rl_38_t1 = TR_50 ;
	7'h7e :
		RG_rl_38_t1 = TR_50 ;
	7'h7f :
		RG_rl_38_t1 = TR_50 ;
	default :
		RG_rl_38_t1 = 9'hx ;
	endcase
always @ ( RG_rl_38_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_221 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_38_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h26 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_38_t = ( ( { 9{ U_570 } } & RG_rl_221 )
		| ( { 9{ U_569 } } & RG_rl_38_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_38_en = ( U_570 | RG_rl_38_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_38_en )
		RG_rl_38 <= RG_rl_38_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_51 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_39_t1 = TR_51 ;
	7'h01 :
		RG_rl_39_t1 = TR_51 ;
	7'h02 :
		RG_rl_39_t1 = TR_51 ;
	7'h03 :
		RG_rl_39_t1 = TR_51 ;
	7'h04 :
		RG_rl_39_t1 = TR_51 ;
	7'h05 :
		RG_rl_39_t1 = TR_51 ;
	7'h06 :
		RG_rl_39_t1 = TR_51 ;
	7'h07 :
		RG_rl_39_t1 = TR_51 ;
	7'h08 :
		RG_rl_39_t1 = TR_51 ;
	7'h09 :
		RG_rl_39_t1 = TR_51 ;
	7'h0a :
		RG_rl_39_t1 = TR_51 ;
	7'h0b :
		RG_rl_39_t1 = TR_51 ;
	7'h0c :
		RG_rl_39_t1 = TR_51 ;
	7'h0d :
		RG_rl_39_t1 = TR_51 ;
	7'h0e :
		RG_rl_39_t1 = TR_51 ;
	7'h0f :
		RG_rl_39_t1 = TR_51 ;
	7'h10 :
		RG_rl_39_t1 = TR_51 ;
	7'h11 :
		RG_rl_39_t1 = TR_51 ;
	7'h12 :
		RG_rl_39_t1 = TR_51 ;
	7'h13 :
		RG_rl_39_t1 = TR_51 ;
	7'h14 :
		RG_rl_39_t1 = TR_51 ;
	7'h15 :
		RG_rl_39_t1 = TR_51 ;
	7'h16 :
		RG_rl_39_t1 = TR_51 ;
	7'h17 :
		RG_rl_39_t1 = TR_51 ;
	7'h18 :
		RG_rl_39_t1 = TR_51 ;
	7'h19 :
		RG_rl_39_t1 = TR_51 ;
	7'h1a :
		RG_rl_39_t1 = TR_51 ;
	7'h1b :
		RG_rl_39_t1 = TR_51 ;
	7'h1c :
		RG_rl_39_t1 = TR_51 ;
	7'h1d :
		RG_rl_39_t1 = TR_51 ;
	7'h1e :
		RG_rl_39_t1 = TR_51 ;
	7'h1f :
		RG_rl_39_t1 = TR_51 ;
	7'h20 :
		RG_rl_39_t1 = TR_51 ;
	7'h21 :
		RG_rl_39_t1 = TR_51 ;
	7'h22 :
		RG_rl_39_t1 = TR_51 ;
	7'h23 :
		RG_rl_39_t1 = TR_51 ;
	7'h24 :
		RG_rl_39_t1 = TR_51 ;
	7'h25 :
		RG_rl_39_t1 = TR_51 ;
	7'h26 :
		RG_rl_39_t1 = TR_51 ;
	7'h27 :
		RG_rl_39_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h28 :
		RG_rl_39_t1 = TR_51 ;
	7'h29 :
		RG_rl_39_t1 = TR_51 ;
	7'h2a :
		RG_rl_39_t1 = TR_51 ;
	7'h2b :
		RG_rl_39_t1 = TR_51 ;
	7'h2c :
		RG_rl_39_t1 = TR_51 ;
	7'h2d :
		RG_rl_39_t1 = TR_51 ;
	7'h2e :
		RG_rl_39_t1 = TR_51 ;
	7'h2f :
		RG_rl_39_t1 = TR_51 ;
	7'h30 :
		RG_rl_39_t1 = TR_51 ;
	7'h31 :
		RG_rl_39_t1 = TR_51 ;
	7'h32 :
		RG_rl_39_t1 = TR_51 ;
	7'h33 :
		RG_rl_39_t1 = TR_51 ;
	7'h34 :
		RG_rl_39_t1 = TR_51 ;
	7'h35 :
		RG_rl_39_t1 = TR_51 ;
	7'h36 :
		RG_rl_39_t1 = TR_51 ;
	7'h37 :
		RG_rl_39_t1 = TR_51 ;
	7'h38 :
		RG_rl_39_t1 = TR_51 ;
	7'h39 :
		RG_rl_39_t1 = TR_51 ;
	7'h3a :
		RG_rl_39_t1 = TR_51 ;
	7'h3b :
		RG_rl_39_t1 = TR_51 ;
	7'h3c :
		RG_rl_39_t1 = TR_51 ;
	7'h3d :
		RG_rl_39_t1 = TR_51 ;
	7'h3e :
		RG_rl_39_t1 = TR_51 ;
	7'h3f :
		RG_rl_39_t1 = TR_51 ;
	7'h40 :
		RG_rl_39_t1 = TR_51 ;
	7'h41 :
		RG_rl_39_t1 = TR_51 ;
	7'h42 :
		RG_rl_39_t1 = TR_51 ;
	7'h43 :
		RG_rl_39_t1 = TR_51 ;
	7'h44 :
		RG_rl_39_t1 = TR_51 ;
	7'h45 :
		RG_rl_39_t1 = TR_51 ;
	7'h46 :
		RG_rl_39_t1 = TR_51 ;
	7'h47 :
		RG_rl_39_t1 = TR_51 ;
	7'h48 :
		RG_rl_39_t1 = TR_51 ;
	7'h49 :
		RG_rl_39_t1 = TR_51 ;
	7'h4a :
		RG_rl_39_t1 = TR_51 ;
	7'h4b :
		RG_rl_39_t1 = TR_51 ;
	7'h4c :
		RG_rl_39_t1 = TR_51 ;
	7'h4d :
		RG_rl_39_t1 = TR_51 ;
	7'h4e :
		RG_rl_39_t1 = TR_51 ;
	7'h4f :
		RG_rl_39_t1 = TR_51 ;
	7'h50 :
		RG_rl_39_t1 = TR_51 ;
	7'h51 :
		RG_rl_39_t1 = TR_51 ;
	7'h52 :
		RG_rl_39_t1 = TR_51 ;
	7'h53 :
		RG_rl_39_t1 = TR_51 ;
	7'h54 :
		RG_rl_39_t1 = TR_51 ;
	7'h55 :
		RG_rl_39_t1 = TR_51 ;
	7'h56 :
		RG_rl_39_t1 = TR_51 ;
	7'h57 :
		RG_rl_39_t1 = TR_51 ;
	7'h58 :
		RG_rl_39_t1 = TR_51 ;
	7'h59 :
		RG_rl_39_t1 = TR_51 ;
	7'h5a :
		RG_rl_39_t1 = TR_51 ;
	7'h5b :
		RG_rl_39_t1 = TR_51 ;
	7'h5c :
		RG_rl_39_t1 = TR_51 ;
	7'h5d :
		RG_rl_39_t1 = TR_51 ;
	7'h5e :
		RG_rl_39_t1 = TR_51 ;
	7'h5f :
		RG_rl_39_t1 = TR_51 ;
	7'h60 :
		RG_rl_39_t1 = TR_51 ;
	7'h61 :
		RG_rl_39_t1 = TR_51 ;
	7'h62 :
		RG_rl_39_t1 = TR_51 ;
	7'h63 :
		RG_rl_39_t1 = TR_51 ;
	7'h64 :
		RG_rl_39_t1 = TR_51 ;
	7'h65 :
		RG_rl_39_t1 = TR_51 ;
	7'h66 :
		RG_rl_39_t1 = TR_51 ;
	7'h67 :
		RG_rl_39_t1 = TR_51 ;
	7'h68 :
		RG_rl_39_t1 = TR_51 ;
	7'h69 :
		RG_rl_39_t1 = TR_51 ;
	7'h6a :
		RG_rl_39_t1 = TR_51 ;
	7'h6b :
		RG_rl_39_t1 = TR_51 ;
	7'h6c :
		RG_rl_39_t1 = TR_51 ;
	7'h6d :
		RG_rl_39_t1 = TR_51 ;
	7'h6e :
		RG_rl_39_t1 = TR_51 ;
	7'h6f :
		RG_rl_39_t1 = TR_51 ;
	7'h70 :
		RG_rl_39_t1 = TR_51 ;
	7'h71 :
		RG_rl_39_t1 = TR_51 ;
	7'h72 :
		RG_rl_39_t1 = TR_51 ;
	7'h73 :
		RG_rl_39_t1 = TR_51 ;
	7'h74 :
		RG_rl_39_t1 = TR_51 ;
	7'h75 :
		RG_rl_39_t1 = TR_51 ;
	7'h76 :
		RG_rl_39_t1 = TR_51 ;
	7'h77 :
		RG_rl_39_t1 = TR_51 ;
	7'h78 :
		RG_rl_39_t1 = TR_51 ;
	7'h79 :
		RG_rl_39_t1 = TR_51 ;
	7'h7a :
		RG_rl_39_t1 = TR_51 ;
	7'h7b :
		RG_rl_39_t1 = TR_51 ;
	7'h7c :
		RG_rl_39_t1 = TR_51 ;
	7'h7d :
		RG_rl_39_t1 = TR_51 ;
	7'h7e :
		RG_rl_39_t1 = TR_51 ;
	7'h7f :
		RG_rl_39_t1 = TR_51 ;
	default :
		RG_rl_39_t1 = 9'hx ;
	endcase
always @ ( RG_rl_39_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_222 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_39_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h27 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_39_t = ( ( { 9{ U_570 } } & RG_rl_222 )
		| ( { 9{ U_569 } } & RG_rl_39_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_39_en = ( U_570 | RG_rl_39_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_39_en )
		RG_rl_39 <= RG_rl_39_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_52 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_40_t1 = TR_52 ;
	7'h01 :
		RG_rl_40_t1 = TR_52 ;
	7'h02 :
		RG_rl_40_t1 = TR_52 ;
	7'h03 :
		RG_rl_40_t1 = TR_52 ;
	7'h04 :
		RG_rl_40_t1 = TR_52 ;
	7'h05 :
		RG_rl_40_t1 = TR_52 ;
	7'h06 :
		RG_rl_40_t1 = TR_52 ;
	7'h07 :
		RG_rl_40_t1 = TR_52 ;
	7'h08 :
		RG_rl_40_t1 = TR_52 ;
	7'h09 :
		RG_rl_40_t1 = TR_52 ;
	7'h0a :
		RG_rl_40_t1 = TR_52 ;
	7'h0b :
		RG_rl_40_t1 = TR_52 ;
	7'h0c :
		RG_rl_40_t1 = TR_52 ;
	7'h0d :
		RG_rl_40_t1 = TR_52 ;
	7'h0e :
		RG_rl_40_t1 = TR_52 ;
	7'h0f :
		RG_rl_40_t1 = TR_52 ;
	7'h10 :
		RG_rl_40_t1 = TR_52 ;
	7'h11 :
		RG_rl_40_t1 = TR_52 ;
	7'h12 :
		RG_rl_40_t1 = TR_52 ;
	7'h13 :
		RG_rl_40_t1 = TR_52 ;
	7'h14 :
		RG_rl_40_t1 = TR_52 ;
	7'h15 :
		RG_rl_40_t1 = TR_52 ;
	7'h16 :
		RG_rl_40_t1 = TR_52 ;
	7'h17 :
		RG_rl_40_t1 = TR_52 ;
	7'h18 :
		RG_rl_40_t1 = TR_52 ;
	7'h19 :
		RG_rl_40_t1 = TR_52 ;
	7'h1a :
		RG_rl_40_t1 = TR_52 ;
	7'h1b :
		RG_rl_40_t1 = TR_52 ;
	7'h1c :
		RG_rl_40_t1 = TR_52 ;
	7'h1d :
		RG_rl_40_t1 = TR_52 ;
	7'h1e :
		RG_rl_40_t1 = TR_52 ;
	7'h1f :
		RG_rl_40_t1 = TR_52 ;
	7'h20 :
		RG_rl_40_t1 = TR_52 ;
	7'h21 :
		RG_rl_40_t1 = TR_52 ;
	7'h22 :
		RG_rl_40_t1 = TR_52 ;
	7'h23 :
		RG_rl_40_t1 = TR_52 ;
	7'h24 :
		RG_rl_40_t1 = TR_52 ;
	7'h25 :
		RG_rl_40_t1 = TR_52 ;
	7'h26 :
		RG_rl_40_t1 = TR_52 ;
	7'h27 :
		RG_rl_40_t1 = TR_52 ;
	7'h28 :
		RG_rl_40_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h29 :
		RG_rl_40_t1 = TR_52 ;
	7'h2a :
		RG_rl_40_t1 = TR_52 ;
	7'h2b :
		RG_rl_40_t1 = TR_52 ;
	7'h2c :
		RG_rl_40_t1 = TR_52 ;
	7'h2d :
		RG_rl_40_t1 = TR_52 ;
	7'h2e :
		RG_rl_40_t1 = TR_52 ;
	7'h2f :
		RG_rl_40_t1 = TR_52 ;
	7'h30 :
		RG_rl_40_t1 = TR_52 ;
	7'h31 :
		RG_rl_40_t1 = TR_52 ;
	7'h32 :
		RG_rl_40_t1 = TR_52 ;
	7'h33 :
		RG_rl_40_t1 = TR_52 ;
	7'h34 :
		RG_rl_40_t1 = TR_52 ;
	7'h35 :
		RG_rl_40_t1 = TR_52 ;
	7'h36 :
		RG_rl_40_t1 = TR_52 ;
	7'h37 :
		RG_rl_40_t1 = TR_52 ;
	7'h38 :
		RG_rl_40_t1 = TR_52 ;
	7'h39 :
		RG_rl_40_t1 = TR_52 ;
	7'h3a :
		RG_rl_40_t1 = TR_52 ;
	7'h3b :
		RG_rl_40_t1 = TR_52 ;
	7'h3c :
		RG_rl_40_t1 = TR_52 ;
	7'h3d :
		RG_rl_40_t1 = TR_52 ;
	7'h3e :
		RG_rl_40_t1 = TR_52 ;
	7'h3f :
		RG_rl_40_t1 = TR_52 ;
	7'h40 :
		RG_rl_40_t1 = TR_52 ;
	7'h41 :
		RG_rl_40_t1 = TR_52 ;
	7'h42 :
		RG_rl_40_t1 = TR_52 ;
	7'h43 :
		RG_rl_40_t1 = TR_52 ;
	7'h44 :
		RG_rl_40_t1 = TR_52 ;
	7'h45 :
		RG_rl_40_t1 = TR_52 ;
	7'h46 :
		RG_rl_40_t1 = TR_52 ;
	7'h47 :
		RG_rl_40_t1 = TR_52 ;
	7'h48 :
		RG_rl_40_t1 = TR_52 ;
	7'h49 :
		RG_rl_40_t1 = TR_52 ;
	7'h4a :
		RG_rl_40_t1 = TR_52 ;
	7'h4b :
		RG_rl_40_t1 = TR_52 ;
	7'h4c :
		RG_rl_40_t1 = TR_52 ;
	7'h4d :
		RG_rl_40_t1 = TR_52 ;
	7'h4e :
		RG_rl_40_t1 = TR_52 ;
	7'h4f :
		RG_rl_40_t1 = TR_52 ;
	7'h50 :
		RG_rl_40_t1 = TR_52 ;
	7'h51 :
		RG_rl_40_t1 = TR_52 ;
	7'h52 :
		RG_rl_40_t1 = TR_52 ;
	7'h53 :
		RG_rl_40_t1 = TR_52 ;
	7'h54 :
		RG_rl_40_t1 = TR_52 ;
	7'h55 :
		RG_rl_40_t1 = TR_52 ;
	7'h56 :
		RG_rl_40_t1 = TR_52 ;
	7'h57 :
		RG_rl_40_t1 = TR_52 ;
	7'h58 :
		RG_rl_40_t1 = TR_52 ;
	7'h59 :
		RG_rl_40_t1 = TR_52 ;
	7'h5a :
		RG_rl_40_t1 = TR_52 ;
	7'h5b :
		RG_rl_40_t1 = TR_52 ;
	7'h5c :
		RG_rl_40_t1 = TR_52 ;
	7'h5d :
		RG_rl_40_t1 = TR_52 ;
	7'h5e :
		RG_rl_40_t1 = TR_52 ;
	7'h5f :
		RG_rl_40_t1 = TR_52 ;
	7'h60 :
		RG_rl_40_t1 = TR_52 ;
	7'h61 :
		RG_rl_40_t1 = TR_52 ;
	7'h62 :
		RG_rl_40_t1 = TR_52 ;
	7'h63 :
		RG_rl_40_t1 = TR_52 ;
	7'h64 :
		RG_rl_40_t1 = TR_52 ;
	7'h65 :
		RG_rl_40_t1 = TR_52 ;
	7'h66 :
		RG_rl_40_t1 = TR_52 ;
	7'h67 :
		RG_rl_40_t1 = TR_52 ;
	7'h68 :
		RG_rl_40_t1 = TR_52 ;
	7'h69 :
		RG_rl_40_t1 = TR_52 ;
	7'h6a :
		RG_rl_40_t1 = TR_52 ;
	7'h6b :
		RG_rl_40_t1 = TR_52 ;
	7'h6c :
		RG_rl_40_t1 = TR_52 ;
	7'h6d :
		RG_rl_40_t1 = TR_52 ;
	7'h6e :
		RG_rl_40_t1 = TR_52 ;
	7'h6f :
		RG_rl_40_t1 = TR_52 ;
	7'h70 :
		RG_rl_40_t1 = TR_52 ;
	7'h71 :
		RG_rl_40_t1 = TR_52 ;
	7'h72 :
		RG_rl_40_t1 = TR_52 ;
	7'h73 :
		RG_rl_40_t1 = TR_52 ;
	7'h74 :
		RG_rl_40_t1 = TR_52 ;
	7'h75 :
		RG_rl_40_t1 = TR_52 ;
	7'h76 :
		RG_rl_40_t1 = TR_52 ;
	7'h77 :
		RG_rl_40_t1 = TR_52 ;
	7'h78 :
		RG_rl_40_t1 = TR_52 ;
	7'h79 :
		RG_rl_40_t1 = TR_52 ;
	7'h7a :
		RG_rl_40_t1 = TR_52 ;
	7'h7b :
		RG_rl_40_t1 = TR_52 ;
	7'h7c :
		RG_rl_40_t1 = TR_52 ;
	7'h7d :
		RG_rl_40_t1 = TR_52 ;
	7'h7e :
		RG_rl_40_t1 = TR_52 ;
	7'h7f :
		RG_rl_40_t1 = TR_52 ;
	default :
		RG_rl_40_t1 = 9'hx ;
	endcase
always @ ( RG_rl_40_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_223 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_40_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h28 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_40_t = ( ( { 9{ U_570 } } & RG_rl_223 )
		| ( { 9{ U_569 } } & RG_rl_40_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_40_en = ( U_570 | RG_rl_40_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_40_en )
		RG_rl_40 <= RG_rl_40_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_53 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_41_t1 = TR_53 ;
	7'h01 :
		RG_rl_41_t1 = TR_53 ;
	7'h02 :
		RG_rl_41_t1 = TR_53 ;
	7'h03 :
		RG_rl_41_t1 = TR_53 ;
	7'h04 :
		RG_rl_41_t1 = TR_53 ;
	7'h05 :
		RG_rl_41_t1 = TR_53 ;
	7'h06 :
		RG_rl_41_t1 = TR_53 ;
	7'h07 :
		RG_rl_41_t1 = TR_53 ;
	7'h08 :
		RG_rl_41_t1 = TR_53 ;
	7'h09 :
		RG_rl_41_t1 = TR_53 ;
	7'h0a :
		RG_rl_41_t1 = TR_53 ;
	7'h0b :
		RG_rl_41_t1 = TR_53 ;
	7'h0c :
		RG_rl_41_t1 = TR_53 ;
	7'h0d :
		RG_rl_41_t1 = TR_53 ;
	7'h0e :
		RG_rl_41_t1 = TR_53 ;
	7'h0f :
		RG_rl_41_t1 = TR_53 ;
	7'h10 :
		RG_rl_41_t1 = TR_53 ;
	7'h11 :
		RG_rl_41_t1 = TR_53 ;
	7'h12 :
		RG_rl_41_t1 = TR_53 ;
	7'h13 :
		RG_rl_41_t1 = TR_53 ;
	7'h14 :
		RG_rl_41_t1 = TR_53 ;
	7'h15 :
		RG_rl_41_t1 = TR_53 ;
	7'h16 :
		RG_rl_41_t1 = TR_53 ;
	7'h17 :
		RG_rl_41_t1 = TR_53 ;
	7'h18 :
		RG_rl_41_t1 = TR_53 ;
	7'h19 :
		RG_rl_41_t1 = TR_53 ;
	7'h1a :
		RG_rl_41_t1 = TR_53 ;
	7'h1b :
		RG_rl_41_t1 = TR_53 ;
	7'h1c :
		RG_rl_41_t1 = TR_53 ;
	7'h1d :
		RG_rl_41_t1 = TR_53 ;
	7'h1e :
		RG_rl_41_t1 = TR_53 ;
	7'h1f :
		RG_rl_41_t1 = TR_53 ;
	7'h20 :
		RG_rl_41_t1 = TR_53 ;
	7'h21 :
		RG_rl_41_t1 = TR_53 ;
	7'h22 :
		RG_rl_41_t1 = TR_53 ;
	7'h23 :
		RG_rl_41_t1 = TR_53 ;
	7'h24 :
		RG_rl_41_t1 = TR_53 ;
	7'h25 :
		RG_rl_41_t1 = TR_53 ;
	7'h26 :
		RG_rl_41_t1 = TR_53 ;
	7'h27 :
		RG_rl_41_t1 = TR_53 ;
	7'h28 :
		RG_rl_41_t1 = TR_53 ;
	7'h29 :
		RG_rl_41_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2a :
		RG_rl_41_t1 = TR_53 ;
	7'h2b :
		RG_rl_41_t1 = TR_53 ;
	7'h2c :
		RG_rl_41_t1 = TR_53 ;
	7'h2d :
		RG_rl_41_t1 = TR_53 ;
	7'h2e :
		RG_rl_41_t1 = TR_53 ;
	7'h2f :
		RG_rl_41_t1 = TR_53 ;
	7'h30 :
		RG_rl_41_t1 = TR_53 ;
	7'h31 :
		RG_rl_41_t1 = TR_53 ;
	7'h32 :
		RG_rl_41_t1 = TR_53 ;
	7'h33 :
		RG_rl_41_t1 = TR_53 ;
	7'h34 :
		RG_rl_41_t1 = TR_53 ;
	7'h35 :
		RG_rl_41_t1 = TR_53 ;
	7'h36 :
		RG_rl_41_t1 = TR_53 ;
	7'h37 :
		RG_rl_41_t1 = TR_53 ;
	7'h38 :
		RG_rl_41_t1 = TR_53 ;
	7'h39 :
		RG_rl_41_t1 = TR_53 ;
	7'h3a :
		RG_rl_41_t1 = TR_53 ;
	7'h3b :
		RG_rl_41_t1 = TR_53 ;
	7'h3c :
		RG_rl_41_t1 = TR_53 ;
	7'h3d :
		RG_rl_41_t1 = TR_53 ;
	7'h3e :
		RG_rl_41_t1 = TR_53 ;
	7'h3f :
		RG_rl_41_t1 = TR_53 ;
	7'h40 :
		RG_rl_41_t1 = TR_53 ;
	7'h41 :
		RG_rl_41_t1 = TR_53 ;
	7'h42 :
		RG_rl_41_t1 = TR_53 ;
	7'h43 :
		RG_rl_41_t1 = TR_53 ;
	7'h44 :
		RG_rl_41_t1 = TR_53 ;
	7'h45 :
		RG_rl_41_t1 = TR_53 ;
	7'h46 :
		RG_rl_41_t1 = TR_53 ;
	7'h47 :
		RG_rl_41_t1 = TR_53 ;
	7'h48 :
		RG_rl_41_t1 = TR_53 ;
	7'h49 :
		RG_rl_41_t1 = TR_53 ;
	7'h4a :
		RG_rl_41_t1 = TR_53 ;
	7'h4b :
		RG_rl_41_t1 = TR_53 ;
	7'h4c :
		RG_rl_41_t1 = TR_53 ;
	7'h4d :
		RG_rl_41_t1 = TR_53 ;
	7'h4e :
		RG_rl_41_t1 = TR_53 ;
	7'h4f :
		RG_rl_41_t1 = TR_53 ;
	7'h50 :
		RG_rl_41_t1 = TR_53 ;
	7'h51 :
		RG_rl_41_t1 = TR_53 ;
	7'h52 :
		RG_rl_41_t1 = TR_53 ;
	7'h53 :
		RG_rl_41_t1 = TR_53 ;
	7'h54 :
		RG_rl_41_t1 = TR_53 ;
	7'h55 :
		RG_rl_41_t1 = TR_53 ;
	7'h56 :
		RG_rl_41_t1 = TR_53 ;
	7'h57 :
		RG_rl_41_t1 = TR_53 ;
	7'h58 :
		RG_rl_41_t1 = TR_53 ;
	7'h59 :
		RG_rl_41_t1 = TR_53 ;
	7'h5a :
		RG_rl_41_t1 = TR_53 ;
	7'h5b :
		RG_rl_41_t1 = TR_53 ;
	7'h5c :
		RG_rl_41_t1 = TR_53 ;
	7'h5d :
		RG_rl_41_t1 = TR_53 ;
	7'h5e :
		RG_rl_41_t1 = TR_53 ;
	7'h5f :
		RG_rl_41_t1 = TR_53 ;
	7'h60 :
		RG_rl_41_t1 = TR_53 ;
	7'h61 :
		RG_rl_41_t1 = TR_53 ;
	7'h62 :
		RG_rl_41_t1 = TR_53 ;
	7'h63 :
		RG_rl_41_t1 = TR_53 ;
	7'h64 :
		RG_rl_41_t1 = TR_53 ;
	7'h65 :
		RG_rl_41_t1 = TR_53 ;
	7'h66 :
		RG_rl_41_t1 = TR_53 ;
	7'h67 :
		RG_rl_41_t1 = TR_53 ;
	7'h68 :
		RG_rl_41_t1 = TR_53 ;
	7'h69 :
		RG_rl_41_t1 = TR_53 ;
	7'h6a :
		RG_rl_41_t1 = TR_53 ;
	7'h6b :
		RG_rl_41_t1 = TR_53 ;
	7'h6c :
		RG_rl_41_t1 = TR_53 ;
	7'h6d :
		RG_rl_41_t1 = TR_53 ;
	7'h6e :
		RG_rl_41_t1 = TR_53 ;
	7'h6f :
		RG_rl_41_t1 = TR_53 ;
	7'h70 :
		RG_rl_41_t1 = TR_53 ;
	7'h71 :
		RG_rl_41_t1 = TR_53 ;
	7'h72 :
		RG_rl_41_t1 = TR_53 ;
	7'h73 :
		RG_rl_41_t1 = TR_53 ;
	7'h74 :
		RG_rl_41_t1 = TR_53 ;
	7'h75 :
		RG_rl_41_t1 = TR_53 ;
	7'h76 :
		RG_rl_41_t1 = TR_53 ;
	7'h77 :
		RG_rl_41_t1 = TR_53 ;
	7'h78 :
		RG_rl_41_t1 = TR_53 ;
	7'h79 :
		RG_rl_41_t1 = TR_53 ;
	7'h7a :
		RG_rl_41_t1 = TR_53 ;
	7'h7b :
		RG_rl_41_t1 = TR_53 ;
	7'h7c :
		RG_rl_41_t1 = TR_53 ;
	7'h7d :
		RG_rl_41_t1 = TR_53 ;
	7'h7e :
		RG_rl_41_t1 = TR_53 ;
	7'h7f :
		RG_rl_41_t1 = TR_53 ;
	default :
		RG_rl_41_t1 = 9'hx ;
	endcase
always @ ( RG_rl_41_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_224 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_41_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h29 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_41_t = ( ( { 9{ U_570 } } & RG_rl_224 )
		| ( { 9{ U_569 } } & RG_rl_41_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_41_en = ( U_570 | RG_rl_41_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_41_en )
		RG_rl_41 <= RG_rl_41_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_54 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_42_t1 = TR_54 ;
	7'h01 :
		RG_rl_42_t1 = TR_54 ;
	7'h02 :
		RG_rl_42_t1 = TR_54 ;
	7'h03 :
		RG_rl_42_t1 = TR_54 ;
	7'h04 :
		RG_rl_42_t1 = TR_54 ;
	7'h05 :
		RG_rl_42_t1 = TR_54 ;
	7'h06 :
		RG_rl_42_t1 = TR_54 ;
	7'h07 :
		RG_rl_42_t1 = TR_54 ;
	7'h08 :
		RG_rl_42_t1 = TR_54 ;
	7'h09 :
		RG_rl_42_t1 = TR_54 ;
	7'h0a :
		RG_rl_42_t1 = TR_54 ;
	7'h0b :
		RG_rl_42_t1 = TR_54 ;
	7'h0c :
		RG_rl_42_t1 = TR_54 ;
	7'h0d :
		RG_rl_42_t1 = TR_54 ;
	7'h0e :
		RG_rl_42_t1 = TR_54 ;
	7'h0f :
		RG_rl_42_t1 = TR_54 ;
	7'h10 :
		RG_rl_42_t1 = TR_54 ;
	7'h11 :
		RG_rl_42_t1 = TR_54 ;
	7'h12 :
		RG_rl_42_t1 = TR_54 ;
	7'h13 :
		RG_rl_42_t1 = TR_54 ;
	7'h14 :
		RG_rl_42_t1 = TR_54 ;
	7'h15 :
		RG_rl_42_t1 = TR_54 ;
	7'h16 :
		RG_rl_42_t1 = TR_54 ;
	7'h17 :
		RG_rl_42_t1 = TR_54 ;
	7'h18 :
		RG_rl_42_t1 = TR_54 ;
	7'h19 :
		RG_rl_42_t1 = TR_54 ;
	7'h1a :
		RG_rl_42_t1 = TR_54 ;
	7'h1b :
		RG_rl_42_t1 = TR_54 ;
	7'h1c :
		RG_rl_42_t1 = TR_54 ;
	7'h1d :
		RG_rl_42_t1 = TR_54 ;
	7'h1e :
		RG_rl_42_t1 = TR_54 ;
	7'h1f :
		RG_rl_42_t1 = TR_54 ;
	7'h20 :
		RG_rl_42_t1 = TR_54 ;
	7'h21 :
		RG_rl_42_t1 = TR_54 ;
	7'h22 :
		RG_rl_42_t1 = TR_54 ;
	7'h23 :
		RG_rl_42_t1 = TR_54 ;
	7'h24 :
		RG_rl_42_t1 = TR_54 ;
	7'h25 :
		RG_rl_42_t1 = TR_54 ;
	7'h26 :
		RG_rl_42_t1 = TR_54 ;
	7'h27 :
		RG_rl_42_t1 = TR_54 ;
	7'h28 :
		RG_rl_42_t1 = TR_54 ;
	7'h29 :
		RG_rl_42_t1 = TR_54 ;
	7'h2a :
		RG_rl_42_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2b :
		RG_rl_42_t1 = TR_54 ;
	7'h2c :
		RG_rl_42_t1 = TR_54 ;
	7'h2d :
		RG_rl_42_t1 = TR_54 ;
	7'h2e :
		RG_rl_42_t1 = TR_54 ;
	7'h2f :
		RG_rl_42_t1 = TR_54 ;
	7'h30 :
		RG_rl_42_t1 = TR_54 ;
	7'h31 :
		RG_rl_42_t1 = TR_54 ;
	7'h32 :
		RG_rl_42_t1 = TR_54 ;
	7'h33 :
		RG_rl_42_t1 = TR_54 ;
	7'h34 :
		RG_rl_42_t1 = TR_54 ;
	7'h35 :
		RG_rl_42_t1 = TR_54 ;
	7'h36 :
		RG_rl_42_t1 = TR_54 ;
	7'h37 :
		RG_rl_42_t1 = TR_54 ;
	7'h38 :
		RG_rl_42_t1 = TR_54 ;
	7'h39 :
		RG_rl_42_t1 = TR_54 ;
	7'h3a :
		RG_rl_42_t1 = TR_54 ;
	7'h3b :
		RG_rl_42_t1 = TR_54 ;
	7'h3c :
		RG_rl_42_t1 = TR_54 ;
	7'h3d :
		RG_rl_42_t1 = TR_54 ;
	7'h3e :
		RG_rl_42_t1 = TR_54 ;
	7'h3f :
		RG_rl_42_t1 = TR_54 ;
	7'h40 :
		RG_rl_42_t1 = TR_54 ;
	7'h41 :
		RG_rl_42_t1 = TR_54 ;
	7'h42 :
		RG_rl_42_t1 = TR_54 ;
	7'h43 :
		RG_rl_42_t1 = TR_54 ;
	7'h44 :
		RG_rl_42_t1 = TR_54 ;
	7'h45 :
		RG_rl_42_t1 = TR_54 ;
	7'h46 :
		RG_rl_42_t1 = TR_54 ;
	7'h47 :
		RG_rl_42_t1 = TR_54 ;
	7'h48 :
		RG_rl_42_t1 = TR_54 ;
	7'h49 :
		RG_rl_42_t1 = TR_54 ;
	7'h4a :
		RG_rl_42_t1 = TR_54 ;
	7'h4b :
		RG_rl_42_t1 = TR_54 ;
	7'h4c :
		RG_rl_42_t1 = TR_54 ;
	7'h4d :
		RG_rl_42_t1 = TR_54 ;
	7'h4e :
		RG_rl_42_t1 = TR_54 ;
	7'h4f :
		RG_rl_42_t1 = TR_54 ;
	7'h50 :
		RG_rl_42_t1 = TR_54 ;
	7'h51 :
		RG_rl_42_t1 = TR_54 ;
	7'h52 :
		RG_rl_42_t1 = TR_54 ;
	7'h53 :
		RG_rl_42_t1 = TR_54 ;
	7'h54 :
		RG_rl_42_t1 = TR_54 ;
	7'h55 :
		RG_rl_42_t1 = TR_54 ;
	7'h56 :
		RG_rl_42_t1 = TR_54 ;
	7'h57 :
		RG_rl_42_t1 = TR_54 ;
	7'h58 :
		RG_rl_42_t1 = TR_54 ;
	7'h59 :
		RG_rl_42_t1 = TR_54 ;
	7'h5a :
		RG_rl_42_t1 = TR_54 ;
	7'h5b :
		RG_rl_42_t1 = TR_54 ;
	7'h5c :
		RG_rl_42_t1 = TR_54 ;
	7'h5d :
		RG_rl_42_t1 = TR_54 ;
	7'h5e :
		RG_rl_42_t1 = TR_54 ;
	7'h5f :
		RG_rl_42_t1 = TR_54 ;
	7'h60 :
		RG_rl_42_t1 = TR_54 ;
	7'h61 :
		RG_rl_42_t1 = TR_54 ;
	7'h62 :
		RG_rl_42_t1 = TR_54 ;
	7'h63 :
		RG_rl_42_t1 = TR_54 ;
	7'h64 :
		RG_rl_42_t1 = TR_54 ;
	7'h65 :
		RG_rl_42_t1 = TR_54 ;
	7'h66 :
		RG_rl_42_t1 = TR_54 ;
	7'h67 :
		RG_rl_42_t1 = TR_54 ;
	7'h68 :
		RG_rl_42_t1 = TR_54 ;
	7'h69 :
		RG_rl_42_t1 = TR_54 ;
	7'h6a :
		RG_rl_42_t1 = TR_54 ;
	7'h6b :
		RG_rl_42_t1 = TR_54 ;
	7'h6c :
		RG_rl_42_t1 = TR_54 ;
	7'h6d :
		RG_rl_42_t1 = TR_54 ;
	7'h6e :
		RG_rl_42_t1 = TR_54 ;
	7'h6f :
		RG_rl_42_t1 = TR_54 ;
	7'h70 :
		RG_rl_42_t1 = TR_54 ;
	7'h71 :
		RG_rl_42_t1 = TR_54 ;
	7'h72 :
		RG_rl_42_t1 = TR_54 ;
	7'h73 :
		RG_rl_42_t1 = TR_54 ;
	7'h74 :
		RG_rl_42_t1 = TR_54 ;
	7'h75 :
		RG_rl_42_t1 = TR_54 ;
	7'h76 :
		RG_rl_42_t1 = TR_54 ;
	7'h77 :
		RG_rl_42_t1 = TR_54 ;
	7'h78 :
		RG_rl_42_t1 = TR_54 ;
	7'h79 :
		RG_rl_42_t1 = TR_54 ;
	7'h7a :
		RG_rl_42_t1 = TR_54 ;
	7'h7b :
		RG_rl_42_t1 = TR_54 ;
	7'h7c :
		RG_rl_42_t1 = TR_54 ;
	7'h7d :
		RG_rl_42_t1 = TR_54 ;
	7'h7e :
		RG_rl_42_t1 = TR_54 ;
	7'h7f :
		RG_rl_42_t1 = TR_54 ;
	default :
		RG_rl_42_t1 = 9'hx ;
	endcase
always @ ( RG_rl_42_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_225 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_42_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h2a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_42_t = ( ( { 9{ U_570 } } & RG_rl_225 )
		| ( { 9{ U_569 } } & RG_rl_42_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_42_en = ( U_570 | RG_rl_42_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_42_en )
		RG_rl_42 <= RG_rl_42_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_55 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_43_t1 = TR_55 ;
	7'h01 :
		RG_rl_43_t1 = TR_55 ;
	7'h02 :
		RG_rl_43_t1 = TR_55 ;
	7'h03 :
		RG_rl_43_t1 = TR_55 ;
	7'h04 :
		RG_rl_43_t1 = TR_55 ;
	7'h05 :
		RG_rl_43_t1 = TR_55 ;
	7'h06 :
		RG_rl_43_t1 = TR_55 ;
	7'h07 :
		RG_rl_43_t1 = TR_55 ;
	7'h08 :
		RG_rl_43_t1 = TR_55 ;
	7'h09 :
		RG_rl_43_t1 = TR_55 ;
	7'h0a :
		RG_rl_43_t1 = TR_55 ;
	7'h0b :
		RG_rl_43_t1 = TR_55 ;
	7'h0c :
		RG_rl_43_t1 = TR_55 ;
	7'h0d :
		RG_rl_43_t1 = TR_55 ;
	7'h0e :
		RG_rl_43_t1 = TR_55 ;
	7'h0f :
		RG_rl_43_t1 = TR_55 ;
	7'h10 :
		RG_rl_43_t1 = TR_55 ;
	7'h11 :
		RG_rl_43_t1 = TR_55 ;
	7'h12 :
		RG_rl_43_t1 = TR_55 ;
	7'h13 :
		RG_rl_43_t1 = TR_55 ;
	7'h14 :
		RG_rl_43_t1 = TR_55 ;
	7'h15 :
		RG_rl_43_t1 = TR_55 ;
	7'h16 :
		RG_rl_43_t1 = TR_55 ;
	7'h17 :
		RG_rl_43_t1 = TR_55 ;
	7'h18 :
		RG_rl_43_t1 = TR_55 ;
	7'h19 :
		RG_rl_43_t1 = TR_55 ;
	7'h1a :
		RG_rl_43_t1 = TR_55 ;
	7'h1b :
		RG_rl_43_t1 = TR_55 ;
	7'h1c :
		RG_rl_43_t1 = TR_55 ;
	7'h1d :
		RG_rl_43_t1 = TR_55 ;
	7'h1e :
		RG_rl_43_t1 = TR_55 ;
	7'h1f :
		RG_rl_43_t1 = TR_55 ;
	7'h20 :
		RG_rl_43_t1 = TR_55 ;
	7'h21 :
		RG_rl_43_t1 = TR_55 ;
	7'h22 :
		RG_rl_43_t1 = TR_55 ;
	7'h23 :
		RG_rl_43_t1 = TR_55 ;
	7'h24 :
		RG_rl_43_t1 = TR_55 ;
	7'h25 :
		RG_rl_43_t1 = TR_55 ;
	7'h26 :
		RG_rl_43_t1 = TR_55 ;
	7'h27 :
		RG_rl_43_t1 = TR_55 ;
	7'h28 :
		RG_rl_43_t1 = TR_55 ;
	7'h29 :
		RG_rl_43_t1 = TR_55 ;
	7'h2a :
		RG_rl_43_t1 = TR_55 ;
	7'h2b :
		RG_rl_43_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2c :
		RG_rl_43_t1 = TR_55 ;
	7'h2d :
		RG_rl_43_t1 = TR_55 ;
	7'h2e :
		RG_rl_43_t1 = TR_55 ;
	7'h2f :
		RG_rl_43_t1 = TR_55 ;
	7'h30 :
		RG_rl_43_t1 = TR_55 ;
	7'h31 :
		RG_rl_43_t1 = TR_55 ;
	7'h32 :
		RG_rl_43_t1 = TR_55 ;
	7'h33 :
		RG_rl_43_t1 = TR_55 ;
	7'h34 :
		RG_rl_43_t1 = TR_55 ;
	7'h35 :
		RG_rl_43_t1 = TR_55 ;
	7'h36 :
		RG_rl_43_t1 = TR_55 ;
	7'h37 :
		RG_rl_43_t1 = TR_55 ;
	7'h38 :
		RG_rl_43_t1 = TR_55 ;
	7'h39 :
		RG_rl_43_t1 = TR_55 ;
	7'h3a :
		RG_rl_43_t1 = TR_55 ;
	7'h3b :
		RG_rl_43_t1 = TR_55 ;
	7'h3c :
		RG_rl_43_t1 = TR_55 ;
	7'h3d :
		RG_rl_43_t1 = TR_55 ;
	7'h3e :
		RG_rl_43_t1 = TR_55 ;
	7'h3f :
		RG_rl_43_t1 = TR_55 ;
	7'h40 :
		RG_rl_43_t1 = TR_55 ;
	7'h41 :
		RG_rl_43_t1 = TR_55 ;
	7'h42 :
		RG_rl_43_t1 = TR_55 ;
	7'h43 :
		RG_rl_43_t1 = TR_55 ;
	7'h44 :
		RG_rl_43_t1 = TR_55 ;
	7'h45 :
		RG_rl_43_t1 = TR_55 ;
	7'h46 :
		RG_rl_43_t1 = TR_55 ;
	7'h47 :
		RG_rl_43_t1 = TR_55 ;
	7'h48 :
		RG_rl_43_t1 = TR_55 ;
	7'h49 :
		RG_rl_43_t1 = TR_55 ;
	7'h4a :
		RG_rl_43_t1 = TR_55 ;
	7'h4b :
		RG_rl_43_t1 = TR_55 ;
	7'h4c :
		RG_rl_43_t1 = TR_55 ;
	7'h4d :
		RG_rl_43_t1 = TR_55 ;
	7'h4e :
		RG_rl_43_t1 = TR_55 ;
	7'h4f :
		RG_rl_43_t1 = TR_55 ;
	7'h50 :
		RG_rl_43_t1 = TR_55 ;
	7'h51 :
		RG_rl_43_t1 = TR_55 ;
	7'h52 :
		RG_rl_43_t1 = TR_55 ;
	7'h53 :
		RG_rl_43_t1 = TR_55 ;
	7'h54 :
		RG_rl_43_t1 = TR_55 ;
	7'h55 :
		RG_rl_43_t1 = TR_55 ;
	7'h56 :
		RG_rl_43_t1 = TR_55 ;
	7'h57 :
		RG_rl_43_t1 = TR_55 ;
	7'h58 :
		RG_rl_43_t1 = TR_55 ;
	7'h59 :
		RG_rl_43_t1 = TR_55 ;
	7'h5a :
		RG_rl_43_t1 = TR_55 ;
	7'h5b :
		RG_rl_43_t1 = TR_55 ;
	7'h5c :
		RG_rl_43_t1 = TR_55 ;
	7'h5d :
		RG_rl_43_t1 = TR_55 ;
	7'h5e :
		RG_rl_43_t1 = TR_55 ;
	7'h5f :
		RG_rl_43_t1 = TR_55 ;
	7'h60 :
		RG_rl_43_t1 = TR_55 ;
	7'h61 :
		RG_rl_43_t1 = TR_55 ;
	7'h62 :
		RG_rl_43_t1 = TR_55 ;
	7'h63 :
		RG_rl_43_t1 = TR_55 ;
	7'h64 :
		RG_rl_43_t1 = TR_55 ;
	7'h65 :
		RG_rl_43_t1 = TR_55 ;
	7'h66 :
		RG_rl_43_t1 = TR_55 ;
	7'h67 :
		RG_rl_43_t1 = TR_55 ;
	7'h68 :
		RG_rl_43_t1 = TR_55 ;
	7'h69 :
		RG_rl_43_t1 = TR_55 ;
	7'h6a :
		RG_rl_43_t1 = TR_55 ;
	7'h6b :
		RG_rl_43_t1 = TR_55 ;
	7'h6c :
		RG_rl_43_t1 = TR_55 ;
	7'h6d :
		RG_rl_43_t1 = TR_55 ;
	7'h6e :
		RG_rl_43_t1 = TR_55 ;
	7'h6f :
		RG_rl_43_t1 = TR_55 ;
	7'h70 :
		RG_rl_43_t1 = TR_55 ;
	7'h71 :
		RG_rl_43_t1 = TR_55 ;
	7'h72 :
		RG_rl_43_t1 = TR_55 ;
	7'h73 :
		RG_rl_43_t1 = TR_55 ;
	7'h74 :
		RG_rl_43_t1 = TR_55 ;
	7'h75 :
		RG_rl_43_t1 = TR_55 ;
	7'h76 :
		RG_rl_43_t1 = TR_55 ;
	7'h77 :
		RG_rl_43_t1 = TR_55 ;
	7'h78 :
		RG_rl_43_t1 = TR_55 ;
	7'h79 :
		RG_rl_43_t1 = TR_55 ;
	7'h7a :
		RG_rl_43_t1 = TR_55 ;
	7'h7b :
		RG_rl_43_t1 = TR_55 ;
	7'h7c :
		RG_rl_43_t1 = TR_55 ;
	7'h7d :
		RG_rl_43_t1 = TR_55 ;
	7'h7e :
		RG_rl_43_t1 = TR_55 ;
	7'h7f :
		RG_rl_43_t1 = TR_55 ;
	default :
		RG_rl_43_t1 = 9'hx ;
	endcase
always @ ( RG_rl_43_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_226 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_43_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h2b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_43_t = ( ( { 9{ U_570 } } & RG_rl_226 )
		| ( { 9{ U_569 } } & RG_rl_43_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_43_en = ( U_570 | RG_rl_43_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_43_en )
		RG_rl_43 <= RG_rl_43_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_56 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_44_t1 = TR_56 ;
	7'h01 :
		RG_rl_44_t1 = TR_56 ;
	7'h02 :
		RG_rl_44_t1 = TR_56 ;
	7'h03 :
		RG_rl_44_t1 = TR_56 ;
	7'h04 :
		RG_rl_44_t1 = TR_56 ;
	7'h05 :
		RG_rl_44_t1 = TR_56 ;
	7'h06 :
		RG_rl_44_t1 = TR_56 ;
	7'h07 :
		RG_rl_44_t1 = TR_56 ;
	7'h08 :
		RG_rl_44_t1 = TR_56 ;
	7'h09 :
		RG_rl_44_t1 = TR_56 ;
	7'h0a :
		RG_rl_44_t1 = TR_56 ;
	7'h0b :
		RG_rl_44_t1 = TR_56 ;
	7'h0c :
		RG_rl_44_t1 = TR_56 ;
	7'h0d :
		RG_rl_44_t1 = TR_56 ;
	7'h0e :
		RG_rl_44_t1 = TR_56 ;
	7'h0f :
		RG_rl_44_t1 = TR_56 ;
	7'h10 :
		RG_rl_44_t1 = TR_56 ;
	7'h11 :
		RG_rl_44_t1 = TR_56 ;
	7'h12 :
		RG_rl_44_t1 = TR_56 ;
	7'h13 :
		RG_rl_44_t1 = TR_56 ;
	7'h14 :
		RG_rl_44_t1 = TR_56 ;
	7'h15 :
		RG_rl_44_t1 = TR_56 ;
	7'h16 :
		RG_rl_44_t1 = TR_56 ;
	7'h17 :
		RG_rl_44_t1 = TR_56 ;
	7'h18 :
		RG_rl_44_t1 = TR_56 ;
	7'h19 :
		RG_rl_44_t1 = TR_56 ;
	7'h1a :
		RG_rl_44_t1 = TR_56 ;
	7'h1b :
		RG_rl_44_t1 = TR_56 ;
	7'h1c :
		RG_rl_44_t1 = TR_56 ;
	7'h1d :
		RG_rl_44_t1 = TR_56 ;
	7'h1e :
		RG_rl_44_t1 = TR_56 ;
	7'h1f :
		RG_rl_44_t1 = TR_56 ;
	7'h20 :
		RG_rl_44_t1 = TR_56 ;
	7'h21 :
		RG_rl_44_t1 = TR_56 ;
	7'h22 :
		RG_rl_44_t1 = TR_56 ;
	7'h23 :
		RG_rl_44_t1 = TR_56 ;
	7'h24 :
		RG_rl_44_t1 = TR_56 ;
	7'h25 :
		RG_rl_44_t1 = TR_56 ;
	7'h26 :
		RG_rl_44_t1 = TR_56 ;
	7'h27 :
		RG_rl_44_t1 = TR_56 ;
	7'h28 :
		RG_rl_44_t1 = TR_56 ;
	7'h29 :
		RG_rl_44_t1 = TR_56 ;
	7'h2a :
		RG_rl_44_t1 = TR_56 ;
	7'h2b :
		RG_rl_44_t1 = TR_56 ;
	7'h2c :
		RG_rl_44_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2d :
		RG_rl_44_t1 = TR_56 ;
	7'h2e :
		RG_rl_44_t1 = TR_56 ;
	7'h2f :
		RG_rl_44_t1 = TR_56 ;
	7'h30 :
		RG_rl_44_t1 = TR_56 ;
	7'h31 :
		RG_rl_44_t1 = TR_56 ;
	7'h32 :
		RG_rl_44_t1 = TR_56 ;
	7'h33 :
		RG_rl_44_t1 = TR_56 ;
	7'h34 :
		RG_rl_44_t1 = TR_56 ;
	7'h35 :
		RG_rl_44_t1 = TR_56 ;
	7'h36 :
		RG_rl_44_t1 = TR_56 ;
	7'h37 :
		RG_rl_44_t1 = TR_56 ;
	7'h38 :
		RG_rl_44_t1 = TR_56 ;
	7'h39 :
		RG_rl_44_t1 = TR_56 ;
	7'h3a :
		RG_rl_44_t1 = TR_56 ;
	7'h3b :
		RG_rl_44_t1 = TR_56 ;
	7'h3c :
		RG_rl_44_t1 = TR_56 ;
	7'h3d :
		RG_rl_44_t1 = TR_56 ;
	7'h3e :
		RG_rl_44_t1 = TR_56 ;
	7'h3f :
		RG_rl_44_t1 = TR_56 ;
	7'h40 :
		RG_rl_44_t1 = TR_56 ;
	7'h41 :
		RG_rl_44_t1 = TR_56 ;
	7'h42 :
		RG_rl_44_t1 = TR_56 ;
	7'h43 :
		RG_rl_44_t1 = TR_56 ;
	7'h44 :
		RG_rl_44_t1 = TR_56 ;
	7'h45 :
		RG_rl_44_t1 = TR_56 ;
	7'h46 :
		RG_rl_44_t1 = TR_56 ;
	7'h47 :
		RG_rl_44_t1 = TR_56 ;
	7'h48 :
		RG_rl_44_t1 = TR_56 ;
	7'h49 :
		RG_rl_44_t1 = TR_56 ;
	7'h4a :
		RG_rl_44_t1 = TR_56 ;
	7'h4b :
		RG_rl_44_t1 = TR_56 ;
	7'h4c :
		RG_rl_44_t1 = TR_56 ;
	7'h4d :
		RG_rl_44_t1 = TR_56 ;
	7'h4e :
		RG_rl_44_t1 = TR_56 ;
	7'h4f :
		RG_rl_44_t1 = TR_56 ;
	7'h50 :
		RG_rl_44_t1 = TR_56 ;
	7'h51 :
		RG_rl_44_t1 = TR_56 ;
	7'h52 :
		RG_rl_44_t1 = TR_56 ;
	7'h53 :
		RG_rl_44_t1 = TR_56 ;
	7'h54 :
		RG_rl_44_t1 = TR_56 ;
	7'h55 :
		RG_rl_44_t1 = TR_56 ;
	7'h56 :
		RG_rl_44_t1 = TR_56 ;
	7'h57 :
		RG_rl_44_t1 = TR_56 ;
	7'h58 :
		RG_rl_44_t1 = TR_56 ;
	7'h59 :
		RG_rl_44_t1 = TR_56 ;
	7'h5a :
		RG_rl_44_t1 = TR_56 ;
	7'h5b :
		RG_rl_44_t1 = TR_56 ;
	7'h5c :
		RG_rl_44_t1 = TR_56 ;
	7'h5d :
		RG_rl_44_t1 = TR_56 ;
	7'h5e :
		RG_rl_44_t1 = TR_56 ;
	7'h5f :
		RG_rl_44_t1 = TR_56 ;
	7'h60 :
		RG_rl_44_t1 = TR_56 ;
	7'h61 :
		RG_rl_44_t1 = TR_56 ;
	7'h62 :
		RG_rl_44_t1 = TR_56 ;
	7'h63 :
		RG_rl_44_t1 = TR_56 ;
	7'h64 :
		RG_rl_44_t1 = TR_56 ;
	7'h65 :
		RG_rl_44_t1 = TR_56 ;
	7'h66 :
		RG_rl_44_t1 = TR_56 ;
	7'h67 :
		RG_rl_44_t1 = TR_56 ;
	7'h68 :
		RG_rl_44_t1 = TR_56 ;
	7'h69 :
		RG_rl_44_t1 = TR_56 ;
	7'h6a :
		RG_rl_44_t1 = TR_56 ;
	7'h6b :
		RG_rl_44_t1 = TR_56 ;
	7'h6c :
		RG_rl_44_t1 = TR_56 ;
	7'h6d :
		RG_rl_44_t1 = TR_56 ;
	7'h6e :
		RG_rl_44_t1 = TR_56 ;
	7'h6f :
		RG_rl_44_t1 = TR_56 ;
	7'h70 :
		RG_rl_44_t1 = TR_56 ;
	7'h71 :
		RG_rl_44_t1 = TR_56 ;
	7'h72 :
		RG_rl_44_t1 = TR_56 ;
	7'h73 :
		RG_rl_44_t1 = TR_56 ;
	7'h74 :
		RG_rl_44_t1 = TR_56 ;
	7'h75 :
		RG_rl_44_t1 = TR_56 ;
	7'h76 :
		RG_rl_44_t1 = TR_56 ;
	7'h77 :
		RG_rl_44_t1 = TR_56 ;
	7'h78 :
		RG_rl_44_t1 = TR_56 ;
	7'h79 :
		RG_rl_44_t1 = TR_56 ;
	7'h7a :
		RG_rl_44_t1 = TR_56 ;
	7'h7b :
		RG_rl_44_t1 = TR_56 ;
	7'h7c :
		RG_rl_44_t1 = TR_56 ;
	7'h7d :
		RG_rl_44_t1 = TR_56 ;
	7'h7e :
		RG_rl_44_t1 = TR_56 ;
	7'h7f :
		RG_rl_44_t1 = TR_56 ;
	default :
		RG_rl_44_t1 = 9'hx ;
	endcase
always @ ( RG_rl_44_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_227 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_44_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h2c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_44_t = ( ( { 9{ U_570 } } & RG_rl_227 )
		| ( { 9{ U_569 } } & RG_rl_44_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_44_en = ( U_570 | RG_rl_44_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_44_en )
		RG_rl_44 <= RG_rl_44_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_57 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_45_t1 = TR_57 ;
	7'h01 :
		RG_rl_45_t1 = TR_57 ;
	7'h02 :
		RG_rl_45_t1 = TR_57 ;
	7'h03 :
		RG_rl_45_t1 = TR_57 ;
	7'h04 :
		RG_rl_45_t1 = TR_57 ;
	7'h05 :
		RG_rl_45_t1 = TR_57 ;
	7'h06 :
		RG_rl_45_t1 = TR_57 ;
	7'h07 :
		RG_rl_45_t1 = TR_57 ;
	7'h08 :
		RG_rl_45_t1 = TR_57 ;
	7'h09 :
		RG_rl_45_t1 = TR_57 ;
	7'h0a :
		RG_rl_45_t1 = TR_57 ;
	7'h0b :
		RG_rl_45_t1 = TR_57 ;
	7'h0c :
		RG_rl_45_t1 = TR_57 ;
	7'h0d :
		RG_rl_45_t1 = TR_57 ;
	7'h0e :
		RG_rl_45_t1 = TR_57 ;
	7'h0f :
		RG_rl_45_t1 = TR_57 ;
	7'h10 :
		RG_rl_45_t1 = TR_57 ;
	7'h11 :
		RG_rl_45_t1 = TR_57 ;
	7'h12 :
		RG_rl_45_t1 = TR_57 ;
	7'h13 :
		RG_rl_45_t1 = TR_57 ;
	7'h14 :
		RG_rl_45_t1 = TR_57 ;
	7'h15 :
		RG_rl_45_t1 = TR_57 ;
	7'h16 :
		RG_rl_45_t1 = TR_57 ;
	7'h17 :
		RG_rl_45_t1 = TR_57 ;
	7'h18 :
		RG_rl_45_t1 = TR_57 ;
	7'h19 :
		RG_rl_45_t1 = TR_57 ;
	7'h1a :
		RG_rl_45_t1 = TR_57 ;
	7'h1b :
		RG_rl_45_t1 = TR_57 ;
	7'h1c :
		RG_rl_45_t1 = TR_57 ;
	7'h1d :
		RG_rl_45_t1 = TR_57 ;
	7'h1e :
		RG_rl_45_t1 = TR_57 ;
	7'h1f :
		RG_rl_45_t1 = TR_57 ;
	7'h20 :
		RG_rl_45_t1 = TR_57 ;
	7'h21 :
		RG_rl_45_t1 = TR_57 ;
	7'h22 :
		RG_rl_45_t1 = TR_57 ;
	7'h23 :
		RG_rl_45_t1 = TR_57 ;
	7'h24 :
		RG_rl_45_t1 = TR_57 ;
	7'h25 :
		RG_rl_45_t1 = TR_57 ;
	7'h26 :
		RG_rl_45_t1 = TR_57 ;
	7'h27 :
		RG_rl_45_t1 = TR_57 ;
	7'h28 :
		RG_rl_45_t1 = TR_57 ;
	7'h29 :
		RG_rl_45_t1 = TR_57 ;
	7'h2a :
		RG_rl_45_t1 = TR_57 ;
	7'h2b :
		RG_rl_45_t1 = TR_57 ;
	7'h2c :
		RG_rl_45_t1 = TR_57 ;
	7'h2d :
		RG_rl_45_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2e :
		RG_rl_45_t1 = TR_57 ;
	7'h2f :
		RG_rl_45_t1 = TR_57 ;
	7'h30 :
		RG_rl_45_t1 = TR_57 ;
	7'h31 :
		RG_rl_45_t1 = TR_57 ;
	7'h32 :
		RG_rl_45_t1 = TR_57 ;
	7'h33 :
		RG_rl_45_t1 = TR_57 ;
	7'h34 :
		RG_rl_45_t1 = TR_57 ;
	7'h35 :
		RG_rl_45_t1 = TR_57 ;
	7'h36 :
		RG_rl_45_t1 = TR_57 ;
	7'h37 :
		RG_rl_45_t1 = TR_57 ;
	7'h38 :
		RG_rl_45_t1 = TR_57 ;
	7'h39 :
		RG_rl_45_t1 = TR_57 ;
	7'h3a :
		RG_rl_45_t1 = TR_57 ;
	7'h3b :
		RG_rl_45_t1 = TR_57 ;
	7'h3c :
		RG_rl_45_t1 = TR_57 ;
	7'h3d :
		RG_rl_45_t1 = TR_57 ;
	7'h3e :
		RG_rl_45_t1 = TR_57 ;
	7'h3f :
		RG_rl_45_t1 = TR_57 ;
	7'h40 :
		RG_rl_45_t1 = TR_57 ;
	7'h41 :
		RG_rl_45_t1 = TR_57 ;
	7'h42 :
		RG_rl_45_t1 = TR_57 ;
	7'h43 :
		RG_rl_45_t1 = TR_57 ;
	7'h44 :
		RG_rl_45_t1 = TR_57 ;
	7'h45 :
		RG_rl_45_t1 = TR_57 ;
	7'h46 :
		RG_rl_45_t1 = TR_57 ;
	7'h47 :
		RG_rl_45_t1 = TR_57 ;
	7'h48 :
		RG_rl_45_t1 = TR_57 ;
	7'h49 :
		RG_rl_45_t1 = TR_57 ;
	7'h4a :
		RG_rl_45_t1 = TR_57 ;
	7'h4b :
		RG_rl_45_t1 = TR_57 ;
	7'h4c :
		RG_rl_45_t1 = TR_57 ;
	7'h4d :
		RG_rl_45_t1 = TR_57 ;
	7'h4e :
		RG_rl_45_t1 = TR_57 ;
	7'h4f :
		RG_rl_45_t1 = TR_57 ;
	7'h50 :
		RG_rl_45_t1 = TR_57 ;
	7'h51 :
		RG_rl_45_t1 = TR_57 ;
	7'h52 :
		RG_rl_45_t1 = TR_57 ;
	7'h53 :
		RG_rl_45_t1 = TR_57 ;
	7'h54 :
		RG_rl_45_t1 = TR_57 ;
	7'h55 :
		RG_rl_45_t1 = TR_57 ;
	7'h56 :
		RG_rl_45_t1 = TR_57 ;
	7'h57 :
		RG_rl_45_t1 = TR_57 ;
	7'h58 :
		RG_rl_45_t1 = TR_57 ;
	7'h59 :
		RG_rl_45_t1 = TR_57 ;
	7'h5a :
		RG_rl_45_t1 = TR_57 ;
	7'h5b :
		RG_rl_45_t1 = TR_57 ;
	7'h5c :
		RG_rl_45_t1 = TR_57 ;
	7'h5d :
		RG_rl_45_t1 = TR_57 ;
	7'h5e :
		RG_rl_45_t1 = TR_57 ;
	7'h5f :
		RG_rl_45_t1 = TR_57 ;
	7'h60 :
		RG_rl_45_t1 = TR_57 ;
	7'h61 :
		RG_rl_45_t1 = TR_57 ;
	7'h62 :
		RG_rl_45_t1 = TR_57 ;
	7'h63 :
		RG_rl_45_t1 = TR_57 ;
	7'h64 :
		RG_rl_45_t1 = TR_57 ;
	7'h65 :
		RG_rl_45_t1 = TR_57 ;
	7'h66 :
		RG_rl_45_t1 = TR_57 ;
	7'h67 :
		RG_rl_45_t1 = TR_57 ;
	7'h68 :
		RG_rl_45_t1 = TR_57 ;
	7'h69 :
		RG_rl_45_t1 = TR_57 ;
	7'h6a :
		RG_rl_45_t1 = TR_57 ;
	7'h6b :
		RG_rl_45_t1 = TR_57 ;
	7'h6c :
		RG_rl_45_t1 = TR_57 ;
	7'h6d :
		RG_rl_45_t1 = TR_57 ;
	7'h6e :
		RG_rl_45_t1 = TR_57 ;
	7'h6f :
		RG_rl_45_t1 = TR_57 ;
	7'h70 :
		RG_rl_45_t1 = TR_57 ;
	7'h71 :
		RG_rl_45_t1 = TR_57 ;
	7'h72 :
		RG_rl_45_t1 = TR_57 ;
	7'h73 :
		RG_rl_45_t1 = TR_57 ;
	7'h74 :
		RG_rl_45_t1 = TR_57 ;
	7'h75 :
		RG_rl_45_t1 = TR_57 ;
	7'h76 :
		RG_rl_45_t1 = TR_57 ;
	7'h77 :
		RG_rl_45_t1 = TR_57 ;
	7'h78 :
		RG_rl_45_t1 = TR_57 ;
	7'h79 :
		RG_rl_45_t1 = TR_57 ;
	7'h7a :
		RG_rl_45_t1 = TR_57 ;
	7'h7b :
		RG_rl_45_t1 = TR_57 ;
	7'h7c :
		RG_rl_45_t1 = TR_57 ;
	7'h7d :
		RG_rl_45_t1 = TR_57 ;
	7'h7e :
		RG_rl_45_t1 = TR_57 ;
	7'h7f :
		RG_rl_45_t1 = TR_57 ;
	default :
		RG_rl_45_t1 = 9'hx ;
	endcase
always @ ( RG_rl_45_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_228 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_45_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h2d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_45_t = ( ( { 9{ U_570 } } & RG_rl_228 )
		| ( { 9{ U_569 } } & RG_rl_45_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_45_en = ( U_570 | RG_rl_45_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_45_en )
		RG_rl_45 <= RG_rl_45_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_58 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_46_t1 = TR_58 ;
	7'h01 :
		RG_rl_46_t1 = TR_58 ;
	7'h02 :
		RG_rl_46_t1 = TR_58 ;
	7'h03 :
		RG_rl_46_t1 = TR_58 ;
	7'h04 :
		RG_rl_46_t1 = TR_58 ;
	7'h05 :
		RG_rl_46_t1 = TR_58 ;
	7'h06 :
		RG_rl_46_t1 = TR_58 ;
	7'h07 :
		RG_rl_46_t1 = TR_58 ;
	7'h08 :
		RG_rl_46_t1 = TR_58 ;
	7'h09 :
		RG_rl_46_t1 = TR_58 ;
	7'h0a :
		RG_rl_46_t1 = TR_58 ;
	7'h0b :
		RG_rl_46_t1 = TR_58 ;
	7'h0c :
		RG_rl_46_t1 = TR_58 ;
	7'h0d :
		RG_rl_46_t1 = TR_58 ;
	7'h0e :
		RG_rl_46_t1 = TR_58 ;
	7'h0f :
		RG_rl_46_t1 = TR_58 ;
	7'h10 :
		RG_rl_46_t1 = TR_58 ;
	7'h11 :
		RG_rl_46_t1 = TR_58 ;
	7'h12 :
		RG_rl_46_t1 = TR_58 ;
	7'h13 :
		RG_rl_46_t1 = TR_58 ;
	7'h14 :
		RG_rl_46_t1 = TR_58 ;
	7'h15 :
		RG_rl_46_t1 = TR_58 ;
	7'h16 :
		RG_rl_46_t1 = TR_58 ;
	7'h17 :
		RG_rl_46_t1 = TR_58 ;
	7'h18 :
		RG_rl_46_t1 = TR_58 ;
	7'h19 :
		RG_rl_46_t1 = TR_58 ;
	7'h1a :
		RG_rl_46_t1 = TR_58 ;
	7'h1b :
		RG_rl_46_t1 = TR_58 ;
	7'h1c :
		RG_rl_46_t1 = TR_58 ;
	7'h1d :
		RG_rl_46_t1 = TR_58 ;
	7'h1e :
		RG_rl_46_t1 = TR_58 ;
	7'h1f :
		RG_rl_46_t1 = TR_58 ;
	7'h20 :
		RG_rl_46_t1 = TR_58 ;
	7'h21 :
		RG_rl_46_t1 = TR_58 ;
	7'h22 :
		RG_rl_46_t1 = TR_58 ;
	7'h23 :
		RG_rl_46_t1 = TR_58 ;
	7'h24 :
		RG_rl_46_t1 = TR_58 ;
	7'h25 :
		RG_rl_46_t1 = TR_58 ;
	7'h26 :
		RG_rl_46_t1 = TR_58 ;
	7'h27 :
		RG_rl_46_t1 = TR_58 ;
	7'h28 :
		RG_rl_46_t1 = TR_58 ;
	7'h29 :
		RG_rl_46_t1 = TR_58 ;
	7'h2a :
		RG_rl_46_t1 = TR_58 ;
	7'h2b :
		RG_rl_46_t1 = TR_58 ;
	7'h2c :
		RG_rl_46_t1 = TR_58 ;
	7'h2d :
		RG_rl_46_t1 = TR_58 ;
	7'h2e :
		RG_rl_46_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h2f :
		RG_rl_46_t1 = TR_58 ;
	7'h30 :
		RG_rl_46_t1 = TR_58 ;
	7'h31 :
		RG_rl_46_t1 = TR_58 ;
	7'h32 :
		RG_rl_46_t1 = TR_58 ;
	7'h33 :
		RG_rl_46_t1 = TR_58 ;
	7'h34 :
		RG_rl_46_t1 = TR_58 ;
	7'h35 :
		RG_rl_46_t1 = TR_58 ;
	7'h36 :
		RG_rl_46_t1 = TR_58 ;
	7'h37 :
		RG_rl_46_t1 = TR_58 ;
	7'h38 :
		RG_rl_46_t1 = TR_58 ;
	7'h39 :
		RG_rl_46_t1 = TR_58 ;
	7'h3a :
		RG_rl_46_t1 = TR_58 ;
	7'h3b :
		RG_rl_46_t1 = TR_58 ;
	7'h3c :
		RG_rl_46_t1 = TR_58 ;
	7'h3d :
		RG_rl_46_t1 = TR_58 ;
	7'h3e :
		RG_rl_46_t1 = TR_58 ;
	7'h3f :
		RG_rl_46_t1 = TR_58 ;
	7'h40 :
		RG_rl_46_t1 = TR_58 ;
	7'h41 :
		RG_rl_46_t1 = TR_58 ;
	7'h42 :
		RG_rl_46_t1 = TR_58 ;
	7'h43 :
		RG_rl_46_t1 = TR_58 ;
	7'h44 :
		RG_rl_46_t1 = TR_58 ;
	7'h45 :
		RG_rl_46_t1 = TR_58 ;
	7'h46 :
		RG_rl_46_t1 = TR_58 ;
	7'h47 :
		RG_rl_46_t1 = TR_58 ;
	7'h48 :
		RG_rl_46_t1 = TR_58 ;
	7'h49 :
		RG_rl_46_t1 = TR_58 ;
	7'h4a :
		RG_rl_46_t1 = TR_58 ;
	7'h4b :
		RG_rl_46_t1 = TR_58 ;
	7'h4c :
		RG_rl_46_t1 = TR_58 ;
	7'h4d :
		RG_rl_46_t1 = TR_58 ;
	7'h4e :
		RG_rl_46_t1 = TR_58 ;
	7'h4f :
		RG_rl_46_t1 = TR_58 ;
	7'h50 :
		RG_rl_46_t1 = TR_58 ;
	7'h51 :
		RG_rl_46_t1 = TR_58 ;
	7'h52 :
		RG_rl_46_t1 = TR_58 ;
	7'h53 :
		RG_rl_46_t1 = TR_58 ;
	7'h54 :
		RG_rl_46_t1 = TR_58 ;
	7'h55 :
		RG_rl_46_t1 = TR_58 ;
	7'h56 :
		RG_rl_46_t1 = TR_58 ;
	7'h57 :
		RG_rl_46_t1 = TR_58 ;
	7'h58 :
		RG_rl_46_t1 = TR_58 ;
	7'h59 :
		RG_rl_46_t1 = TR_58 ;
	7'h5a :
		RG_rl_46_t1 = TR_58 ;
	7'h5b :
		RG_rl_46_t1 = TR_58 ;
	7'h5c :
		RG_rl_46_t1 = TR_58 ;
	7'h5d :
		RG_rl_46_t1 = TR_58 ;
	7'h5e :
		RG_rl_46_t1 = TR_58 ;
	7'h5f :
		RG_rl_46_t1 = TR_58 ;
	7'h60 :
		RG_rl_46_t1 = TR_58 ;
	7'h61 :
		RG_rl_46_t1 = TR_58 ;
	7'h62 :
		RG_rl_46_t1 = TR_58 ;
	7'h63 :
		RG_rl_46_t1 = TR_58 ;
	7'h64 :
		RG_rl_46_t1 = TR_58 ;
	7'h65 :
		RG_rl_46_t1 = TR_58 ;
	7'h66 :
		RG_rl_46_t1 = TR_58 ;
	7'h67 :
		RG_rl_46_t1 = TR_58 ;
	7'h68 :
		RG_rl_46_t1 = TR_58 ;
	7'h69 :
		RG_rl_46_t1 = TR_58 ;
	7'h6a :
		RG_rl_46_t1 = TR_58 ;
	7'h6b :
		RG_rl_46_t1 = TR_58 ;
	7'h6c :
		RG_rl_46_t1 = TR_58 ;
	7'h6d :
		RG_rl_46_t1 = TR_58 ;
	7'h6e :
		RG_rl_46_t1 = TR_58 ;
	7'h6f :
		RG_rl_46_t1 = TR_58 ;
	7'h70 :
		RG_rl_46_t1 = TR_58 ;
	7'h71 :
		RG_rl_46_t1 = TR_58 ;
	7'h72 :
		RG_rl_46_t1 = TR_58 ;
	7'h73 :
		RG_rl_46_t1 = TR_58 ;
	7'h74 :
		RG_rl_46_t1 = TR_58 ;
	7'h75 :
		RG_rl_46_t1 = TR_58 ;
	7'h76 :
		RG_rl_46_t1 = TR_58 ;
	7'h77 :
		RG_rl_46_t1 = TR_58 ;
	7'h78 :
		RG_rl_46_t1 = TR_58 ;
	7'h79 :
		RG_rl_46_t1 = TR_58 ;
	7'h7a :
		RG_rl_46_t1 = TR_58 ;
	7'h7b :
		RG_rl_46_t1 = TR_58 ;
	7'h7c :
		RG_rl_46_t1 = TR_58 ;
	7'h7d :
		RG_rl_46_t1 = TR_58 ;
	7'h7e :
		RG_rl_46_t1 = TR_58 ;
	7'h7f :
		RG_rl_46_t1 = TR_58 ;
	default :
		RG_rl_46_t1 = 9'hx ;
	endcase
always @ ( RG_rl_46_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_229 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_46_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h2e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_46_t = ( ( { 9{ U_570 } } & RG_rl_229 )
		| ( { 9{ U_569 } } & RG_rl_46_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_46_en = ( U_570 | RG_rl_46_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_46_en )
		RG_rl_46 <= RG_rl_46_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_59 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_47_t1 = TR_59 ;
	7'h01 :
		RG_rl_47_t1 = TR_59 ;
	7'h02 :
		RG_rl_47_t1 = TR_59 ;
	7'h03 :
		RG_rl_47_t1 = TR_59 ;
	7'h04 :
		RG_rl_47_t1 = TR_59 ;
	7'h05 :
		RG_rl_47_t1 = TR_59 ;
	7'h06 :
		RG_rl_47_t1 = TR_59 ;
	7'h07 :
		RG_rl_47_t1 = TR_59 ;
	7'h08 :
		RG_rl_47_t1 = TR_59 ;
	7'h09 :
		RG_rl_47_t1 = TR_59 ;
	7'h0a :
		RG_rl_47_t1 = TR_59 ;
	7'h0b :
		RG_rl_47_t1 = TR_59 ;
	7'h0c :
		RG_rl_47_t1 = TR_59 ;
	7'h0d :
		RG_rl_47_t1 = TR_59 ;
	7'h0e :
		RG_rl_47_t1 = TR_59 ;
	7'h0f :
		RG_rl_47_t1 = TR_59 ;
	7'h10 :
		RG_rl_47_t1 = TR_59 ;
	7'h11 :
		RG_rl_47_t1 = TR_59 ;
	7'h12 :
		RG_rl_47_t1 = TR_59 ;
	7'h13 :
		RG_rl_47_t1 = TR_59 ;
	7'h14 :
		RG_rl_47_t1 = TR_59 ;
	7'h15 :
		RG_rl_47_t1 = TR_59 ;
	7'h16 :
		RG_rl_47_t1 = TR_59 ;
	7'h17 :
		RG_rl_47_t1 = TR_59 ;
	7'h18 :
		RG_rl_47_t1 = TR_59 ;
	7'h19 :
		RG_rl_47_t1 = TR_59 ;
	7'h1a :
		RG_rl_47_t1 = TR_59 ;
	7'h1b :
		RG_rl_47_t1 = TR_59 ;
	7'h1c :
		RG_rl_47_t1 = TR_59 ;
	7'h1d :
		RG_rl_47_t1 = TR_59 ;
	7'h1e :
		RG_rl_47_t1 = TR_59 ;
	7'h1f :
		RG_rl_47_t1 = TR_59 ;
	7'h20 :
		RG_rl_47_t1 = TR_59 ;
	7'h21 :
		RG_rl_47_t1 = TR_59 ;
	7'h22 :
		RG_rl_47_t1 = TR_59 ;
	7'h23 :
		RG_rl_47_t1 = TR_59 ;
	7'h24 :
		RG_rl_47_t1 = TR_59 ;
	7'h25 :
		RG_rl_47_t1 = TR_59 ;
	7'h26 :
		RG_rl_47_t1 = TR_59 ;
	7'h27 :
		RG_rl_47_t1 = TR_59 ;
	7'h28 :
		RG_rl_47_t1 = TR_59 ;
	7'h29 :
		RG_rl_47_t1 = TR_59 ;
	7'h2a :
		RG_rl_47_t1 = TR_59 ;
	7'h2b :
		RG_rl_47_t1 = TR_59 ;
	7'h2c :
		RG_rl_47_t1 = TR_59 ;
	7'h2d :
		RG_rl_47_t1 = TR_59 ;
	7'h2e :
		RG_rl_47_t1 = TR_59 ;
	7'h2f :
		RG_rl_47_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h30 :
		RG_rl_47_t1 = TR_59 ;
	7'h31 :
		RG_rl_47_t1 = TR_59 ;
	7'h32 :
		RG_rl_47_t1 = TR_59 ;
	7'h33 :
		RG_rl_47_t1 = TR_59 ;
	7'h34 :
		RG_rl_47_t1 = TR_59 ;
	7'h35 :
		RG_rl_47_t1 = TR_59 ;
	7'h36 :
		RG_rl_47_t1 = TR_59 ;
	7'h37 :
		RG_rl_47_t1 = TR_59 ;
	7'h38 :
		RG_rl_47_t1 = TR_59 ;
	7'h39 :
		RG_rl_47_t1 = TR_59 ;
	7'h3a :
		RG_rl_47_t1 = TR_59 ;
	7'h3b :
		RG_rl_47_t1 = TR_59 ;
	7'h3c :
		RG_rl_47_t1 = TR_59 ;
	7'h3d :
		RG_rl_47_t1 = TR_59 ;
	7'h3e :
		RG_rl_47_t1 = TR_59 ;
	7'h3f :
		RG_rl_47_t1 = TR_59 ;
	7'h40 :
		RG_rl_47_t1 = TR_59 ;
	7'h41 :
		RG_rl_47_t1 = TR_59 ;
	7'h42 :
		RG_rl_47_t1 = TR_59 ;
	7'h43 :
		RG_rl_47_t1 = TR_59 ;
	7'h44 :
		RG_rl_47_t1 = TR_59 ;
	7'h45 :
		RG_rl_47_t1 = TR_59 ;
	7'h46 :
		RG_rl_47_t1 = TR_59 ;
	7'h47 :
		RG_rl_47_t1 = TR_59 ;
	7'h48 :
		RG_rl_47_t1 = TR_59 ;
	7'h49 :
		RG_rl_47_t1 = TR_59 ;
	7'h4a :
		RG_rl_47_t1 = TR_59 ;
	7'h4b :
		RG_rl_47_t1 = TR_59 ;
	7'h4c :
		RG_rl_47_t1 = TR_59 ;
	7'h4d :
		RG_rl_47_t1 = TR_59 ;
	7'h4e :
		RG_rl_47_t1 = TR_59 ;
	7'h4f :
		RG_rl_47_t1 = TR_59 ;
	7'h50 :
		RG_rl_47_t1 = TR_59 ;
	7'h51 :
		RG_rl_47_t1 = TR_59 ;
	7'h52 :
		RG_rl_47_t1 = TR_59 ;
	7'h53 :
		RG_rl_47_t1 = TR_59 ;
	7'h54 :
		RG_rl_47_t1 = TR_59 ;
	7'h55 :
		RG_rl_47_t1 = TR_59 ;
	7'h56 :
		RG_rl_47_t1 = TR_59 ;
	7'h57 :
		RG_rl_47_t1 = TR_59 ;
	7'h58 :
		RG_rl_47_t1 = TR_59 ;
	7'h59 :
		RG_rl_47_t1 = TR_59 ;
	7'h5a :
		RG_rl_47_t1 = TR_59 ;
	7'h5b :
		RG_rl_47_t1 = TR_59 ;
	7'h5c :
		RG_rl_47_t1 = TR_59 ;
	7'h5d :
		RG_rl_47_t1 = TR_59 ;
	7'h5e :
		RG_rl_47_t1 = TR_59 ;
	7'h5f :
		RG_rl_47_t1 = TR_59 ;
	7'h60 :
		RG_rl_47_t1 = TR_59 ;
	7'h61 :
		RG_rl_47_t1 = TR_59 ;
	7'h62 :
		RG_rl_47_t1 = TR_59 ;
	7'h63 :
		RG_rl_47_t1 = TR_59 ;
	7'h64 :
		RG_rl_47_t1 = TR_59 ;
	7'h65 :
		RG_rl_47_t1 = TR_59 ;
	7'h66 :
		RG_rl_47_t1 = TR_59 ;
	7'h67 :
		RG_rl_47_t1 = TR_59 ;
	7'h68 :
		RG_rl_47_t1 = TR_59 ;
	7'h69 :
		RG_rl_47_t1 = TR_59 ;
	7'h6a :
		RG_rl_47_t1 = TR_59 ;
	7'h6b :
		RG_rl_47_t1 = TR_59 ;
	7'h6c :
		RG_rl_47_t1 = TR_59 ;
	7'h6d :
		RG_rl_47_t1 = TR_59 ;
	7'h6e :
		RG_rl_47_t1 = TR_59 ;
	7'h6f :
		RG_rl_47_t1 = TR_59 ;
	7'h70 :
		RG_rl_47_t1 = TR_59 ;
	7'h71 :
		RG_rl_47_t1 = TR_59 ;
	7'h72 :
		RG_rl_47_t1 = TR_59 ;
	7'h73 :
		RG_rl_47_t1 = TR_59 ;
	7'h74 :
		RG_rl_47_t1 = TR_59 ;
	7'h75 :
		RG_rl_47_t1 = TR_59 ;
	7'h76 :
		RG_rl_47_t1 = TR_59 ;
	7'h77 :
		RG_rl_47_t1 = TR_59 ;
	7'h78 :
		RG_rl_47_t1 = TR_59 ;
	7'h79 :
		RG_rl_47_t1 = TR_59 ;
	7'h7a :
		RG_rl_47_t1 = TR_59 ;
	7'h7b :
		RG_rl_47_t1 = TR_59 ;
	7'h7c :
		RG_rl_47_t1 = TR_59 ;
	7'h7d :
		RG_rl_47_t1 = TR_59 ;
	7'h7e :
		RG_rl_47_t1 = TR_59 ;
	7'h7f :
		RG_rl_47_t1 = TR_59 ;
	default :
		RG_rl_47_t1 = 9'hx ;
	endcase
always @ ( RG_rl_47_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_230 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_47_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h2f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_47_t = ( ( { 9{ U_570 } } & RG_rl_230 )
		| ( { 9{ U_569 } } & RG_rl_47_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_47_en = ( U_570 | RG_rl_47_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_47_en )
		RG_rl_47 <= RG_rl_47_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_60 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_48_t1 = TR_60 ;
	7'h01 :
		RG_rl_48_t1 = TR_60 ;
	7'h02 :
		RG_rl_48_t1 = TR_60 ;
	7'h03 :
		RG_rl_48_t1 = TR_60 ;
	7'h04 :
		RG_rl_48_t1 = TR_60 ;
	7'h05 :
		RG_rl_48_t1 = TR_60 ;
	7'h06 :
		RG_rl_48_t1 = TR_60 ;
	7'h07 :
		RG_rl_48_t1 = TR_60 ;
	7'h08 :
		RG_rl_48_t1 = TR_60 ;
	7'h09 :
		RG_rl_48_t1 = TR_60 ;
	7'h0a :
		RG_rl_48_t1 = TR_60 ;
	7'h0b :
		RG_rl_48_t1 = TR_60 ;
	7'h0c :
		RG_rl_48_t1 = TR_60 ;
	7'h0d :
		RG_rl_48_t1 = TR_60 ;
	7'h0e :
		RG_rl_48_t1 = TR_60 ;
	7'h0f :
		RG_rl_48_t1 = TR_60 ;
	7'h10 :
		RG_rl_48_t1 = TR_60 ;
	7'h11 :
		RG_rl_48_t1 = TR_60 ;
	7'h12 :
		RG_rl_48_t1 = TR_60 ;
	7'h13 :
		RG_rl_48_t1 = TR_60 ;
	7'h14 :
		RG_rl_48_t1 = TR_60 ;
	7'h15 :
		RG_rl_48_t1 = TR_60 ;
	7'h16 :
		RG_rl_48_t1 = TR_60 ;
	7'h17 :
		RG_rl_48_t1 = TR_60 ;
	7'h18 :
		RG_rl_48_t1 = TR_60 ;
	7'h19 :
		RG_rl_48_t1 = TR_60 ;
	7'h1a :
		RG_rl_48_t1 = TR_60 ;
	7'h1b :
		RG_rl_48_t1 = TR_60 ;
	7'h1c :
		RG_rl_48_t1 = TR_60 ;
	7'h1d :
		RG_rl_48_t1 = TR_60 ;
	7'h1e :
		RG_rl_48_t1 = TR_60 ;
	7'h1f :
		RG_rl_48_t1 = TR_60 ;
	7'h20 :
		RG_rl_48_t1 = TR_60 ;
	7'h21 :
		RG_rl_48_t1 = TR_60 ;
	7'h22 :
		RG_rl_48_t1 = TR_60 ;
	7'h23 :
		RG_rl_48_t1 = TR_60 ;
	7'h24 :
		RG_rl_48_t1 = TR_60 ;
	7'h25 :
		RG_rl_48_t1 = TR_60 ;
	7'h26 :
		RG_rl_48_t1 = TR_60 ;
	7'h27 :
		RG_rl_48_t1 = TR_60 ;
	7'h28 :
		RG_rl_48_t1 = TR_60 ;
	7'h29 :
		RG_rl_48_t1 = TR_60 ;
	7'h2a :
		RG_rl_48_t1 = TR_60 ;
	7'h2b :
		RG_rl_48_t1 = TR_60 ;
	7'h2c :
		RG_rl_48_t1 = TR_60 ;
	7'h2d :
		RG_rl_48_t1 = TR_60 ;
	7'h2e :
		RG_rl_48_t1 = TR_60 ;
	7'h2f :
		RG_rl_48_t1 = TR_60 ;
	7'h30 :
		RG_rl_48_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h31 :
		RG_rl_48_t1 = TR_60 ;
	7'h32 :
		RG_rl_48_t1 = TR_60 ;
	7'h33 :
		RG_rl_48_t1 = TR_60 ;
	7'h34 :
		RG_rl_48_t1 = TR_60 ;
	7'h35 :
		RG_rl_48_t1 = TR_60 ;
	7'h36 :
		RG_rl_48_t1 = TR_60 ;
	7'h37 :
		RG_rl_48_t1 = TR_60 ;
	7'h38 :
		RG_rl_48_t1 = TR_60 ;
	7'h39 :
		RG_rl_48_t1 = TR_60 ;
	7'h3a :
		RG_rl_48_t1 = TR_60 ;
	7'h3b :
		RG_rl_48_t1 = TR_60 ;
	7'h3c :
		RG_rl_48_t1 = TR_60 ;
	7'h3d :
		RG_rl_48_t1 = TR_60 ;
	7'h3e :
		RG_rl_48_t1 = TR_60 ;
	7'h3f :
		RG_rl_48_t1 = TR_60 ;
	7'h40 :
		RG_rl_48_t1 = TR_60 ;
	7'h41 :
		RG_rl_48_t1 = TR_60 ;
	7'h42 :
		RG_rl_48_t1 = TR_60 ;
	7'h43 :
		RG_rl_48_t1 = TR_60 ;
	7'h44 :
		RG_rl_48_t1 = TR_60 ;
	7'h45 :
		RG_rl_48_t1 = TR_60 ;
	7'h46 :
		RG_rl_48_t1 = TR_60 ;
	7'h47 :
		RG_rl_48_t1 = TR_60 ;
	7'h48 :
		RG_rl_48_t1 = TR_60 ;
	7'h49 :
		RG_rl_48_t1 = TR_60 ;
	7'h4a :
		RG_rl_48_t1 = TR_60 ;
	7'h4b :
		RG_rl_48_t1 = TR_60 ;
	7'h4c :
		RG_rl_48_t1 = TR_60 ;
	7'h4d :
		RG_rl_48_t1 = TR_60 ;
	7'h4e :
		RG_rl_48_t1 = TR_60 ;
	7'h4f :
		RG_rl_48_t1 = TR_60 ;
	7'h50 :
		RG_rl_48_t1 = TR_60 ;
	7'h51 :
		RG_rl_48_t1 = TR_60 ;
	7'h52 :
		RG_rl_48_t1 = TR_60 ;
	7'h53 :
		RG_rl_48_t1 = TR_60 ;
	7'h54 :
		RG_rl_48_t1 = TR_60 ;
	7'h55 :
		RG_rl_48_t1 = TR_60 ;
	7'h56 :
		RG_rl_48_t1 = TR_60 ;
	7'h57 :
		RG_rl_48_t1 = TR_60 ;
	7'h58 :
		RG_rl_48_t1 = TR_60 ;
	7'h59 :
		RG_rl_48_t1 = TR_60 ;
	7'h5a :
		RG_rl_48_t1 = TR_60 ;
	7'h5b :
		RG_rl_48_t1 = TR_60 ;
	7'h5c :
		RG_rl_48_t1 = TR_60 ;
	7'h5d :
		RG_rl_48_t1 = TR_60 ;
	7'h5e :
		RG_rl_48_t1 = TR_60 ;
	7'h5f :
		RG_rl_48_t1 = TR_60 ;
	7'h60 :
		RG_rl_48_t1 = TR_60 ;
	7'h61 :
		RG_rl_48_t1 = TR_60 ;
	7'h62 :
		RG_rl_48_t1 = TR_60 ;
	7'h63 :
		RG_rl_48_t1 = TR_60 ;
	7'h64 :
		RG_rl_48_t1 = TR_60 ;
	7'h65 :
		RG_rl_48_t1 = TR_60 ;
	7'h66 :
		RG_rl_48_t1 = TR_60 ;
	7'h67 :
		RG_rl_48_t1 = TR_60 ;
	7'h68 :
		RG_rl_48_t1 = TR_60 ;
	7'h69 :
		RG_rl_48_t1 = TR_60 ;
	7'h6a :
		RG_rl_48_t1 = TR_60 ;
	7'h6b :
		RG_rl_48_t1 = TR_60 ;
	7'h6c :
		RG_rl_48_t1 = TR_60 ;
	7'h6d :
		RG_rl_48_t1 = TR_60 ;
	7'h6e :
		RG_rl_48_t1 = TR_60 ;
	7'h6f :
		RG_rl_48_t1 = TR_60 ;
	7'h70 :
		RG_rl_48_t1 = TR_60 ;
	7'h71 :
		RG_rl_48_t1 = TR_60 ;
	7'h72 :
		RG_rl_48_t1 = TR_60 ;
	7'h73 :
		RG_rl_48_t1 = TR_60 ;
	7'h74 :
		RG_rl_48_t1 = TR_60 ;
	7'h75 :
		RG_rl_48_t1 = TR_60 ;
	7'h76 :
		RG_rl_48_t1 = TR_60 ;
	7'h77 :
		RG_rl_48_t1 = TR_60 ;
	7'h78 :
		RG_rl_48_t1 = TR_60 ;
	7'h79 :
		RG_rl_48_t1 = TR_60 ;
	7'h7a :
		RG_rl_48_t1 = TR_60 ;
	7'h7b :
		RG_rl_48_t1 = TR_60 ;
	7'h7c :
		RG_rl_48_t1 = TR_60 ;
	7'h7d :
		RG_rl_48_t1 = TR_60 ;
	7'h7e :
		RG_rl_48_t1 = TR_60 ;
	7'h7f :
		RG_rl_48_t1 = TR_60 ;
	default :
		RG_rl_48_t1 = 9'hx ;
	endcase
always @ ( RG_rl_48_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_231 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_48_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h30 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_48_t = ( ( { 9{ U_570 } } & RG_rl_231 )
		| ( { 9{ U_569 } } & RG_rl_48_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_48_en = ( U_570 | RG_rl_48_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_48_en )
		RG_rl_48 <= RG_rl_48_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_61 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_49_t1 = TR_61 ;
	7'h01 :
		RG_rl_49_t1 = TR_61 ;
	7'h02 :
		RG_rl_49_t1 = TR_61 ;
	7'h03 :
		RG_rl_49_t1 = TR_61 ;
	7'h04 :
		RG_rl_49_t1 = TR_61 ;
	7'h05 :
		RG_rl_49_t1 = TR_61 ;
	7'h06 :
		RG_rl_49_t1 = TR_61 ;
	7'h07 :
		RG_rl_49_t1 = TR_61 ;
	7'h08 :
		RG_rl_49_t1 = TR_61 ;
	7'h09 :
		RG_rl_49_t1 = TR_61 ;
	7'h0a :
		RG_rl_49_t1 = TR_61 ;
	7'h0b :
		RG_rl_49_t1 = TR_61 ;
	7'h0c :
		RG_rl_49_t1 = TR_61 ;
	7'h0d :
		RG_rl_49_t1 = TR_61 ;
	7'h0e :
		RG_rl_49_t1 = TR_61 ;
	7'h0f :
		RG_rl_49_t1 = TR_61 ;
	7'h10 :
		RG_rl_49_t1 = TR_61 ;
	7'h11 :
		RG_rl_49_t1 = TR_61 ;
	7'h12 :
		RG_rl_49_t1 = TR_61 ;
	7'h13 :
		RG_rl_49_t1 = TR_61 ;
	7'h14 :
		RG_rl_49_t1 = TR_61 ;
	7'h15 :
		RG_rl_49_t1 = TR_61 ;
	7'h16 :
		RG_rl_49_t1 = TR_61 ;
	7'h17 :
		RG_rl_49_t1 = TR_61 ;
	7'h18 :
		RG_rl_49_t1 = TR_61 ;
	7'h19 :
		RG_rl_49_t1 = TR_61 ;
	7'h1a :
		RG_rl_49_t1 = TR_61 ;
	7'h1b :
		RG_rl_49_t1 = TR_61 ;
	7'h1c :
		RG_rl_49_t1 = TR_61 ;
	7'h1d :
		RG_rl_49_t1 = TR_61 ;
	7'h1e :
		RG_rl_49_t1 = TR_61 ;
	7'h1f :
		RG_rl_49_t1 = TR_61 ;
	7'h20 :
		RG_rl_49_t1 = TR_61 ;
	7'h21 :
		RG_rl_49_t1 = TR_61 ;
	7'h22 :
		RG_rl_49_t1 = TR_61 ;
	7'h23 :
		RG_rl_49_t1 = TR_61 ;
	7'h24 :
		RG_rl_49_t1 = TR_61 ;
	7'h25 :
		RG_rl_49_t1 = TR_61 ;
	7'h26 :
		RG_rl_49_t1 = TR_61 ;
	7'h27 :
		RG_rl_49_t1 = TR_61 ;
	7'h28 :
		RG_rl_49_t1 = TR_61 ;
	7'h29 :
		RG_rl_49_t1 = TR_61 ;
	7'h2a :
		RG_rl_49_t1 = TR_61 ;
	7'h2b :
		RG_rl_49_t1 = TR_61 ;
	7'h2c :
		RG_rl_49_t1 = TR_61 ;
	7'h2d :
		RG_rl_49_t1 = TR_61 ;
	7'h2e :
		RG_rl_49_t1 = TR_61 ;
	7'h2f :
		RG_rl_49_t1 = TR_61 ;
	7'h30 :
		RG_rl_49_t1 = TR_61 ;
	7'h31 :
		RG_rl_49_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h32 :
		RG_rl_49_t1 = TR_61 ;
	7'h33 :
		RG_rl_49_t1 = TR_61 ;
	7'h34 :
		RG_rl_49_t1 = TR_61 ;
	7'h35 :
		RG_rl_49_t1 = TR_61 ;
	7'h36 :
		RG_rl_49_t1 = TR_61 ;
	7'h37 :
		RG_rl_49_t1 = TR_61 ;
	7'h38 :
		RG_rl_49_t1 = TR_61 ;
	7'h39 :
		RG_rl_49_t1 = TR_61 ;
	7'h3a :
		RG_rl_49_t1 = TR_61 ;
	7'h3b :
		RG_rl_49_t1 = TR_61 ;
	7'h3c :
		RG_rl_49_t1 = TR_61 ;
	7'h3d :
		RG_rl_49_t1 = TR_61 ;
	7'h3e :
		RG_rl_49_t1 = TR_61 ;
	7'h3f :
		RG_rl_49_t1 = TR_61 ;
	7'h40 :
		RG_rl_49_t1 = TR_61 ;
	7'h41 :
		RG_rl_49_t1 = TR_61 ;
	7'h42 :
		RG_rl_49_t1 = TR_61 ;
	7'h43 :
		RG_rl_49_t1 = TR_61 ;
	7'h44 :
		RG_rl_49_t1 = TR_61 ;
	7'h45 :
		RG_rl_49_t1 = TR_61 ;
	7'h46 :
		RG_rl_49_t1 = TR_61 ;
	7'h47 :
		RG_rl_49_t1 = TR_61 ;
	7'h48 :
		RG_rl_49_t1 = TR_61 ;
	7'h49 :
		RG_rl_49_t1 = TR_61 ;
	7'h4a :
		RG_rl_49_t1 = TR_61 ;
	7'h4b :
		RG_rl_49_t1 = TR_61 ;
	7'h4c :
		RG_rl_49_t1 = TR_61 ;
	7'h4d :
		RG_rl_49_t1 = TR_61 ;
	7'h4e :
		RG_rl_49_t1 = TR_61 ;
	7'h4f :
		RG_rl_49_t1 = TR_61 ;
	7'h50 :
		RG_rl_49_t1 = TR_61 ;
	7'h51 :
		RG_rl_49_t1 = TR_61 ;
	7'h52 :
		RG_rl_49_t1 = TR_61 ;
	7'h53 :
		RG_rl_49_t1 = TR_61 ;
	7'h54 :
		RG_rl_49_t1 = TR_61 ;
	7'h55 :
		RG_rl_49_t1 = TR_61 ;
	7'h56 :
		RG_rl_49_t1 = TR_61 ;
	7'h57 :
		RG_rl_49_t1 = TR_61 ;
	7'h58 :
		RG_rl_49_t1 = TR_61 ;
	7'h59 :
		RG_rl_49_t1 = TR_61 ;
	7'h5a :
		RG_rl_49_t1 = TR_61 ;
	7'h5b :
		RG_rl_49_t1 = TR_61 ;
	7'h5c :
		RG_rl_49_t1 = TR_61 ;
	7'h5d :
		RG_rl_49_t1 = TR_61 ;
	7'h5e :
		RG_rl_49_t1 = TR_61 ;
	7'h5f :
		RG_rl_49_t1 = TR_61 ;
	7'h60 :
		RG_rl_49_t1 = TR_61 ;
	7'h61 :
		RG_rl_49_t1 = TR_61 ;
	7'h62 :
		RG_rl_49_t1 = TR_61 ;
	7'h63 :
		RG_rl_49_t1 = TR_61 ;
	7'h64 :
		RG_rl_49_t1 = TR_61 ;
	7'h65 :
		RG_rl_49_t1 = TR_61 ;
	7'h66 :
		RG_rl_49_t1 = TR_61 ;
	7'h67 :
		RG_rl_49_t1 = TR_61 ;
	7'h68 :
		RG_rl_49_t1 = TR_61 ;
	7'h69 :
		RG_rl_49_t1 = TR_61 ;
	7'h6a :
		RG_rl_49_t1 = TR_61 ;
	7'h6b :
		RG_rl_49_t1 = TR_61 ;
	7'h6c :
		RG_rl_49_t1 = TR_61 ;
	7'h6d :
		RG_rl_49_t1 = TR_61 ;
	7'h6e :
		RG_rl_49_t1 = TR_61 ;
	7'h6f :
		RG_rl_49_t1 = TR_61 ;
	7'h70 :
		RG_rl_49_t1 = TR_61 ;
	7'h71 :
		RG_rl_49_t1 = TR_61 ;
	7'h72 :
		RG_rl_49_t1 = TR_61 ;
	7'h73 :
		RG_rl_49_t1 = TR_61 ;
	7'h74 :
		RG_rl_49_t1 = TR_61 ;
	7'h75 :
		RG_rl_49_t1 = TR_61 ;
	7'h76 :
		RG_rl_49_t1 = TR_61 ;
	7'h77 :
		RG_rl_49_t1 = TR_61 ;
	7'h78 :
		RG_rl_49_t1 = TR_61 ;
	7'h79 :
		RG_rl_49_t1 = TR_61 ;
	7'h7a :
		RG_rl_49_t1 = TR_61 ;
	7'h7b :
		RG_rl_49_t1 = TR_61 ;
	7'h7c :
		RG_rl_49_t1 = TR_61 ;
	7'h7d :
		RG_rl_49_t1 = TR_61 ;
	7'h7e :
		RG_rl_49_t1 = TR_61 ;
	7'h7f :
		RG_rl_49_t1 = TR_61 ;
	default :
		RG_rl_49_t1 = 9'hx ;
	endcase
always @ ( RG_rl_49_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_232 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_49_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h31 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_49_t = ( ( { 9{ U_570 } } & RG_rl_232 )
		| ( { 9{ U_569 } } & RG_rl_49_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_49_en = ( U_570 | RG_rl_49_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_49_en )
		RG_rl_49 <= RG_rl_49_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_62 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_50_t1 = TR_62 ;
	7'h01 :
		RG_rl_50_t1 = TR_62 ;
	7'h02 :
		RG_rl_50_t1 = TR_62 ;
	7'h03 :
		RG_rl_50_t1 = TR_62 ;
	7'h04 :
		RG_rl_50_t1 = TR_62 ;
	7'h05 :
		RG_rl_50_t1 = TR_62 ;
	7'h06 :
		RG_rl_50_t1 = TR_62 ;
	7'h07 :
		RG_rl_50_t1 = TR_62 ;
	7'h08 :
		RG_rl_50_t1 = TR_62 ;
	7'h09 :
		RG_rl_50_t1 = TR_62 ;
	7'h0a :
		RG_rl_50_t1 = TR_62 ;
	7'h0b :
		RG_rl_50_t1 = TR_62 ;
	7'h0c :
		RG_rl_50_t1 = TR_62 ;
	7'h0d :
		RG_rl_50_t1 = TR_62 ;
	7'h0e :
		RG_rl_50_t1 = TR_62 ;
	7'h0f :
		RG_rl_50_t1 = TR_62 ;
	7'h10 :
		RG_rl_50_t1 = TR_62 ;
	7'h11 :
		RG_rl_50_t1 = TR_62 ;
	7'h12 :
		RG_rl_50_t1 = TR_62 ;
	7'h13 :
		RG_rl_50_t1 = TR_62 ;
	7'h14 :
		RG_rl_50_t1 = TR_62 ;
	7'h15 :
		RG_rl_50_t1 = TR_62 ;
	7'h16 :
		RG_rl_50_t1 = TR_62 ;
	7'h17 :
		RG_rl_50_t1 = TR_62 ;
	7'h18 :
		RG_rl_50_t1 = TR_62 ;
	7'h19 :
		RG_rl_50_t1 = TR_62 ;
	7'h1a :
		RG_rl_50_t1 = TR_62 ;
	7'h1b :
		RG_rl_50_t1 = TR_62 ;
	7'h1c :
		RG_rl_50_t1 = TR_62 ;
	7'h1d :
		RG_rl_50_t1 = TR_62 ;
	7'h1e :
		RG_rl_50_t1 = TR_62 ;
	7'h1f :
		RG_rl_50_t1 = TR_62 ;
	7'h20 :
		RG_rl_50_t1 = TR_62 ;
	7'h21 :
		RG_rl_50_t1 = TR_62 ;
	7'h22 :
		RG_rl_50_t1 = TR_62 ;
	7'h23 :
		RG_rl_50_t1 = TR_62 ;
	7'h24 :
		RG_rl_50_t1 = TR_62 ;
	7'h25 :
		RG_rl_50_t1 = TR_62 ;
	7'h26 :
		RG_rl_50_t1 = TR_62 ;
	7'h27 :
		RG_rl_50_t1 = TR_62 ;
	7'h28 :
		RG_rl_50_t1 = TR_62 ;
	7'h29 :
		RG_rl_50_t1 = TR_62 ;
	7'h2a :
		RG_rl_50_t1 = TR_62 ;
	7'h2b :
		RG_rl_50_t1 = TR_62 ;
	7'h2c :
		RG_rl_50_t1 = TR_62 ;
	7'h2d :
		RG_rl_50_t1 = TR_62 ;
	7'h2e :
		RG_rl_50_t1 = TR_62 ;
	7'h2f :
		RG_rl_50_t1 = TR_62 ;
	7'h30 :
		RG_rl_50_t1 = TR_62 ;
	7'h31 :
		RG_rl_50_t1 = TR_62 ;
	7'h32 :
		RG_rl_50_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h33 :
		RG_rl_50_t1 = TR_62 ;
	7'h34 :
		RG_rl_50_t1 = TR_62 ;
	7'h35 :
		RG_rl_50_t1 = TR_62 ;
	7'h36 :
		RG_rl_50_t1 = TR_62 ;
	7'h37 :
		RG_rl_50_t1 = TR_62 ;
	7'h38 :
		RG_rl_50_t1 = TR_62 ;
	7'h39 :
		RG_rl_50_t1 = TR_62 ;
	7'h3a :
		RG_rl_50_t1 = TR_62 ;
	7'h3b :
		RG_rl_50_t1 = TR_62 ;
	7'h3c :
		RG_rl_50_t1 = TR_62 ;
	7'h3d :
		RG_rl_50_t1 = TR_62 ;
	7'h3e :
		RG_rl_50_t1 = TR_62 ;
	7'h3f :
		RG_rl_50_t1 = TR_62 ;
	7'h40 :
		RG_rl_50_t1 = TR_62 ;
	7'h41 :
		RG_rl_50_t1 = TR_62 ;
	7'h42 :
		RG_rl_50_t1 = TR_62 ;
	7'h43 :
		RG_rl_50_t1 = TR_62 ;
	7'h44 :
		RG_rl_50_t1 = TR_62 ;
	7'h45 :
		RG_rl_50_t1 = TR_62 ;
	7'h46 :
		RG_rl_50_t1 = TR_62 ;
	7'h47 :
		RG_rl_50_t1 = TR_62 ;
	7'h48 :
		RG_rl_50_t1 = TR_62 ;
	7'h49 :
		RG_rl_50_t1 = TR_62 ;
	7'h4a :
		RG_rl_50_t1 = TR_62 ;
	7'h4b :
		RG_rl_50_t1 = TR_62 ;
	7'h4c :
		RG_rl_50_t1 = TR_62 ;
	7'h4d :
		RG_rl_50_t1 = TR_62 ;
	7'h4e :
		RG_rl_50_t1 = TR_62 ;
	7'h4f :
		RG_rl_50_t1 = TR_62 ;
	7'h50 :
		RG_rl_50_t1 = TR_62 ;
	7'h51 :
		RG_rl_50_t1 = TR_62 ;
	7'h52 :
		RG_rl_50_t1 = TR_62 ;
	7'h53 :
		RG_rl_50_t1 = TR_62 ;
	7'h54 :
		RG_rl_50_t1 = TR_62 ;
	7'h55 :
		RG_rl_50_t1 = TR_62 ;
	7'h56 :
		RG_rl_50_t1 = TR_62 ;
	7'h57 :
		RG_rl_50_t1 = TR_62 ;
	7'h58 :
		RG_rl_50_t1 = TR_62 ;
	7'h59 :
		RG_rl_50_t1 = TR_62 ;
	7'h5a :
		RG_rl_50_t1 = TR_62 ;
	7'h5b :
		RG_rl_50_t1 = TR_62 ;
	7'h5c :
		RG_rl_50_t1 = TR_62 ;
	7'h5d :
		RG_rl_50_t1 = TR_62 ;
	7'h5e :
		RG_rl_50_t1 = TR_62 ;
	7'h5f :
		RG_rl_50_t1 = TR_62 ;
	7'h60 :
		RG_rl_50_t1 = TR_62 ;
	7'h61 :
		RG_rl_50_t1 = TR_62 ;
	7'h62 :
		RG_rl_50_t1 = TR_62 ;
	7'h63 :
		RG_rl_50_t1 = TR_62 ;
	7'h64 :
		RG_rl_50_t1 = TR_62 ;
	7'h65 :
		RG_rl_50_t1 = TR_62 ;
	7'h66 :
		RG_rl_50_t1 = TR_62 ;
	7'h67 :
		RG_rl_50_t1 = TR_62 ;
	7'h68 :
		RG_rl_50_t1 = TR_62 ;
	7'h69 :
		RG_rl_50_t1 = TR_62 ;
	7'h6a :
		RG_rl_50_t1 = TR_62 ;
	7'h6b :
		RG_rl_50_t1 = TR_62 ;
	7'h6c :
		RG_rl_50_t1 = TR_62 ;
	7'h6d :
		RG_rl_50_t1 = TR_62 ;
	7'h6e :
		RG_rl_50_t1 = TR_62 ;
	7'h6f :
		RG_rl_50_t1 = TR_62 ;
	7'h70 :
		RG_rl_50_t1 = TR_62 ;
	7'h71 :
		RG_rl_50_t1 = TR_62 ;
	7'h72 :
		RG_rl_50_t1 = TR_62 ;
	7'h73 :
		RG_rl_50_t1 = TR_62 ;
	7'h74 :
		RG_rl_50_t1 = TR_62 ;
	7'h75 :
		RG_rl_50_t1 = TR_62 ;
	7'h76 :
		RG_rl_50_t1 = TR_62 ;
	7'h77 :
		RG_rl_50_t1 = TR_62 ;
	7'h78 :
		RG_rl_50_t1 = TR_62 ;
	7'h79 :
		RG_rl_50_t1 = TR_62 ;
	7'h7a :
		RG_rl_50_t1 = TR_62 ;
	7'h7b :
		RG_rl_50_t1 = TR_62 ;
	7'h7c :
		RG_rl_50_t1 = TR_62 ;
	7'h7d :
		RG_rl_50_t1 = TR_62 ;
	7'h7e :
		RG_rl_50_t1 = TR_62 ;
	7'h7f :
		RG_rl_50_t1 = TR_62 ;
	default :
		RG_rl_50_t1 = 9'hx ;
	endcase
always @ ( RG_rl_50_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_233 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_50_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h32 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_50_t = ( ( { 9{ U_570 } } & RG_rl_233 )
		| ( { 9{ U_569 } } & RG_rl_50_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_50_en = ( U_570 | RG_rl_50_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_50_en )
		RG_rl_50 <= RG_rl_50_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_63 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_51_t1 = TR_63 ;
	7'h01 :
		RG_rl_51_t1 = TR_63 ;
	7'h02 :
		RG_rl_51_t1 = TR_63 ;
	7'h03 :
		RG_rl_51_t1 = TR_63 ;
	7'h04 :
		RG_rl_51_t1 = TR_63 ;
	7'h05 :
		RG_rl_51_t1 = TR_63 ;
	7'h06 :
		RG_rl_51_t1 = TR_63 ;
	7'h07 :
		RG_rl_51_t1 = TR_63 ;
	7'h08 :
		RG_rl_51_t1 = TR_63 ;
	7'h09 :
		RG_rl_51_t1 = TR_63 ;
	7'h0a :
		RG_rl_51_t1 = TR_63 ;
	7'h0b :
		RG_rl_51_t1 = TR_63 ;
	7'h0c :
		RG_rl_51_t1 = TR_63 ;
	7'h0d :
		RG_rl_51_t1 = TR_63 ;
	7'h0e :
		RG_rl_51_t1 = TR_63 ;
	7'h0f :
		RG_rl_51_t1 = TR_63 ;
	7'h10 :
		RG_rl_51_t1 = TR_63 ;
	7'h11 :
		RG_rl_51_t1 = TR_63 ;
	7'h12 :
		RG_rl_51_t1 = TR_63 ;
	7'h13 :
		RG_rl_51_t1 = TR_63 ;
	7'h14 :
		RG_rl_51_t1 = TR_63 ;
	7'h15 :
		RG_rl_51_t1 = TR_63 ;
	7'h16 :
		RG_rl_51_t1 = TR_63 ;
	7'h17 :
		RG_rl_51_t1 = TR_63 ;
	7'h18 :
		RG_rl_51_t1 = TR_63 ;
	7'h19 :
		RG_rl_51_t1 = TR_63 ;
	7'h1a :
		RG_rl_51_t1 = TR_63 ;
	7'h1b :
		RG_rl_51_t1 = TR_63 ;
	7'h1c :
		RG_rl_51_t1 = TR_63 ;
	7'h1d :
		RG_rl_51_t1 = TR_63 ;
	7'h1e :
		RG_rl_51_t1 = TR_63 ;
	7'h1f :
		RG_rl_51_t1 = TR_63 ;
	7'h20 :
		RG_rl_51_t1 = TR_63 ;
	7'h21 :
		RG_rl_51_t1 = TR_63 ;
	7'h22 :
		RG_rl_51_t1 = TR_63 ;
	7'h23 :
		RG_rl_51_t1 = TR_63 ;
	7'h24 :
		RG_rl_51_t1 = TR_63 ;
	7'h25 :
		RG_rl_51_t1 = TR_63 ;
	7'h26 :
		RG_rl_51_t1 = TR_63 ;
	7'h27 :
		RG_rl_51_t1 = TR_63 ;
	7'h28 :
		RG_rl_51_t1 = TR_63 ;
	7'h29 :
		RG_rl_51_t1 = TR_63 ;
	7'h2a :
		RG_rl_51_t1 = TR_63 ;
	7'h2b :
		RG_rl_51_t1 = TR_63 ;
	7'h2c :
		RG_rl_51_t1 = TR_63 ;
	7'h2d :
		RG_rl_51_t1 = TR_63 ;
	7'h2e :
		RG_rl_51_t1 = TR_63 ;
	7'h2f :
		RG_rl_51_t1 = TR_63 ;
	7'h30 :
		RG_rl_51_t1 = TR_63 ;
	7'h31 :
		RG_rl_51_t1 = TR_63 ;
	7'h32 :
		RG_rl_51_t1 = TR_63 ;
	7'h33 :
		RG_rl_51_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h34 :
		RG_rl_51_t1 = TR_63 ;
	7'h35 :
		RG_rl_51_t1 = TR_63 ;
	7'h36 :
		RG_rl_51_t1 = TR_63 ;
	7'h37 :
		RG_rl_51_t1 = TR_63 ;
	7'h38 :
		RG_rl_51_t1 = TR_63 ;
	7'h39 :
		RG_rl_51_t1 = TR_63 ;
	7'h3a :
		RG_rl_51_t1 = TR_63 ;
	7'h3b :
		RG_rl_51_t1 = TR_63 ;
	7'h3c :
		RG_rl_51_t1 = TR_63 ;
	7'h3d :
		RG_rl_51_t1 = TR_63 ;
	7'h3e :
		RG_rl_51_t1 = TR_63 ;
	7'h3f :
		RG_rl_51_t1 = TR_63 ;
	7'h40 :
		RG_rl_51_t1 = TR_63 ;
	7'h41 :
		RG_rl_51_t1 = TR_63 ;
	7'h42 :
		RG_rl_51_t1 = TR_63 ;
	7'h43 :
		RG_rl_51_t1 = TR_63 ;
	7'h44 :
		RG_rl_51_t1 = TR_63 ;
	7'h45 :
		RG_rl_51_t1 = TR_63 ;
	7'h46 :
		RG_rl_51_t1 = TR_63 ;
	7'h47 :
		RG_rl_51_t1 = TR_63 ;
	7'h48 :
		RG_rl_51_t1 = TR_63 ;
	7'h49 :
		RG_rl_51_t1 = TR_63 ;
	7'h4a :
		RG_rl_51_t1 = TR_63 ;
	7'h4b :
		RG_rl_51_t1 = TR_63 ;
	7'h4c :
		RG_rl_51_t1 = TR_63 ;
	7'h4d :
		RG_rl_51_t1 = TR_63 ;
	7'h4e :
		RG_rl_51_t1 = TR_63 ;
	7'h4f :
		RG_rl_51_t1 = TR_63 ;
	7'h50 :
		RG_rl_51_t1 = TR_63 ;
	7'h51 :
		RG_rl_51_t1 = TR_63 ;
	7'h52 :
		RG_rl_51_t1 = TR_63 ;
	7'h53 :
		RG_rl_51_t1 = TR_63 ;
	7'h54 :
		RG_rl_51_t1 = TR_63 ;
	7'h55 :
		RG_rl_51_t1 = TR_63 ;
	7'h56 :
		RG_rl_51_t1 = TR_63 ;
	7'h57 :
		RG_rl_51_t1 = TR_63 ;
	7'h58 :
		RG_rl_51_t1 = TR_63 ;
	7'h59 :
		RG_rl_51_t1 = TR_63 ;
	7'h5a :
		RG_rl_51_t1 = TR_63 ;
	7'h5b :
		RG_rl_51_t1 = TR_63 ;
	7'h5c :
		RG_rl_51_t1 = TR_63 ;
	7'h5d :
		RG_rl_51_t1 = TR_63 ;
	7'h5e :
		RG_rl_51_t1 = TR_63 ;
	7'h5f :
		RG_rl_51_t1 = TR_63 ;
	7'h60 :
		RG_rl_51_t1 = TR_63 ;
	7'h61 :
		RG_rl_51_t1 = TR_63 ;
	7'h62 :
		RG_rl_51_t1 = TR_63 ;
	7'h63 :
		RG_rl_51_t1 = TR_63 ;
	7'h64 :
		RG_rl_51_t1 = TR_63 ;
	7'h65 :
		RG_rl_51_t1 = TR_63 ;
	7'h66 :
		RG_rl_51_t1 = TR_63 ;
	7'h67 :
		RG_rl_51_t1 = TR_63 ;
	7'h68 :
		RG_rl_51_t1 = TR_63 ;
	7'h69 :
		RG_rl_51_t1 = TR_63 ;
	7'h6a :
		RG_rl_51_t1 = TR_63 ;
	7'h6b :
		RG_rl_51_t1 = TR_63 ;
	7'h6c :
		RG_rl_51_t1 = TR_63 ;
	7'h6d :
		RG_rl_51_t1 = TR_63 ;
	7'h6e :
		RG_rl_51_t1 = TR_63 ;
	7'h6f :
		RG_rl_51_t1 = TR_63 ;
	7'h70 :
		RG_rl_51_t1 = TR_63 ;
	7'h71 :
		RG_rl_51_t1 = TR_63 ;
	7'h72 :
		RG_rl_51_t1 = TR_63 ;
	7'h73 :
		RG_rl_51_t1 = TR_63 ;
	7'h74 :
		RG_rl_51_t1 = TR_63 ;
	7'h75 :
		RG_rl_51_t1 = TR_63 ;
	7'h76 :
		RG_rl_51_t1 = TR_63 ;
	7'h77 :
		RG_rl_51_t1 = TR_63 ;
	7'h78 :
		RG_rl_51_t1 = TR_63 ;
	7'h79 :
		RG_rl_51_t1 = TR_63 ;
	7'h7a :
		RG_rl_51_t1 = TR_63 ;
	7'h7b :
		RG_rl_51_t1 = TR_63 ;
	7'h7c :
		RG_rl_51_t1 = TR_63 ;
	7'h7d :
		RG_rl_51_t1 = TR_63 ;
	7'h7e :
		RG_rl_51_t1 = TR_63 ;
	7'h7f :
		RG_rl_51_t1 = TR_63 ;
	default :
		RG_rl_51_t1 = 9'hx ;
	endcase
always @ ( RG_rl_51_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_234 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_51_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h33 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_51_t = ( ( { 9{ U_570 } } & RG_rl_234 )
		| ( { 9{ U_569 } } & RG_rl_51_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_51_en = ( U_570 | RG_rl_51_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_51_en )
		RG_rl_51 <= RG_rl_51_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_64 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_52_t1 = TR_64 ;
	7'h01 :
		RG_rl_52_t1 = TR_64 ;
	7'h02 :
		RG_rl_52_t1 = TR_64 ;
	7'h03 :
		RG_rl_52_t1 = TR_64 ;
	7'h04 :
		RG_rl_52_t1 = TR_64 ;
	7'h05 :
		RG_rl_52_t1 = TR_64 ;
	7'h06 :
		RG_rl_52_t1 = TR_64 ;
	7'h07 :
		RG_rl_52_t1 = TR_64 ;
	7'h08 :
		RG_rl_52_t1 = TR_64 ;
	7'h09 :
		RG_rl_52_t1 = TR_64 ;
	7'h0a :
		RG_rl_52_t1 = TR_64 ;
	7'h0b :
		RG_rl_52_t1 = TR_64 ;
	7'h0c :
		RG_rl_52_t1 = TR_64 ;
	7'h0d :
		RG_rl_52_t1 = TR_64 ;
	7'h0e :
		RG_rl_52_t1 = TR_64 ;
	7'h0f :
		RG_rl_52_t1 = TR_64 ;
	7'h10 :
		RG_rl_52_t1 = TR_64 ;
	7'h11 :
		RG_rl_52_t1 = TR_64 ;
	7'h12 :
		RG_rl_52_t1 = TR_64 ;
	7'h13 :
		RG_rl_52_t1 = TR_64 ;
	7'h14 :
		RG_rl_52_t1 = TR_64 ;
	7'h15 :
		RG_rl_52_t1 = TR_64 ;
	7'h16 :
		RG_rl_52_t1 = TR_64 ;
	7'h17 :
		RG_rl_52_t1 = TR_64 ;
	7'h18 :
		RG_rl_52_t1 = TR_64 ;
	7'h19 :
		RG_rl_52_t1 = TR_64 ;
	7'h1a :
		RG_rl_52_t1 = TR_64 ;
	7'h1b :
		RG_rl_52_t1 = TR_64 ;
	7'h1c :
		RG_rl_52_t1 = TR_64 ;
	7'h1d :
		RG_rl_52_t1 = TR_64 ;
	7'h1e :
		RG_rl_52_t1 = TR_64 ;
	7'h1f :
		RG_rl_52_t1 = TR_64 ;
	7'h20 :
		RG_rl_52_t1 = TR_64 ;
	7'h21 :
		RG_rl_52_t1 = TR_64 ;
	7'h22 :
		RG_rl_52_t1 = TR_64 ;
	7'h23 :
		RG_rl_52_t1 = TR_64 ;
	7'h24 :
		RG_rl_52_t1 = TR_64 ;
	7'h25 :
		RG_rl_52_t1 = TR_64 ;
	7'h26 :
		RG_rl_52_t1 = TR_64 ;
	7'h27 :
		RG_rl_52_t1 = TR_64 ;
	7'h28 :
		RG_rl_52_t1 = TR_64 ;
	7'h29 :
		RG_rl_52_t1 = TR_64 ;
	7'h2a :
		RG_rl_52_t1 = TR_64 ;
	7'h2b :
		RG_rl_52_t1 = TR_64 ;
	7'h2c :
		RG_rl_52_t1 = TR_64 ;
	7'h2d :
		RG_rl_52_t1 = TR_64 ;
	7'h2e :
		RG_rl_52_t1 = TR_64 ;
	7'h2f :
		RG_rl_52_t1 = TR_64 ;
	7'h30 :
		RG_rl_52_t1 = TR_64 ;
	7'h31 :
		RG_rl_52_t1 = TR_64 ;
	7'h32 :
		RG_rl_52_t1 = TR_64 ;
	7'h33 :
		RG_rl_52_t1 = TR_64 ;
	7'h34 :
		RG_rl_52_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h35 :
		RG_rl_52_t1 = TR_64 ;
	7'h36 :
		RG_rl_52_t1 = TR_64 ;
	7'h37 :
		RG_rl_52_t1 = TR_64 ;
	7'h38 :
		RG_rl_52_t1 = TR_64 ;
	7'h39 :
		RG_rl_52_t1 = TR_64 ;
	7'h3a :
		RG_rl_52_t1 = TR_64 ;
	7'h3b :
		RG_rl_52_t1 = TR_64 ;
	7'h3c :
		RG_rl_52_t1 = TR_64 ;
	7'h3d :
		RG_rl_52_t1 = TR_64 ;
	7'h3e :
		RG_rl_52_t1 = TR_64 ;
	7'h3f :
		RG_rl_52_t1 = TR_64 ;
	7'h40 :
		RG_rl_52_t1 = TR_64 ;
	7'h41 :
		RG_rl_52_t1 = TR_64 ;
	7'h42 :
		RG_rl_52_t1 = TR_64 ;
	7'h43 :
		RG_rl_52_t1 = TR_64 ;
	7'h44 :
		RG_rl_52_t1 = TR_64 ;
	7'h45 :
		RG_rl_52_t1 = TR_64 ;
	7'h46 :
		RG_rl_52_t1 = TR_64 ;
	7'h47 :
		RG_rl_52_t1 = TR_64 ;
	7'h48 :
		RG_rl_52_t1 = TR_64 ;
	7'h49 :
		RG_rl_52_t1 = TR_64 ;
	7'h4a :
		RG_rl_52_t1 = TR_64 ;
	7'h4b :
		RG_rl_52_t1 = TR_64 ;
	7'h4c :
		RG_rl_52_t1 = TR_64 ;
	7'h4d :
		RG_rl_52_t1 = TR_64 ;
	7'h4e :
		RG_rl_52_t1 = TR_64 ;
	7'h4f :
		RG_rl_52_t1 = TR_64 ;
	7'h50 :
		RG_rl_52_t1 = TR_64 ;
	7'h51 :
		RG_rl_52_t1 = TR_64 ;
	7'h52 :
		RG_rl_52_t1 = TR_64 ;
	7'h53 :
		RG_rl_52_t1 = TR_64 ;
	7'h54 :
		RG_rl_52_t1 = TR_64 ;
	7'h55 :
		RG_rl_52_t1 = TR_64 ;
	7'h56 :
		RG_rl_52_t1 = TR_64 ;
	7'h57 :
		RG_rl_52_t1 = TR_64 ;
	7'h58 :
		RG_rl_52_t1 = TR_64 ;
	7'h59 :
		RG_rl_52_t1 = TR_64 ;
	7'h5a :
		RG_rl_52_t1 = TR_64 ;
	7'h5b :
		RG_rl_52_t1 = TR_64 ;
	7'h5c :
		RG_rl_52_t1 = TR_64 ;
	7'h5d :
		RG_rl_52_t1 = TR_64 ;
	7'h5e :
		RG_rl_52_t1 = TR_64 ;
	7'h5f :
		RG_rl_52_t1 = TR_64 ;
	7'h60 :
		RG_rl_52_t1 = TR_64 ;
	7'h61 :
		RG_rl_52_t1 = TR_64 ;
	7'h62 :
		RG_rl_52_t1 = TR_64 ;
	7'h63 :
		RG_rl_52_t1 = TR_64 ;
	7'h64 :
		RG_rl_52_t1 = TR_64 ;
	7'h65 :
		RG_rl_52_t1 = TR_64 ;
	7'h66 :
		RG_rl_52_t1 = TR_64 ;
	7'h67 :
		RG_rl_52_t1 = TR_64 ;
	7'h68 :
		RG_rl_52_t1 = TR_64 ;
	7'h69 :
		RG_rl_52_t1 = TR_64 ;
	7'h6a :
		RG_rl_52_t1 = TR_64 ;
	7'h6b :
		RG_rl_52_t1 = TR_64 ;
	7'h6c :
		RG_rl_52_t1 = TR_64 ;
	7'h6d :
		RG_rl_52_t1 = TR_64 ;
	7'h6e :
		RG_rl_52_t1 = TR_64 ;
	7'h6f :
		RG_rl_52_t1 = TR_64 ;
	7'h70 :
		RG_rl_52_t1 = TR_64 ;
	7'h71 :
		RG_rl_52_t1 = TR_64 ;
	7'h72 :
		RG_rl_52_t1 = TR_64 ;
	7'h73 :
		RG_rl_52_t1 = TR_64 ;
	7'h74 :
		RG_rl_52_t1 = TR_64 ;
	7'h75 :
		RG_rl_52_t1 = TR_64 ;
	7'h76 :
		RG_rl_52_t1 = TR_64 ;
	7'h77 :
		RG_rl_52_t1 = TR_64 ;
	7'h78 :
		RG_rl_52_t1 = TR_64 ;
	7'h79 :
		RG_rl_52_t1 = TR_64 ;
	7'h7a :
		RG_rl_52_t1 = TR_64 ;
	7'h7b :
		RG_rl_52_t1 = TR_64 ;
	7'h7c :
		RG_rl_52_t1 = TR_64 ;
	7'h7d :
		RG_rl_52_t1 = TR_64 ;
	7'h7e :
		RG_rl_52_t1 = TR_64 ;
	7'h7f :
		RG_rl_52_t1 = TR_64 ;
	default :
		RG_rl_52_t1 = 9'hx ;
	endcase
always @ ( RG_rl_52_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_235 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_52_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h34 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_52_t = ( ( { 9{ U_570 } } & RG_rl_235 )
		| ( { 9{ U_569 } } & RG_rl_52_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_52_en = ( U_570 | RG_rl_52_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_52_en )
		RG_rl_52 <= RG_rl_52_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_65 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_53_t1 = TR_65 ;
	7'h01 :
		RG_rl_53_t1 = TR_65 ;
	7'h02 :
		RG_rl_53_t1 = TR_65 ;
	7'h03 :
		RG_rl_53_t1 = TR_65 ;
	7'h04 :
		RG_rl_53_t1 = TR_65 ;
	7'h05 :
		RG_rl_53_t1 = TR_65 ;
	7'h06 :
		RG_rl_53_t1 = TR_65 ;
	7'h07 :
		RG_rl_53_t1 = TR_65 ;
	7'h08 :
		RG_rl_53_t1 = TR_65 ;
	7'h09 :
		RG_rl_53_t1 = TR_65 ;
	7'h0a :
		RG_rl_53_t1 = TR_65 ;
	7'h0b :
		RG_rl_53_t1 = TR_65 ;
	7'h0c :
		RG_rl_53_t1 = TR_65 ;
	7'h0d :
		RG_rl_53_t1 = TR_65 ;
	7'h0e :
		RG_rl_53_t1 = TR_65 ;
	7'h0f :
		RG_rl_53_t1 = TR_65 ;
	7'h10 :
		RG_rl_53_t1 = TR_65 ;
	7'h11 :
		RG_rl_53_t1 = TR_65 ;
	7'h12 :
		RG_rl_53_t1 = TR_65 ;
	7'h13 :
		RG_rl_53_t1 = TR_65 ;
	7'h14 :
		RG_rl_53_t1 = TR_65 ;
	7'h15 :
		RG_rl_53_t1 = TR_65 ;
	7'h16 :
		RG_rl_53_t1 = TR_65 ;
	7'h17 :
		RG_rl_53_t1 = TR_65 ;
	7'h18 :
		RG_rl_53_t1 = TR_65 ;
	7'h19 :
		RG_rl_53_t1 = TR_65 ;
	7'h1a :
		RG_rl_53_t1 = TR_65 ;
	7'h1b :
		RG_rl_53_t1 = TR_65 ;
	7'h1c :
		RG_rl_53_t1 = TR_65 ;
	7'h1d :
		RG_rl_53_t1 = TR_65 ;
	7'h1e :
		RG_rl_53_t1 = TR_65 ;
	7'h1f :
		RG_rl_53_t1 = TR_65 ;
	7'h20 :
		RG_rl_53_t1 = TR_65 ;
	7'h21 :
		RG_rl_53_t1 = TR_65 ;
	7'h22 :
		RG_rl_53_t1 = TR_65 ;
	7'h23 :
		RG_rl_53_t1 = TR_65 ;
	7'h24 :
		RG_rl_53_t1 = TR_65 ;
	7'h25 :
		RG_rl_53_t1 = TR_65 ;
	7'h26 :
		RG_rl_53_t1 = TR_65 ;
	7'h27 :
		RG_rl_53_t1 = TR_65 ;
	7'h28 :
		RG_rl_53_t1 = TR_65 ;
	7'h29 :
		RG_rl_53_t1 = TR_65 ;
	7'h2a :
		RG_rl_53_t1 = TR_65 ;
	7'h2b :
		RG_rl_53_t1 = TR_65 ;
	7'h2c :
		RG_rl_53_t1 = TR_65 ;
	7'h2d :
		RG_rl_53_t1 = TR_65 ;
	7'h2e :
		RG_rl_53_t1 = TR_65 ;
	7'h2f :
		RG_rl_53_t1 = TR_65 ;
	7'h30 :
		RG_rl_53_t1 = TR_65 ;
	7'h31 :
		RG_rl_53_t1 = TR_65 ;
	7'h32 :
		RG_rl_53_t1 = TR_65 ;
	7'h33 :
		RG_rl_53_t1 = TR_65 ;
	7'h34 :
		RG_rl_53_t1 = TR_65 ;
	7'h35 :
		RG_rl_53_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h36 :
		RG_rl_53_t1 = TR_65 ;
	7'h37 :
		RG_rl_53_t1 = TR_65 ;
	7'h38 :
		RG_rl_53_t1 = TR_65 ;
	7'h39 :
		RG_rl_53_t1 = TR_65 ;
	7'h3a :
		RG_rl_53_t1 = TR_65 ;
	7'h3b :
		RG_rl_53_t1 = TR_65 ;
	7'h3c :
		RG_rl_53_t1 = TR_65 ;
	7'h3d :
		RG_rl_53_t1 = TR_65 ;
	7'h3e :
		RG_rl_53_t1 = TR_65 ;
	7'h3f :
		RG_rl_53_t1 = TR_65 ;
	7'h40 :
		RG_rl_53_t1 = TR_65 ;
	7'h41 :
		RG_rl_53_t1 = TR_65 ;
	7'h42 :
		RG_rl_53_t1 = TR_65 ;
	7'h43 :
		RG_rl_53_t1 = TR_65 ;
	7'h44 :
		RG_rl_53_t1 = TR_65 ;
	7'h45 :
		RG_rl_53_t1 = TR_65 ;
	7'h46 :
		RG_rl_53_t1 = TR_65 ;
	7'h47 :
		RG_rl_53_t1 = TR_65 ;
	7'h48 :
		RG_rl_53_t1 = TR_65 ;
	7'h49 :
		RG_rl_53_t1 = TR_65 ;
	7'h4a :
		RG_rl_53_t1 = TR_65 ;
	7'h4b :
		RG_rl_53_t1 = TR_65 ;
	7'h4c :
		RG_rl_53_t1 = TR_65 ;
	7'h4d :
		RG_rl_53_t1 = TR_65 ;
	7'h4e :
		RG_rl_53_t1 = TR_65 ;
	7'h4f :
		RG_rl_53_t1 = TR_65 ;
	7'h50 :
		RG_rl_53_t1 = TR_65 ;
	7'h51 :
		RG_rl_53_t1 = TR_65 ;
	7'h52 :
		RG_rl_53_t1 = TR_65 ;
	7'h53 :
		RG_rl_53_t1 = TR_65 ;
	7'h54 :
		RG_rl_53_t1 = TR_65 ;
	7'h55 :
		RG_rl_53_t1 = TR_65 ;
	7'h56 :
		RG_rl_53_t1 = TR_65 ;
	7'h57 :
		RG_rl_53_t1 = TR_65 ;
	7'h58 :
		RG_rl_53_t1 = TR_65 ;
	7'h59 :
		RG_rl_53_t1 = TR_65 ;
	7'h5a :
		RG_rl_53_t1 = TR_65 ;
	7'h5b :
		RG_rl_53_t1 = TR_65 ;
	7'h5c :
		RG_rl_53_t1 = TR_65 ;
	7'h5d :
		RG_rl_53_t1 = TR_65 ;
	7'h5e :
		RG_rl_53_t1 = TR_65 ;
	7'h5f :
		RG_rl_53_t1 = TR_65 ;
	7'h60 :
		RG_rl_53_t1 = TR_65 ;
	7'h61 :
		RG_rl_53_t1 = TR_65 ;
	7'h62 :
		RG_rl_53_t1 = TR_65 ;
	7'h63 :
		RG_rl_53_t1 = TR_65 ;
	7'h64 :
		RG_rl_53_t1 = TR_65 ;
	7'h65 :
		RG_rl_53_t1 = TR_65 ;
	7'h66 :
		RG_rl_53_t1 = TR_65 ;
	7'h67 :
		RG_rl_53_t1 = TR_65 ;
	7'h68 :
		RG_rl_53_t1 = TR_65 ;
	7'h69 :
		RG_rl_53_t1 = TR_65 ;
	7'h6a :
		RG_rl_53_t1 = TR_65 ;
	7'h6b :
		RG_rl_53_t1 = TR_65 ;
	7'h6c :
		RG_rl_53_t1 = TR_65 ;
	7'h6d :
		RG_rl_53_t1 = TR_65 ;
	7'h6e :
		RG_rl_53_t1 = TR_65 ;
	7'h6f :
		RG_rl_53_t1 = TR_65 ;
	7'h70 :
		RG_rl_53_t1 = TR_65 ;
	7'h71 :
		RG_rl_53_t1 = TR_65 ;
	7'h72 :
		RG_rl_53_t1 = TR_65 ;
	7'h73 :
		RG_rl_53_t1 = TR_65 ;
	7'h74 :
		RG_rl_53_t1 = TR_65 ;
	7'h75 :
		RG_rl_53_t1 = TR_65 ;
	7'h76 :
		RG_rl_53_t1 = TR_65 ;
	7'h77 :
		RG_rl_53_t1 = TR_65 ;
	7'h78 :
		RG_rl_53_t1 = TR_65 ;
	7'h79 :
		RG_rl_53_t1 = TR_65 ;
	7'h7a :
		RG_rl_53_t1 = TR_65 ;
	7'h7b :
		RG_rl_53_t1 = TR_65 ;
	7'h7c :
		RG_rl_53_t1 = TR_65 ;
	7'h7d :
		RG_rl_53_t1 = TR_65 ;
	7'h7e :
		RG_rl_53_t1 = TR_65 ;
	7'h7f :
		RG_rl_53_t1 = TR_65 ;
	default :
		RG_rl_53_t1 = 9'hx ;
	endcase
always @ ( RG_rl_53_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_236 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_53_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h35 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_53_t = ( ( { 9{ U_570 } } & RG_rl_236 )
		| ( { 9{ U_569 } } & RG_rl_53_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_53_en = ( U_570 | RG_rl_53_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_53_en )
		RG_rl_53 <= RG_rl_53_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_66 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_54_t1 = TR_66 ;
	7'h01 :
		RG_rl_54_t1 = TR_66 ;
	7'h02 :
		RG_rl_54_t1 = TR_66 ;
	7'h03 :
		RG_rl_54_t1 = TR_66 ;
	7'h04 :
		RG_rl_54_t1 = TR_66 ;
	7'h05 :
		RG_rl_54_t1 = TR_66 ;
	7'h06 :
		RG_rl_54_t1 = TR_66 ;
	7'h07 :
		RG_rl_54_t1 = TR_66 ;
	7'h08 :
		RG_rl_54_t1 = TR_66 ;
	7'h09 :
		RG_rl_54_t1 = TR_66 ;
	7'h0a :
		RG_rl_54_t1 = TR_66 ;
	7'h0b :
		RG_rl_54_t1 = TR_66 ;
	7'h0c :
		RG_rl_54_t1 = TR_66 ;
	7'h0d :
		RG_rl_54_t1 = TR_66 ;
	7'h0e :
		RG_rl_54_t1 = TR_66 ;
	7'h0f :
		RG_rl_54_t1 = TR_66 ;
	7'h10 :
		RG_rl_54_t1 = TR_66 ;
	7'h11 :
		RG_rl_54_t1 = TR_66 ;
	7'h12 :
		RG_rl_54_t1 = TR_66 ;
	7'h13 :
		RG_rl_54_t1 = TR_66 ;
	7'h14 :
		RG_rl_54_t1 = TR_66 ;
	7'h15 :
		RG_rl_54_t1 = TR_66 ;
	7'h16 :
		RG_rl_54_t1 = TR_66 ;
	7'h17 :
		RG_rl_54_t1 = TR_66 ;
	7'h18 :
		RG_rl_54_t1 = TR_66 ;
	7'h19 :
		RG_rl_54_t1 = TR_66 ;
	7'h1a :
		RG_rl_54_t1 = TR_66 ;
	7'h1b :
		RG_rl_54_t1 = TR_66 ;
	7'h1c :
		RG_rl_54_t1 = TR_66 ;
	7'h1d :
		RG_rl_54_t1 = TR_66 ;
	7'h1e :
		RG_rl_54_t1 = TR_66 ;
	7'h1f :
		RG_rl_54_t1 = TR_66 ;
	7'h20 :
		RG_rl_54_t1 = TR_66 ;
	7'h21 :
		RG_rl_54_t1 = TR_66 ;
	7'h22 :
		RG_rl_54_t1 = TR_66 ;
	7'h23 :
		RG_rl_54_t1 = TR_66 ;
	7'h24 :
		RG_rl_54_t1 = TR_66 ;
	7'h25 :
		RG_rl_54_t1 = TR_66 ;
	7'h26 :
		RG_rl_54_t1 = TR_66 ;
	7'h27 :
		RG_rl_54_t1 = TR_66 ;
	7'h28 :
		RG_rl_54_t1 = TR_66 ;
	7'h29 :
		RG_rl_54_t1 = TR_66 ;
	7'h2a :
		RG_rl_54_t1 = TR_66 ;
	7'h2b :
		RG_rl_54_t1 = TR_66 ;
	7'h2c :
		RG_rl_54_t1 = TR_66 ;
	7'h2d :
		RG_rl_54_t1 = TR_66 ;
	7'h2e :
		RG_rl_54_t1 = TR_66 ;
	7'h2f :
		RG_rl_54_t1 = TR_66 ;
	7'h30 :
		RG_rl_54_t1 = TR_66 ;
	7'h31 :
		RG_rl_54_t1 = TR_66 ;
	7'h32 :
		RG_rl_54_t1 = TR_66 ;
	7'h33 :
		RG_rl_54_t1 = TR_66 ;
	7'h34 :
		RG_rl_54_t1 = TR_66 ;
	7'h35 :
		RG_rl_54_t1 = TR_66 ;
	7'h36 :
		RG_rl_54_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h37 :
		RG_rl_54_t1 = TR_66 ;
	7'h38 :
		RG_rl_54_t1 = TR_66 ;
	7'h39 :
		RG_rl_54_t1 = TR_66 ;
	7'h3a :
		RG_rl_54_t1 = TR_66 ;
	7'h3b :
		RG_rl_54_t1 = TR_66 ;
	7'h3c :
		RG_rl_54_t1 = TR_66 ;
	7'h3d :
		RG_rl_54_t1 = TR_66 ;
	7'h3e :
		RG_rl_54_t1 = TR_66 ;
	7'h3f :
		RG_rl_54_t1 = TR_66 ;
	7'h40 :
		RG_rl_54_t1 = TR_66 ;
	7'h41 :
		RG_rl_54_t1 = TR_66 ;
	7'h42 :
		RG_rl_54_t1 = TR_66 ;
	7'h43 :
		RG_rl_54_t1 = TR_66 ;
	7'h44 :
		RG_rl_54_t1 = TR_66 ;
	7'h45 :
		RG_rl_54_t1 = TR_66 ;
	7'h46 :
		RG_rl_54_t1 = TR_66 ;
	7'h47 :
		RG_rl_54_t1 = TR_66 ;
	7'h48 :
		RG_rl_54_t1 = TR_66 ;
	7'h49 :
		RG_rl_54_t1 = TR_66 ;
	7'h4a :
		RG_rl_54_t1 = TR_66 ;
	7'h4b :
		RG_rl_54_t1 = TR_66 ;
	7'h4c :
		RG_rl_54_t1 = TR_66 ;
	7'h4d :
		RG_rl_54_t1 = TR_66 ;
	7'h4e :
		RG_rl_54_t1 = TR_66 ;
	7'h4f :
		RG_rl_54_t1 = TR_66 ;
	7'h50 :
		RG_rl_54_t1 = TR_66 ;
	7'h51 :
		RG_rl_54_t1 = TR_66 ;
	7'h52 :
		RG_rl_54_t1 = TR_66 ;
	7'h53 :
		RG_rl_54_t1 = TR_66 ;
	7'h54 :
		RG_rl_54_t1 = TR_66 ;
	7'h55 :
		RG_rl_54_t1 = TR_66 ;
	7'h56 :
		RG_rl_54_t1 = TR_66 ;
	7'h57 :
		RG_rl_54_t1 = TR_66 ;
	7'h58 :
		RG_rl_54_t1 = TR_66 ;
	7'h59 :
		RG_rl_54_t1 = TR_66 ;
	7'h5a :
		RG_rl_54_t1 = TR_66 ;
	7'h5b :
		RG_rl_54_t1 = TR_66 ;
	7'h5c :
		RG_rl_54_t1 = TR_66 ;
	7'h5d :
		RG_rl_54_t1 = TR_66 ;
	7'h5e :
		RG_rl_54_t1 = TR_66 ;
	7'h5f :
		RG_rl_54_t1 = TR_66 ;
	7'h60 :
		RG_rl_54_t1 = TR_66 ;
	7'h61 :
		RG_rl_54_t1 = TR_66 ;
	7'h62 :
		RG_rl_54_t1 = TR_66 ;
	7'h63 :
		RG_rl_54_t1 = TR_66 ;
	7'h64 :
		RG_rl_54_t1 = TR_66 ;
	7'h65 :
		RG_rl_54_t1 = TR_66 ;
	7'h66 :
		RG_rl_54_t1 = TR_66 ;
	7'h67 :
		RG_rl_54_t1 = TR_66 ;
	7'h68 :
		RG_rl_54_t1 = TR_66 ;
	7'h69 :
		RG_rl_54_t1 = TR_66 ;
	7'h6a :
		RG_rl_54_t1 = TR_66 ;
	7'h6b :
		RG_rl_54_t1 = TR_66 ;
	7'h6c :
		RG_rl_54_t1 = TR_66 ;
	7'h6d :
		RG_rl_54_t1 = TR_66 ;
	7'h6e :
		RG_rl_54_t1 = TR_66 ;
	7'h6f :
		RG_rl_54_t1 = TR_66 ;
	7'h70 :
		RG_rl_54_t1 = TR_66 ;
	7'h71 :
		RG_rl_54_t1 = TR_66 ;
	7'h72 :
		RG_rl_54_t1 = TR_66 ;
	7'h73 :
		RG_rl_54_t1 = TR_66 ;
	7'h74 :
		RG_rl_54_t1 = TR_66 ;
	7'h75 :
		RG_rl_54_t1 = TR_66 ;
	7'h76 :
		RG_rl_54_t1 = TR_66 ;
	7'h77 :
		RG_rl_54_t1 = TR_66 ;
	7'h78 :
		RG_rl_54_t1 = TR_66 ;
	7'h79 :
		RG_rl_54_t1 = TR_66 ;
	7'h7a :
		RG_rl_54_t1 = TR_66 ;
	7'h7b :
		RG_rl_54_t1 = TR_66 ;
	7'h7c :
		RG_rl_54_t1 = TR_66 ;
	7'h7d :
		RG_rl_54_t1 = TR_66 ;
	7'h7e :
		RG_rl_54_t1 = TR_66 ;
	7'h7f :
		RG_rl_54_t1 = TR_66 ;
	default :
		RG_rl_54_t1 = 9'hx ;
	endcase
always @ ( RG_rl_54_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_237 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_54_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h36 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_54_t = ( ( { 9{ U_570 } } & RG_rl_237 )
		| ( { 9{ U_569 } } & RG_rl_54_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_54_en = ( U_570 | RG_rl_54_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_54_en )
		RG_rl_54 <= RG_rl_54_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_67 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_55_t1 = TR_67 ;
	7'h01 :
		RG_rl_55_t1 = TR_67 ;
	7'h02 :
		RG_rl_55_t1 = TR_67 ;
	7'h03 :
		RG_rl_55_t1 = TR_67 ;
	7'h04 :
		RG_rl_55_t1 = TR_67 ;
	7'h05 :
		RG_rl_55_t1 = TR_67 ;
	7'h06 :
		RG_rl_55_t1 = TR_67 ;
	7'h07 :
		RG_rl_55_t1 = TR_67 ;
	7'h08 :
		RG_rl_55_t1 = TR_67 ;
	7'h09 :
		RG_rl_55_t1 = TR_67 ;
	7'h0a :
		RG_rl_55_t1 = TR_67 ;
	7'h0b :
		RG_rl_55_t1 = TR_67 ;
	7'h0c :
		RG_rl_55_t1 = TR_67 ;
	7'h0d :
		RG_rl_55_t1 = TR_67 ;
	7'h0e :
		RG_rl_55_t1 = TR_67 ;
	7'h0f :
		RG_rl_55_t1 = TR_67 ;
	7'h10 :
		RG_rl_55_t1 = TR_67 ;
	7'h11 :
		RG_rl_55_t1 = TR_67 ;
	7'h12 :
		RG_rl_55_t1 = TR_67 ;
	7'h13 :
		RG_rl_55_t1 = TR_67 ;
	7'h14 :
		RG_rl_55_t1 = TR_67 ;
	7'h15 :
		RG_rl_55_t1 = TR_67 ;
	7'h16 :
		RG_rl_55_t1 = TR_67 ;
	7'h17 :
		RG_rl_55_t1 = TR_67 ;
	7'h18 :
		RG_rl_55_t1 = TR_67 ;
	7'h19 :
		RG_rl_55_t1 = TR_67 ;
	7'h1a :
		RG_rl_55_t1 = TR_67 ;
	7'h1b :
		RG_rl_55_t1 = TR_67 ;
	7'h1c :
		RG_rl_55_t1 = TR_67 ;
	7'h1d :
		RG_rl_55_t1 = TR_67 ;
	7'h1e :
		RG_rl_55_t1 = TR_67 ;
	7'h1f :
		RG_rl_55_t1 = TR_67 ;
	7'h20 :
		RG_rl_55_t1 = TR_67 ;
	7'h21 :
		RG_rl_55_t1 = TR_67 ;
	7'h22 :
		RG_rl_55_t1 = TR_67 ;
	7'h23 :
		RG_rl_55_t1 = TR_67 ;
	7'h24 :
		RG_rl_55_t1 = TR_67 ;
	7'h25 :
		RG_rl_55_t1 = TR_67 ;
	7'h26 :
		RG_rl_55_t1 = TR_67 ;
	7'h27 :
		RG_rl_55_t1 = TR_67 ;
	7'h28 :
		RG_rl_55_t1 = TR_67 ;
	7'h29 :
		RG_rl_55_t1 = TR_67 ;
	7'h2a :
		RG_rl_55_t1 = TR_67 ;
	7'h2b :
		RG_rl_55_t1 = TR_67 ;
	7'h2c :
		RG_rl_55_t1 = TR_67 ;
	7'h2d :
		RG_rl_55_t1 = TR_67 ;
	7'h2e :
		RG_rl_55_t1 = TR_67 ;
	7'h2f :
		RG_rl_55_t1 = TR_67 ;
	7'h30 :
		RG_rl_55_t1 = TR_67 ;
	7'h31 :
		RG_rl_55_t1 = TR_67 ;
	7'h32 :
		RG_rl_55_t1 = TR_67 ;
	7'h33 :
		RG_rl_55_t1 = TR_67 ;
	7'h34 :
		RG_rl_55_t1 = TR_67 ;
	7'h35 :
		RG_rl_55_t1 = TR_67 ;
	7'h36 :
		RG_rl_55_t1 = TR_67 ;
	7'h37 :
		RG_rl_55_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h38 :
		RG_rl_55_t1 = TR_67 ;
	7'h39 :
		RG_rl_55_t1 = TR_67 ;
	7'h3a :
		RG_rl_55_t1 = TR_67 ;
	7'h3b :
		RG_rl_55_t1 = TR_67 ;
	7'h3c :
		RG_rl_55_t1 = TR_67 ;
	7'h3d :
		RG_rl_55_t1 = TR_67 ;
	7'h3e :
		RG_rl_55_t1 = TR_67 ;
	7'h3f :
		RG_rl_55_t1 = TR_67 ;
	7'h40 :
		RG_rl_55_t1 = TR_67 ;
	7'h41 :
		RG_rl_55_t1 = TR_67 ;
	7'h42 :
		RG_rl_55_t1 = TR_67 ;
	7'h43 :
		RG_rl_55_t1 = TR_67 ;
	7'h44 :
		RG_rl_55_t1 = TR_67 ;
	7'h45 :
		RG_rl_55_t1 = TR_67 ;
	7'h46 :
		RG_rl_55_t1 = TR_67 ;
	7'h47 :
		RG_rl_55_t1 = TR_67 ;
	7'h48 :
		RG_rl_55_t1 = TR_67 ;
	7'h49 :
		RG_rl_55_t1 = TR_67 ;
	7'h4a :
		RG_rl_55_t1 = TR_67 ;
	7'h4b :
		RG_rl_55_t1 = TR_67 ;
	7'h4c :
		RG_rl_55_t1 = TR_67 ;
	7'h4d :
		RG_rl_55_t1 = TR_67 ;
	7'h4e :
		RG_rl_55_t1 = TR_67 ;
	7'h4f :
		RG_rl_55_t1 = TR_67 ;
	7'h50 :
		RG_rl_55_t1 = TR_67 ;
	7'h51 :
		RG_rl_55_t1 = TR_67 ;
	7'h52 :
		RG_rl_55_t1 = TR_67 ;
	7'h53 :
		RG_rl_55_t1 = TR_67 ;
	7'h54 :
		RG_rl_55_t1 = TR_67 ;
	7'h55 :
		RG_rl_55_t1 = TR_67 ;
	7'h56 :
		RG_rl_55_t1 = TR_67 ;
	7'h57 :
		RG_rl_55_t1 = TR_67 ;
	7'h58 :
		RG_rl_55_t1 = TR_67 ;
	7'h59 :
		RG_rl_55_t1 = TR_67 ;
	7'h5a :
		RG_rl_55_t1 = TR_67 ;
	7'h5b :
		RG_rl_55_t1 = TR_67 ;
	7'h5c :
		RG_rl_55_t1 = TR_67 ;
	7'h5d :
		RG_rl_55_t1 = TR_67 ;
	7'h5e :
		RG_rl_55_t1 = TR_67 ;
	7'h5f :
		RG_rl_55_t1 = TR_67 ;
	7'h60 :
		RG_rl_55_t1 = TR_67 ;
	7'h61 :
		RG_rl_55_t1 = TR_67 ;
	7'h62 :
		RG_rl_55_t1 = TR_67 ;
	7'h63 :
		RG_rl_55_t1 = TR_67 ;
	7'h64 :
		RG_rl_55_t1 = TR_67 ;
	7'h65 :
		RG_rl_55_t1 = TR_67 ;
	7'h66 :
		RG_rl_55_t1 = TR_67 ;
	7'h67 :
		RG_rl_55_t1 = TR_67 ;
	7'h68 :
		RG_rl_55_t1 = TR_67 ;
	7'h69 :
		RG_rl_55_t1 = TR_67 ;
	7'h6a :
		RG_rl_55_t1 = TR_67 ;
	7'h6b :
		RG_rl_55_t1 = TR_67 ;
	7'h6c :
		RG_rl_55_t1 = TR_67 ;
	7'h6d :
		RG_rl_55_t1 = TR_67 ;
	7'h6e :
		RG_rl_55_t1 = TR_67 ;
	7'h6f :
		RG_rl_55_t1 = TR_67 ;
	7'h70 :
		RG_rl_55_t1 = TR_67 ;
	7'h71 :
		RG_rl_55_t1 = TR_67 ;
	7'h72 :
		RG_rl_55_t1 = TR_67 ;
	7'h73 :
		RG_rl_55_t1 = TR_67 ;
	7'h74 :
		RG_rl_55_t1 = TR_67 ;
	7'h75 :
		RG_rl_55_t1 = TR_67 ;
	7'h76 :
		RG_rl_55_t1 = TR_67 ;
	7'h77 :
		RG_rl_55_t1 = TR_67 ;
	7'h78 :
		RG_rl_55_t1 = TR_67 ;
	7'h79 :
		RG_rl_55_t1 = TR_67 ;
	7'h7a :
		RG_rl_55_t1 = TR_67 ;
	7'h7b :
		RG_rl_55_t1 = TR_67 ;
	7'h7c :
		RG_rl_55_t1 = TR_67 ;
	7'h7d :
		RG_rl_55_t1 = TR_67 ;
	7'h7e :
		RG_rl_55_t1 = TR_67 ;
	7'h7f :
		RG_rl_55_t1 = TR_67 ;
	default :
		RG_rl_55_t1 = 9'hx ;
	endcase
always @ ( RG_rl_55_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_238 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_55_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h37 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_55_t = ( ( { 9{ U_570 } } & RG_rl_238 )
		| ( { 9{ U_569 } } & RG_rl_55_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_55_en = ( U_570 | RG_rl_55_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_55_en )
		RG_rl_55 <= RG_rl_55_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_68 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_56_t1 = TR_68 ;
	7'h01 :
		RG_rl_56_t1 = TR_68 ;
	7'h02 :
		RG_rl_56_t1 = TR_68 ;
	7'h03 :
		RG_rl_56_t1 = TR_68 ;
	7'h04 :
		RG_rl_56_t1 = TR_68 ;
	7'h05 :
		RG_rl_56_t1 = TR_68 ;
	7'h06 :
		RG_rl_56_t1 = TR_68 ;
	7'h07 :
		RG_rl_56_t1 = TR_68 ;
	7'h08 :
		RG_rl_56_t1 = TR_68 ;
	7'h09 :
		RG_rl_56_t1 = TR_68 ;
	7'h0a :
		RG_rl_56_t1 = TR_68 ;
	7'h0b :
		RG_rl_56_t1 = TR_68 ;
	7'h0c :
		RG_rl_56_t1 = TR_68 ;
	7'h0d :
		RG_rl_56_t1 = TR_68 ;
	7'h0e :
		RG_rl_56_t1 = TR_68 ;
	7'h0f :
		RG_rl_56_t1 = TR_68 ;
	7'h10 :
		RG_rl_56_t1 = TR_68 ;
	7'h11 :
		RG_rl_56_t1 = TR_68 ;
	7'h12 :
		RG_rl_56_t1 = TR_68 ;
	7'h13 :
		RG_rl_56_t1 = TR_68 ;
	7'h14 :
		RG_rl_56_t1 = TR_68 ;
	7'h15 :
		RG_rl_56_t1 = TR_68 ;
	7'h16 :
		RG_rl_56_t1 = TR_68 ;
	7'h17 :
		RG_rl_56_t1 = TR_68 ;
	7'h18 :
		RG_rl_56_t1 = TR_68 ;
	7'h19 :
		RG_rl_56_t1 = TR_68 ;
	7'h1a :
		RG_rl_56_t1 = TR_68 ;
	7'h1b :
		RG_rl_56_t1 = TR_68 ;
	7'h1c :
		RG_rl_56_t1 = TR_68 ;
	7'h1d :
		RG_rl_56_t1 = TR_68 ;
	7'h1e :
		RG_rl_56_t1 = TR_68 ;
	7'h1f :
		RG_rl_56_t1 = TR_68 ;
	7'h20 :
		RG_rl_56_t1 = TR_68 ;
	7'h21 :
		RG_rl_56_t1 = TR_68 ;
	7'h22 :
		RG_rl_56_t1 = TR_68 ;
	7'h23 :
		RG_rl_56_t1 = TR_68 ;
	7'h24 :
		RG_rl_56_t1 = TR_68 ;
	7'h25 :
		RG_rl_56_t1 = TR_68 ;
	7'h26 :
		RG_rl_56_t1 = TR_68 ;
	7'h27 :
		RG_rl_56_t1 = TR_68 ;
	7'h28 :
		RG_rl_56_t1 = TR_68 ;
	7'h29 :
		RG_rl_56_t1 = TR_68 ;
	7'h2a :
		RG_rl_56_t1 = TR_68 ;
	7'h2b :
		RG_rl_56_t1 = TR_68 ;
	7'h2c :
		RG_rl_56_t1 = TR_68 ;
	7'h2d :
		RG_rl_56_t1 = TR_68 ;
	7'h2e :
		RG_rl_56_t1 = TR_68 ;
	7'h2f :
		RG_rl_56_t1 = TR_68 ;
	7'h30 :
		RG_rl_56_t1 = TR_68 ;
	7'h31 :
		RG_rl_56_t1 = TR_68 ;
	7'h32 :
		RG_rl_56_t1 = TR_68 ;
	7'h33 :
		RG_rl_56_t1 = TR_68 ;
	7'h34 :
		RG_rl_56_t1 = TR_68 ;
	7'h35 :
		RG_rl_56_t1 = TR_68 ;
	7'h36 :
		RG_rl_56_t1 = TR_68 ;
	7'h37 :
		RG_rl_56_t1 = TR_68 ;
	7'h38 :
		RG_rl_56_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h39 :
		RG_rl_56_t1 = TR_68 ;
	7'h3a :
		RG_rl_56_t1 = TR_68 ;
	7'h3b :
		RG_rl_56_t1 = TR_68 ;
	7'h3c :
		RG_rl_56_t1 = TR_68 ;
	7'h3d :
		RG_rl_56_t1 = TR_68 ;
	7'h3e :
		RG_rl_56_t1 = TR_68 ;
	7'h3f :
		RG_rl_56_t1 = TR_68 ;
	7'h40 :
		RG_rl_56_t1 = TR_68 ;
	7'h41 :
		RG_rl_56_t1 = TR_68 ;
	7'h42 :
		RG_rl_56_t1 = TR_68 ;
	7'h43 :
		RG_rl_56_t1 = TR_68 ;
	7'h44 :
		RG_rl_56_t1 = TR_68 ;
	7'h45 :
		RG_rl_56_t1 = TR_68 ;
	7'h46 :
		RG_rl_56_t1 = TR_68 ;
	7'h47 :
		RG_rl_56_t1 = TR_68 ;
	7'h48 :
		RG_rl_56_t1 = TR_68 ;
	7'h49 :
		RG_rl_56_t1 = TR_68 ;
	7'h4a :
		RG_rl_56_t1 = TR_68 ;
	7'h4b :
		RG_rl_56_t1 = TR_68 ;
	7'h4c :
		RG_rl_56_t1 = TR_68 ;
	7'h4d :
		RG_rl_56_t1 = TR_68 ;
	7'h4e :
		RG_rl_56_t1 = TR_68 ;
	7'h4f :
		RG_rl_56_t1 = TR_68 ;
	7'h50 :
		RG_rl_56_t1 = TR_68 ;
	7'h51 :
		RG_rl_56_t1 = TR_68 ;
	7'h52 :
		RG_rl_56_t1 = TR_68 ;
	7'h53 :
		RG_rl_56_t1 = TR_68 ;
	7'h54 :
		RG_rl_56_t1 = TR_68 ;
	7'h55 :
		RG_rl_56_t1 = TR_68 ;
	7'h56 :
		RG_rl_56_t1 = TR_68 ;
	7'h57 :
		RG_rl_56_t1 = TR_68 ;
	7'h58 :
		RG_rl_56_t1 = TR_68 ;
	7'h59 :
		RG_rl_56_t1 = TR_68 ;
	7'h5a :
		RG_rl_56_t1 = TR_68 ;
	7'h5b :
		RG_rl_56_t1 = TR_68 ;
	7'h5c :
		RG_rl_56_t1 = TR_68 ;
	7'h5d :
		RG_rl_56_t1 = TR_68 ;
	7'h5e :
		RG_rl_56_t1 = TR_68 ;
	7'h5f :
		RG_rl_56_t1 = TR_68 ;
	7'h60 :
		RG_rl_56_t1 = TR_68 ;
	7'h61 :
		RG_rl_56_t1 = TR_68 ;
	7'h62 :
		RG_rl_56_t1 = TR_68 ;
	7'h63 :
		RG_rl_56_t1 = TR_68 ;
	7'h64 :
		RG_rl_56_t1 = TR_68 ;
	7'h65 :
		RG_rl_56_t1 = TR_68 ;
	7'h66 :
		RG_rl_56_t1 = TR_68 ;
	7'h67 :
		RG_rl_56_t1 = TR_68 ;
	7'h68 :
		RG_rl_56_t1 = TR_68 ;
	7'h69 :
		RG_rl_56_t1 = TR_68 ;
	7'h6a :
		RG_rl_56_t1 = TR_68 ;
	7'h6b :
		RG_rl_56_t1 = TR_68 ;
	7'h6c :
		RG_rl_56_t1 = TR_68 ;
	7'h6d :
		RG_rl_56_t1 = TR_68 ;
	7'h6e :
		RG_rl_56_t1 = TR_68 ;
	7'h6f :
		RG_rl_56_t1 = TR_68 ;
	7'h70 :
		RG_rl_56_t1 = TR_68 ;
	7'h71 :
		RG_rl_56_t1 = TR_68 ;
	7'h72 :
		RG_rl_56_t1 = TR_68 ;
	7'h73 :
		RG_rl_56_t1 = TR_68 ;
	7'h74 :
		RG_rl_56_t1 = TR_68 ;
	7'h75 :
		RG_rl_56_t1 = TR_68 ;
	7'h76 :
		RG_rl_56_t1 = TR_68 ;
	7'h77 :
		RG_rl_56_t1 = TR_68 ;
	7'h78 :
		RG_rl_56_t1 = TR_68 ;
	7'h79 :
		RG_rl_56_t1 = TR_68 ;
	7'h7a :
		RG_rl_56_t1 = TR_68 ;
	7'h7b :
		RG_rl_56_t1 = TR_68 ;
	7'h7c :
		RG_rl_56_t1 = TR_68 ;
	7'h7d :
		RG_rl_56_t1 = TR_68 ;
	7'h7e :
		RG_rl_56_t1 = TR_68 ;
	7'h7f :
		RG_rl_56_t1 = TR_68 ;
	default :
		RG_rl_56_t1 = 9'hx ;
	endcase
always @ ( RG_rl_56_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_239 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_56_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h38 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_56_t = ( ( { 9{ U_570 } } & RG_rl_239 )
		| ( { 9{ U_569 } } & RG_rl_56_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_56_en = ( U_570 | RG_rl_56_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_56_en )
		RG_rl_56 <= RG_rl_56_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_69 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_57_t1 = TR_69 ;
	7'h01 :
		RG_rl_57_t1 = TR_69 ;
	7'h02 :
		RG_rl_57_t1 = TR_69 ;
	7'h03 :
		RG_rl_57_t1 = TR_69 ;
	7'h04 :
		RG_rl_57_t1 = TR_69 ;
	7'h05 :
		RG_rl_57_t1 = TR_69 ;
	7'h06 :
		RG_rl_57_t1 = TR_69 ;
	7'h07 :
		RG_rl_57_t1 = TR_69 ;
	7'h08 :
		RG_rl_57_t1 = TR_69 ;
	7'h09 :
		RG_rl_57_t1 = TR_69 ;
	7'h0a :
		RG_rl_57_t1 = TR_69 ;
	7'h0b :
		RG_rl_57_t1 = TR_69 ;
	7'h0c :
		RG_rl_57_t1 = TR_69 ;
	7'h0d :
		RG_rl_57_t1 = TR_69 ;
	7'h0e :
		RG_rl_57_t1 = TR_69 ;
	7'h0f :
		RG_rl_57_t1 = TR_69 ;
	7'h10 :
		RG_rl_57_t1 = TR_69 ;
	7'h11 :
		RG_rl_57_t1 = TR_69 ;
	7'h12 :
		RG_rl_57_t1 = TR_69 ;
	7'h13 :
		RG_rl_57_t1 = TR_69 ;
	7'h14 :
		RG_rl_57_t1 = TR_69 ;
	7'h15 :
		RG_rl_57_t1 = TR_69 ;
	7'h16 :
		RG_rl_57_t1 = TR_69 ;
	7'h17 :
		RG_rl_57_t1 = TR_69 ;
	7'h18 :
		RG_rl_57_t1 = TR_69 ;
	7'h19 :
		RG_rl_57_t1 = TR_69 ;
	7'h1a :
		RG_rl_57_t1 = TR_69 ;
	7'h1b :
		RG_rl_57_t1 = TR_69 ;
	7'h1c :
		RG_rl_57_t1 = TR_69 ;
	7'h1d :
		RG_rl_57_t1 = TR_69 ;
	7'h1e :
		RG_rl_57_t1 = TR_69 ;
	7'h1f :
		RG_rl_57_t1 = TR_69 ;
	7'h20 :
		RG_rl_57_t1 = TR_69 ;
	7'h21 :
		RG_rl_57_t1 = TR_69 ;
	7'h22 :
		RG_rl_57_t1 = TR_69 ;
	7'h23 :
		RG_rl_57_t1 = TR_69 ;
	7'h24 :
		RG_rl_57_t1 = TR_69 ;
	7'h25 :
		RG_rl_57_t1 = TR_69 ;
	7'h26 :
		RG_rl_57_t1 = TR_69 ;
	7'h27 :
		RG_rl_57_t1 = TR_69 ;
	7'h28 :
		RG_rl_57_t1 = TR_69 ;
	7'h29 :
		RG_rl_57_t1 = TR_69 ;
	7'h2a :
		RG_rl_57_t1 = TR_69 ;
	7'h2b :
		RG_rl_57_t1 = TR_69 ;
	7'h2c :
		RG_rl_57_t1 = TR_69 ;
	7'h2d :
		RG_rl_57_t1 = TR_69 ;
	7'h2e :
		RG_rl_57_t1 = TR_69 ;
	7'h2f :
		RG_rl_57_t1 = TR_69 ;
	7'h30 :
		RG_rl_57_t1 = TR_69 ;
	7'h31 :
		RG_rl_57_t1 = TR_69 ;
	7'h32 :
		RG_rl_57_t1 = TR_69 ;
	7'h33 :
		RG_rl_57_t1 = TR_69 ;
	7'h34 :
		RG_rl_57_t1 = TR_69 ;
	7'h35 :
		RG_rl_57_t1 = TR_69 ;
	7'h36 :
		RG_rl_57_t1 = TR_69 ;
	7'h37 :
		RG_rl_57_t1 = TR_69 ;
	7'h38 :
		RG_rl_57_t1 = TR_69 ;
	7'h39 :
		RG_rl_57_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3a :
		RG_rl_57_t1 = TR_69 ;
	7'h3b :
		RG_rl_57_t1 = TR_69 ;
	7'h3c :
		RG_rl_57_t1 = TR_69 ;
	7'h3d :
		RG_rl_57_t1 = TR_69 ;
	7'h3e :
		RG_rl_57_t1 = TR_69 ;
	7'h3f :
		RG_rl_57_t1 = TR_69 ;
	7'h40 :
		RG_rl_57_t1 = TR_69 ;
	7'h41 :
		RG_rl_57_t1 = TR_69 ;
	7'h42 :
		RG_rl_57_t1 = TR_69 ;
	7'h43 :
		RG_rl_57_t1 = TR_69 ;
	7'h44 :
		RG_rl_57_t1 = TR_69 ;
	7'h45 :
		RG_rl_57_t1 = TR_69 ;
	7'h46 :
		RG_rl_57_t1 = TR_69 ;
	7'h47 :
		RG_rl_57_t1 = TR_69 ;
	7'h48 :
		RG_rl_57_t1 = TR_69 ;
	7'h49 :
		RG_rl_57_t1 = TR_69 ;
	7'h4a :
		RG_rl_57_t1 = TR_69 ;
	7'h4b :
		RG_rl_57_t1 = TR_69 ;
	7'h4c :
		RG_rl_57_t1 = TR_69 ;
	7'h4d :
		RG_rl_57_t1 = TR_69 ;
	7'h4e :
		RG_rl_57_t1 = TR_69 ;
	7'h4f :
		RG_rl_57_t1 = TR_69 ;
	7'h50 :
		RG_rl_57_t1 = TR_69 ;
	7'h51 :
		RG_rl_57_t1 = TR_69 ;
	7'h52 :
		RG_rl_57_t1 = TR_69 ;
	7'h53 :
		RG_rl_57_t1 = TR_69 ;
	7'h54 :
		RG_rl_57_t1 = TR_69 ;
	7'h55 :
		RG_rl_57_t1 = TR_69 ;
	7'h56 :
		RG_rl_57_t1 = TR_69 ;
	7'h57 :
		RG_rl_57_t1 = TR_69 ;
	7'h58 :
		RG_rl_57_t1 = TR_69 ;
	7'h59 :
		RG_rl_57_t1 = TR_69 ;
	7'h5a :
		RG_rl_57_t1 = TR_69 ;
	7'h5b :
		RG_rl_57_t1 = TR_69 ;
	7'h5c :
		RG_rl_57_t1 = TR_69 ;
	7'h5d :
		RG_rl_57_t1 = TR_69 ;
	7'h5e :
		RG_rl_57_t1 = TR_69 ;
	7'h5f :
		RG_rl_57_t1 = TR_69 ;
	7'h60 :
		RG_rl_57_t1 = TR_69 ;
	7'h61 :
		RG_rl_57_t1 = TR_69 ;
	7'h62 :
		RG_rl_57_t1 = TR_69 ;
	7'h63 :
		RG_rl_57_t1 = TR_69 ;
	7'h64 :
		RG_rl_57_t1 = TR_69 ;
	7'h65 :
		RG_rl_57_t1 = TR_69 ;
	7'h66 :
		RG_rl_57_t1 = TR_69 ;
	7'h67 :
		RG_rl_57_t1 = TR_69 ;
	7'h68 :
		RG_rl_57_t1 = TR_69 ;
	7'h69 :
		RG_rl_57_t1 = TR_69 ;
	7'h6a :
		RG_rl_57_t1 = TR_69 ;
	7'h6b :
		RG_rl_57_t1 = TR_69 ;
	7'h6c :
		RG_rl_57_t1 = TR_69 ;
	7'h6d :
		RG_rl_57_t1 = TR_69 ;
	7'h6e :
		RG_rl_57_t1 = TR_69 ;
	7'h6f :
		RG_rl_57_t1 = TR_69 ;
	7'h70 :
		RG_rl_57_t1 = TR_69 ;
	7'h71 :
		RG_rl_57_t1 = TR_69 ;
	7'h72 :
		RG_rl_57_t1 = TR_69 ;
	7'h73 :
		RG_rl_57_t1 = TR_69 ;
	7'h74 :
		RG_rl_57_t1 = TR_69 ;
	7'h75 :
		RG_rl_57_t1 = TR_69 ;
	7'h76 :
		RG_rl_57_t1 = TR_69 ;
	7'h77 :
		RG_rl_57_t1 = TR_69 ;
	7'h78 :
		RG_rl_57_t1 = TR_69 ;
	7'h79 :
		RG_rl_57_t1 = TR_69 ;
	7'h7a :
		RG_rl_57_t1 = TR_69 ;
	7'h7b :
		RG_rl_57_t1 = TR_69 ;
	7'h7c :
		RG_rl_57_t1 = TR_69 ;
	7'h7d :
		RG_rl_57_t1 = TR_69 ;
	7'h7e :
		RG_rl_57_t1 = TR_69 ;
	7'h7f :
		RG_rl_57_t1 = TR_69 ;
	default :
		RG_rl_57_t1 = 9'hx ;
	endcase
always @ ( RG_rl_57_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_240 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_57_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h39 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_57_t = ( ( { 9{ U_570 } } & RG_rl_240 )
		| ( { 9{ U_569 } } & RG_rl_57_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_57_en = ( U_570 | RG_rl_57_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_57_en )
		RG_rl_57 <= RG_rl_57_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_70 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_58_t1 = TR_70 ;
	7'h01 :
		RG_rl_58_t1 = TR_70 ;
	7'h02 :
		RG_rl_58_t1 = TR_70 ;
	7'h03 :
		RG_rl_58_t1 = TR_70 ;
	7'h04 :
		RG_rl_58_t1 = TR_70 ;
	7'h05 :
		RG_rl_58_t1 = TR_70 ;
	7'h06 :
		RG_rl_58_t1 = TR_70 ;
	7'h07 :
		RG_rl_58_t1 = TR_70 ;
	7'h08 :
		RG_rl_58_t1 = TR_70 ;
	7'h09 :
		RG_rl_58_t1 = TR_70 ;
	7'h0a :
		RG_rl_58_t1 = TR_70 ;
	7'h0b :
		RG_rl_58_t1 = TR_70 ;
	7'h0c :
		RG_rl_58_t1 = TR_70 ;
	7'h0d :
		RG_rl_58_t1 = TR_70 ;
	7'h0e :
		RG_rl_58_t1 = TR_70 ;
	7'h0f :
		RG_rl_58_t1 = TR_70 ;
	7'h10 :
		RG_rl_58_t1 = TR_70 ;
	7'h11 :
		RG_rl_58_t1 = TR_70 ;
	7'h12 :
		RG_rl_58_t1 = TR_70 ;
	7'h13 :
		RG_rl_58_t1 = TR_70 ;
	7'h14 :
		RG_rl_58_t1 = TR_70 ;
	7'h15 :
		RG_rl_58_t1 = TR_70 ;
	7'h16 :
		RG_rl_58_t1 = TR_70 ;
	7'h17 :
		RG_rl_58_t1 = TR_70 ;
	7'h18 :
		RG_rl_58_t1 = TR_70 ;
	7'h19 :
		RG_rl_58_t1 = TR_70 ;
	7'h1a :
		RG_rl_58_t1 = TR_70 ;
	7'h1b :
		RG_rl_58_t1 = TR_70 ;
	7'h1c :
		RG_rl_58_t1 = TR_70 ;
	7'h1d :
		RG_rl_58_t1 = TR_70 ;
	7'h1e :
		RG_rl_58_t1 = TR_70 ;
	7'h1f :
		RG_rl_58_t1 = TR_70 ;
	7'h20 :
		RG_rl_58_t1 = TR_70 ;
	7'h21 :
		RG_rl_58_t1 = TR_70 ;
	7'h22 :
		RG_rl_58_t1 = TR_70 ;
	7'h23 :
		RG_rl_58_t1 = TR_70 ;
	7'h24 :
		RG_rl_58_t1 = TR_70 ;
	7'h25 :
		RG_rl_58_t1 = TR_70 ;
	7'h26 :
		RG_rl_58_t1 = TR_70 ;
	7'h27 :
		RG_rl_58_t1 = TR_70 ;
	7'h28 :
		RG_rl_58_t1 = TR_70 ;
	7'h29 :
		RG_rl_58_t1 = TR_70 ;
	7'h2a :
		RG_rl_58_t1 = TR_70 ;
	7'h2b :
		RG_rl_58_t1 = TR_70 ;
	7'h2c :
		RG_rl_58_t1 = TR_70 ;
	7'h2d :
		RG_rl_58_t1 = TR_70 ;
	7'h2e :
		RG_rl_58_t1 = TR_70 ;
	7'h2f :
		RG_rl_58_t1 = TR_70 ;
	7'h30 :
		RG_rl_58_t1 = TR_70 ;
	7'h31 :
		RG_rl_58_t1 = TR_70 ;
	7'h32 :
		RG_rl_58_t1 = TR_70 ;
	7'h33 :
		RG_rl_58_t1 = TR_70 ;
	7'h34 :
		RG_rl_58_t1 = TR_70 ;
	7'h35 :
		RG_rl_58_t1 = TR_70 ;
	7'h36 :
		RG_rl_58_t1 = TR_70 ;
	7'h37 :
		RG_rl_58_t1 = TR_70 ;
	7'h38 :
		RG_rl_58_t1 = TR_70 ;
	7'h39 :
		RG_rl_58_t1 = TR_70 ;
	7'h3a :
		RG_rl_58_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3b :
		RG_rl_58_t1 = TR_70 ;
	7'h3c :
		RG_rl_58_t1 = TR_70 ;
	7'h3d :
		RG_rl_58_t1 = TR_70 ;
	7'h3e :
		RG_rl_58_t1 = TR_70 ;
	7'h3f :
		RG_rl_58_t1 = TR_70 ;
	7'h40 :
		RG_rl_58_t1 = TR_70 ;
	7'h41 :
		RG_rl_58_t1 = TR_70 ;
	7'h42 :
		RG_rl_58_t1 = TR_70 ;
	7'h43 :
		RG_rl_58_t1 = TR_70 ;
	7'h44 :
		RG_rl_58_t1 = TR_70 ;
	7'h45 :
		RG_rl_58_t1 = TR_70 ;
	7'h46 :
		RG_rl_58_t1 = TR_70 ;
	7'h47 :
		RG_rl_58_t1 = TR_70 ;
	7'h48 :
		RG_rl_58_t1 = TR_70 ;
	7'h49 :
		RG_rl_58_t1 = TR_70 ;
	7'h4a :
		RG_rl_58_t1 = TR_70 ;
	7'h4b :
		RG_rl_58_t1 = TR_70 ;
	7'h4c :
		RG_rl_58_t1 = TR_70 ;
	7'h4d :
		RG_rl_58_t1 = TR_70 ;
	7'h4e :
		RG_rl_58_t1 = TR_70 ;
	7'h4f :
		RG_rl_58_t1 = TR_70 ;
	7'h50 :
		RG_rl_58_t1 = TR_70 ;
	7'h51 :
		RG_rl_58_t1 = TR_70 ;
	7'h52 :
		RG_rl_58_t1 = TR_70 ;
	7'h53 :
		RG_rl_58_t1 = TR_70 ;
	7'h54 :
		RG_rl_58_t1 = TR_70 ;
	7'h55 :
		RG_rl_58_t1 = TR_70 ;
	7'h56 :
		RG_rl_58_t1 = TR_70 ;
	7'h57 :
		RG_rl_58_t1 = TR_70 ;
	7'h58 :
		RG_rl_58_t1 = TR_70 ;
	7'h59 :
		RG_rl_58_t1 = TR_70 ;
	7'h5a :
		RG_rl_58_t1 = TR_70 ;
	7'h5b :
		RG_rl_58_t1 = TR_70 ;
	7'h5c :
		RG_rl_58_t1 = TR_70 ;
	7'h5d :
		RG_rl_58_t1 = TR_70 ;
	7'h5e :
		RG_rl_58_t1 = TR_70 ;
	7'h5f :
		RG_rl_58_t1 = TR_70 ;
	7'h60 :
		RG_rl_58_t1 = TR_70 ;
	7'h61 :
		RG_rl_58_t1 = TR_70 ;
	7'h62 :
		RG_rl_58_t1 = TR_70 ;
	7'h63 :
		RG_rl_58_t1 = TR_70 ;
	7'h64 :
		RG_rl_58_t1 = TR_70 ;
	7'h65 :
		RG_rl_58_t1 = TR_70 ;
	7'h66 :
		RG_rl_58_t1 = TR_70 ;
	7'h67 :
		RG_rl_58_t1 = TR_70 ;
	7'h68 :
		RG_rl_58_t1 = TR_70 ;
	7'h69 :
		RG_rl_58_t1 = TR_70 ;
	7'h6a :
		RG_rl_58_t1 = TR_70 ;
	7'h6b :
		RG_rl_58_t1 = TR_70 ;
	7'h6c :
		RG_rl_58_t1 = TR_70 ;
	7'h6d :
		RG_rl_58_t1 = TR_70 ;
	7'h6e :
		RG_rl_58_t1 = TR_70 ;
	7'h6f :
		RG_rl_58_t1 = TR_70 ;
	7'h70 :
		RG_rl_58_t1 = TR_70 ;
	7'h71 :
		RG_rl_58_t1 = TR_70 ;
	7'h72 :
		RG_rl_58_t1 = TR_70 ;
	7'h73 :
		RG_rl_58_t1 = TR_70 ;
	7'h74 :
		RG_rl_58_t1 = TR_70 ;
	7'h75 :
		RG_rl_58_t1 = TR_70 ;
	7'h76 :
		RG_rl_58_t1 = TR_70 ;
	7'h77 :
		RG_rl_58_t1 = TR_70 ;
	7'h78 :
		RG_rl_58_t1 = TR_70 ;
	7'h79 :
		RG_rl_58_t1 = TR_70 ;
	7'h7a :
		RG_rl_58_t1 = TR_70 ;
	7'h7b :
		RG_rl_58_t1 = TR_70 ;
	7'h7c :
		RG_rl_58_t1 = TR_70 ;
	7'h7d :
		RG_rl_58_t1 = TR_70 ;
	7'h7e :
		RG_rl_58_t1 = TR_70 ;
	7'h7f :
		RG_rl_58_t1 = TR_70 ;
	default :
		RG_rl_58_t1 = 9'hx ;
	endcase
always @ ( RG_rl_58_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_241 or U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_58_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h3a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_58_t = ( ( { 9{ U_570 } } & RG_rl_241 )
		| ( { 9{ U_569 } } & RG_rl_58_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_58_en = ( U_570 | RG_rl_58_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_58_en )
		RG_rl_58 <= RG_rl_58_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_71 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_59_t1 = TR_71 ;
	7'h01 :
		RG_rl_59_t1 = TR_71 ;
	7'h02 :
		RG_rl_59_t1 = TR_71 ;
	7'h03 :
		RG_rl_59_t1 = TR_71 ;
	7'h04 :
		RG_rl_59_t1 = TR_71 ;
	7'h05 :
		RG_rl_59_t1 = TR_71 ;
	7'h06 :
		RG_rl_59_t1 = TR_71 ;
	7'h07 :
		RG_rl_59_t1 = TR_71 ;
	7'h08 :
		RG_rl_59_t1 = TR_71 ;
	7'h09 :
		RG_rl_59_t1 = TR_71 ;
	7'h0a :
		RG_rl_59_t1 = TR_71 ;
	7'h0b :
		RG_rl_59_t1 = TR_71 ;
	7'h0c :
		RG_rl_59_t1 = TR_71 ;
	7'h0d :
		RG_rl_59_t1 = TR_71 ;
	7'h0e :
		RG_rl_59_t1 = TR_71 ;
	7'h0f :
		RG_rl_59_t1 = TR_71 ;
	7'h10 :
		RG_rl_59_t1 = TR_71 ;
	7'h11 :
		RG_rl_59_t1 = TR_71 ;
	7'h12 :
		RG_rl_59_t1 = TR_71 ;
	7'h13 :
		RG_rl_59_t1 = TR_71 ;
	7'h14 :
		RG_rl_59_t1 = TR_71 ;
	7'h15 :
		RG_rl_59_t1 = TR_71 ;
	7'h16 :
		RG_rl_59_t1 = TR_71 ;
	7'h17 :
		RG_rl_59_t1 = TR_71 ;
	7'h18 :
		RG_rl_59_t1 = TR_71 ;
	7'h19 :
		RG_rl_59_t1 = TR_71 ;
	7'h1a :
		RG_rl_59_t1 = TR_71 ;
	7'h1b :
		RG_rl_59_t1 = TR_71 ;
	7'h1c :
		RG_rl_59_t1 = TR_71 ;
	7'h1d :
		RG_rl_59_t1 = TR_71 ;
	7'h1e :
		RG_rl_59_t1 = TR_71 ;
	7'h1f :
		RG_rl_59_t1 = TR_71 ;
	7'h20 :
		RG_rl_59_t1 = TR_71 ;
	7'h21 :
		RG_rl_59_t1 = TR_71 ;
	7'h22 :
		RG_rl_59_t1 = TR_71 ;
	7'h23 :
		RG_rl_59_t1 = TR_71 ;
	7'h24 :
		RG_rl_59_t1 = TR_71 ;
	7'h25 :
		RG_rl_59_t1 = TR_71 ;
	7'h26 :
		RG_rl_59_t1 = TR_71 ;
	7'h27 :
		RG_rl_59_t1 = TR_71 ;
	7'h28 :
		RG_rl_59_t1 = TR_71 ;
	7'h29 :
		RG_rl_59_t1 = TR_71 ;
	7'h2a :
		RG_rl_59_t1 = TR_71 ;
	7'h2b :
		RG_rl_59_t1 = TR_71 ;
	7'h2c :
		RG_rl_59_t1 = TR_71 ;
	7'h2d :
		RG_rl_59_t1 = TR_71 ;
	7'h2e :
		RG_rl_59_t1 = TR_71 ;
	7'h2f :
		RG_rl_59_t1 = TR_71 ;
	7'h30 :
		RG_rl_59_t1 = TR_71 ;
	7'h31 :
		RG_rl_59_t1 = TR_71 ;
	7'h32 :
		RG_rl_59_t1 = TR_71 ;
	7'h33 :
		RG_rl_59_t1 = TR_71 ;
	7'h34 :
		RG_rl_59_t1 = TR_71 ;
	7'h35 :
		RG_rl_59_t1 = TR_71 ;
	7'h36 :
		RG_rl_59_t1 = TR_71 ;
	7'h37 :
		RG_rl_59_t1 = TR_71 ;
	7'h38 :
		RG_rl_59_t1 = TR_71 ;
	7'h39 :
		RG_rl_59_t1 = TR_71 ;
	7'h3a :
		RG_rl_59_t1 = TR_71 ;
	7'h3b :
		RG_rl_59_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3c :
		RG_rl_59_t1 = TR_71 ;
	7'h3d :
		RG_rl_59_t1 = TR_71 ;
	7'h3e :
		RG_rl_59_t1 = TR_71 ;
	7'h3f :
		RG_rl_59_t1 = TR_71 ;
	7'h40 :
		RG_rl_59_t1 = TR_71 ;
	7'h41 :
		RG_rl_59_t1 = TR_71 ;
	7'h42 :
		RG_rl_59_t1 = TR_71 ;
	7'h43 :
		RG_rl_59_t1 = TR_71 ;
	7'h44 :
		RG_rl_59_t1 = TR_71 ;
	7'h45 :
		RG_rl_59_t1 = TR_71 ;
	7'h46 :
		RG_rl_59_t1 = TR_71 ;
	7'h47 :
		RG_rl_59_t1 = TR_71 ;
	7'h48 :
		RG_rl_59_t1 = TR_71 ;
	7'h49 :
		RG_rl_59_t1 = TR_71 ;
	7'h4a :
		RG_rl_59_t1 = TR_71 ;
	7'h4b :
		RG_rl_59_t1 = TR_71 ;
	7'h4c :
		RG_rl_59_t1 = TR_71 ;
	7'h4d :
		RG_rl_59_t1 = TR_71 ;
	7'h4e :
		RG_rl_59_t1 = TR_71 ;
	7'h4f :
		RG_rl_59_t1 = TR_71 ;
	7'h50 :
		RG_rl_59_t1 = TR_71 ;
	7'h51 :
		RG_rl_59_t1 = TR_71 ;
	7'h52 :
		RG_rl_59_t1 = TR_71 ;
	7'h53 :
		RG_rl_59_t1 = TR_71 ;
	7'h54 :
		RG_rl_59_t1 = TR_71 ;
	7'h55 :
		RG_rl_59_t1 = TR_71 ;
	7'h56 :
		RG_rl_59_t1 = TR_71 ;
	7'h57 :
		RG_rl_59_t1 = TR_71 ;
	7'h58 :
		RG_rl_59_t1 = TR_71 ;
	7'h59 :
		RG_rl_59_t1 = TR_71 ;
	7'h5a :
		RG_rl_59_t1 = TR_71 ;
	7'h5b :
		RG_rl_59_t1 = TR_71 ;
	7'h5c :
		RG_rl_59_t1 = TR_71 ;
	7'h5d :
		RG_rl_59_t1 = TR_71 ;
	7'h5e :
		RG_rl_59_t1 = TR_71 ;
	7'h5f :
		RG_rl_59_t1 = TR_71 ;
	7'h60 :
		RG_rl_59_t1 = TR_71 ;
	7'h61 :
		RG_rl_59_t1 = TR_71 ;
	7'h62 :
		RG_rl_59_t1 = TR_71 ;
	7'h63 :
		RG_rl_59_t1 = TR_71 ;
	7'h64 :
		RG_rl_59_t1 = TR_71 ;
	7'h65 :
		RG_rl_59_t1 = TR_71 ;
	7'h66 :
		RG_rl_59_t1 = TR_71 ;
	7'h67 :
		RG_rl_59_t1 = TR_71 ;
	7'h68 :
		RG_rl_59_t1 = TR_71 ;
	7'h69 :
		RG_rl_59_t1 = TR_71 ;
	7'h6a :
		RG_rl_59_t1 = TR_71 ;
	7'h6b :
		RG_rl_59_t1 = TR_71 ;
	7'h6c :
		RG_rl_59_t1 = TR_71 ;
	7'h6d :
		RG_rl_59_t1 = TR_71 ;
	7'h6e :
		RG_rl_59_t1 = TR_71 ;
	7'h6f :
		RG_rl_59_t1 = TR_71 ;
	7'h70 :
		RG_rl_59_t1 = TR_71 ;
	7'h71 :
		RG_rl_59_t1 = TR_71 ;
	7'h72 :
		RG_rl_59_t1 = TR_71 ;
	7'h73 :
		RG_rl_59_t1 = TR_71 ;
	7'h74 :
		RG_rl_59_t1 = TR_71 ;
	7'h75 :
		RG_rl_59_t1 = TR_71 ;
	7'h76 :
		RG_rl_59_t1 = TR_71 ;
	7'h77 :
		RG_rl_59_t1 = TR_71 ;
	7'h78 :
		RG_rl_59_t1 = TR_71 ;
	7'h79 :
		RG_rl_59_t1 = TR_71 ;
	7'h7a :
		RG_rl_59_t1 = TR_71 ;
	7'h7b :
		RG_rl_59_t1 = TR_71 ;
	7'h7c :
		RG_rl_59_t1 = TR_71 ;
	7'h7d :
		RG_rl_59_t1 = TR_71 ;
	7'h7e :
		RG_rl_59_t1 = TR_71 ;
	7'h7f :
		RG_rl_59_t1 = TR_71 ;
	default :
		RG_rl_59_t1 = 9'hx ;
	endcase
always @ ( RG_rl_59_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_59_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h3b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_59_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl )
		| ( { 9{ U_569 } } & RG_rl_59_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_59_en = ( U_570 | RG_rl_59_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_59_en )
		RG_rl_59 <= RG_rl_59_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_72 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_60_t1 = TR_72 ;
	7'h01 :
		RG_rl_60_t1 = TR_72 ;
	7'h02 :
		RG_rl_60_t1 = TR_72 ;
	7'h03 :
		RG_rl_60_t1 = TR_72 ;
	7'h04 :
		RG_rl_60_t1 = TR_72 ;
	7'h05 :
		RG_rl_60_t1 = TR_72 ;
	7'h06 :
		RG_rl_60_t1 = TR_72 ;
	7'h07 :
		RG_rl_60_t1 = TR_72 ;
	7'h08 :
		RG_rl_60_t1 = TR_72 ;
	7'h09 :
		RG_rl_60_t1 = TR_72 ;
	7'h0a :
		RG_rl_60_t1 = TR_72 ;
	7'h0b :
		RG_rl_60_t1 = TR_72 ;
	7'h0c :
		RG_rl_60_t1 = TR_72 ;
	7'h0d :
		RG_rl_60_t1 = TR_72 ;
	7'h0e :
		RG_rl_60_t1 = TR_72 ;
	7'h0f :
		RG_rl_60_t1 = TR_72 ;
	7'h10 :
		RG_rl_60_t1 = TR_72 ;
	7'h11 :
		RG_rl_60_t1 = TR_72 ;
	7'h12 :
		RG_rl_60_t1 = TR_72 ;
	7'h13 :
		RG_rl_60_t1 = TR_72 ;
	7'h14 :
		RG_rl_60_t1 = TR_72 ;
	7'h15 :
		RG_rl_60_t1 = TR_72 ;
	7'h16 :
		RG_rl_60_t1 = TR_72 ;
	7'h17 :
		RG_rl_60_t1 = TR_72 ;
	7'h18 :
		RG_rl_60_t1 = TR_72 ;
	7'h19 :
		RG_rl_60_t1 = TR_72 ;
	7'h1a :
		RG_rl_60_t1 = TR_72 ;
	7'h1b :
		RG_rl_60_t1 = TR_72 ;
	7'h1c :
		RG_rl_60_t1 = TR_72 ;
	7'h1d :
		RG_rl_60_t1 = TR_72 ;
	7'h1e :
		RG_rl_60_t1 = TR_72 ;
	7'h1f :
		RG_rl_60_t1 = TR_72 ;
	7'h20 :
		RG_rl_60_t1 = TR_72 ;
	7'h21 :
		RG_rl_60_t1 = TR_72 ;
	7'h22 :
		RG_rl_60_t1 = TR_72 ;
	7'h23 :
		RG_rl_60_t1 = TR_72 ;
	7'h24 :
		RG_rl_60_t1 = TR_72 ;
	7'h25 :
		RG_rl_60_t1 = TR_72 ;
	7'h26 :
		RG_rl_60_t1 = TR_72 ;
	7'h27 :
		RG_rl_60_t1 = TR_72 ;
	7'h28 :
		RG_rl_60_t1 = TR_72 ;
	7'h29 :
		RG_rl_60_t1 = TR_72 ;
	7'h2a :
		RG_rl_60_t1 = TR_72 ;
	7'h2b :
		RG_rl_60_t1 = TR_72 ;
	7'h2c :
		RG_rl_60_t1 = TR_72 ;
	7'h2d :
		RG_rl_60_t1 = TR_72 ;
	7'h2e :
		RG_rl_60_t1 = TR_72 ;
	7'h2f :
		RG_rl_60_t1 = TR_72 ;
	7'h30 :
		RG_rl_60_t1 = TR_72 ;
	7'h31 :
		RG_rl_60_t1 = TR_72 ;
	7'h32 :
		RG_rl_60_t1 = TR_72 ;
	7'h33 :
		RG_rl_60_t1 = TR_72 ;
	7'h34 :
		RG_rl_60_t1 = TR_72 ;
	7'h35 :
		RG_rl_60_t1 = TR_72 ;
	7'h36 :
		RG_rl_60_t1 = TR_72 ;
	7'h37 :
		RG_rl_60_t1 = TR_72 ;
	7'h38 :
		RG_rl_60_t1 = TR_72 ;
	7'h39 :
		RG_rl_60_t1 = TR_72 ;
	7'h3a :
		RG_rl_60_t1 = TR_72 ;
	7'h3b :
		RG_rl_60_t1 = TR_72 ;
	7'h3c :
		RG_rl_60_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3d :
		RG_rl_60_t1 = TR_72 ;
	7'h3e :
		RG_rl_60_t1 = TR_72 ;
	7'h3f :
		RG_rl_60_t1 = TR_72 ;
	7'h40 :
		RG_rl_60_t1 = TR_72 ;
	7'h41 :
		RG_rl_60_t1 = TR_72 ;
	7'h42 :
		RG_rl_60_t1 = TR_72 ;
	7'h43 :
		RG_rl_60_t1 = TR_72 ;
	7'h44 :
		RG_rl_60_t1 = TR_72 ;
	7'h45 :
		RG_rl_60_t1 = TR_72 ;
	7'h46 :
		RG_rl_60_t1 = TR_72 ;
	7'h47 :
		RG_rl_60_t1 = TR_72 ;
	7'h48 :
		RG_rl_60_t1 = TR_72 ;
	7'h49 :
		RG_rl_60_t1 = TR_72 ;
	7'h4a :
		RG_rl_60_t1 = TR_72 ;
	7'h4b :
		RG_rl_60_t1 = TR_72 ;
	7'h4c :
		RG_rl_60_t1 = TR_72 ;
	7'h4d :
		RG_rl_60_t1 = TR_72 ;
	7'h4e :
		RG_rl_60_t1 = TR_72 ;
	7'h4f :
		RG_rl_60_t1 = TR_72 ;
	7'h50 :
		RG_rl_60_t1 = TR_72 ;
	7'h51 :
		RG_rl_60_t1 = TR_72 ;
	7'h52 :
		RG_rl_60_t1 = TR_72 ;
	7'h53 :
		RG_rl_60_t1 = TR_72 ;
	7'h54 :
		RG_rl_60_t1 = TR_72 ;
	7'h55 :
		RG_rl_60_t1 = TR_72 ;
	7'h56 :
		RG_rl_60_t1 = TR_72 ;
	7'h57 :
		RG_rl_60_t1 = TR_72 ;
	7'h58 :
		RG_rl_60_t1 = TR_72 ;
	7'h59 :
		RG_rl_60_t1 = TR_72 ;
	7'h5a :
		RG_rl_60_t1 = TR_72 ;
	7'h5b :
		RG_rl_60_t1 = TR_72 ;
	7'h5c :
		RG_rl_60_t1 = TR_72 ;
	7'h5d :
		RG_rl_60_t1 = TR_72 ;
	7'h5e :
		RG_rl_60_t1 = TR_72 ;
	7'h5f :
		RG_rl_60_t1 = TR_72 ;
	7'h60 :
		RG_rl_60_t1 = TR_72 ;
	7'h61 :
		RG_rl_60_t1 = TR_72 ;
	7'h62 :
		RG_rl_60_t1 = TR_72 ;
	7'h63 :
		RG_rl_60_t1 = TR_72 ;
	7'h64 :
		RG_rl_60_t1 = TR_72 ;
	7'h65 :
		RG_rl_60_t1 = TR_72 ;
	7'h66 :
		RG_rl_60_t1 = TR_72 ;
	7'h67 :
		RG_rl_60_t1 = TR_72 ;
	7'h68 :
		RG_rl_60_t1 = TR_72 ;
	7'h69 :
		RG_rl_60_t1 = TR_72 ;
	7'h6a :
		RG_rl_60_t1 = TR_72 ;
	7'h6b :
		RG_rl_60_t1 = TR_72 ;
	7'h6c :
		RG_rl_60_t1 = TR_72 ;
	7'h6d :
		RG_rl_60_t1 = TR_72 ;
	7'h6e :
		RG_rl_60_t1 = TR_72 ;
	7'h6f :
		RG_rl_60_t1 = TR_72 ;
	7'h70 :
		RG_rl_60_t1 = TR_72 ;
	7'h71 :
		RG_rl_60_t1 = TR_72 ;
	7'h72 :
		RG_rl_60_t1 = TR_72 ;
	7'h73 :
		RG_rl_60_t1 = TR_72 ;
	7'h74 :
		RG_rl_60_t1 = TR_72 ;
	7'h75 :
		RG_rl_60_t1 = TR_72 ;
	7'h76 :
		RG_rl_60_t1 = TR_72 ;
	7'h77 :
		RG_rl_60_t1 = TR_72 ;
	7'h78 :
		RG_rl_60_t1 = TR_72 ;
	7'h79 :
		RG_rl_60_t1 = TR_72 ;
	7'h7a :
		RG_rl_60_t1 = TR_72 ;
	7'h7b :
		RG_rl_60_t1 = TR_72 ;
	7'h7c :
		RG_rl_60_t1 = TR_72 ;
	7'h7d :
		RG_rl_60_t1 = TR_72 ;
	7'h7e :
		RG_rl_60_t1 = TR_72 ;
	7'h7f :
		RG_rl_60_t1 = TR_72 ;
	default :
		RG_rl_60_t1 = 9'hx ;
	endcase
always @ ( RG_rl_60_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_1 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_60_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h3c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_60_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_1 )
		| ( { 9{ U_569 } } & RG_rl_60_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_60_en = ( U_570 | RG_rl_60_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_60_en )
		RG_rl_60 <= RG_rl_60_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_73 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_61_t1 = TR_73 ;
	7'h01 :
		RG_rl_61_t1 = TR_73 ;
	7'h02 :
		RG_rl_61_t1 = TR_73 ;
	7'h03 :
		RG_rl_61_t1 = TR_73 ;
	7'h04 :
		RG_rl_61_t1 = TR_73 ;
	7'h05 :
		RG_rl_61_t1 = TR_73 ;
	7'h06 :
		RG_rl_61_t1 = TR_73 ;
	7'h07 :
		RG_rl_61_t1 = TR_73 ;
	7'h08 :
		RG_rl_61_t1 = TR_73 ;
	7'h09 :
		RG_rl_61_t1 = TR_73 ;
	7'h0a :
		RG_rl_61_t1 = TR_73 ;
	7'h0b :
		RG_rl_61_t1 = TR_73 ;
	7'h0c :
		RG_rl_61_t1 = TR_73 ;
	7'h0d :
		RG_rl_61_t1 = TR_73 ;
	7'h0e :
		RG_rl_61_t1 = TR_73 ;
	7'h0f :
		RG_rl_61_t1 = TR_73 ;
	7'h10 :
		RG_rl_61_t1 = TR_73 ;
	7'h11 :
		RG_rl_61_t1 = TR_73 ;
	7'h12 :
		RG_rl_61_t1 = TR_73 ;
	7'h13 :
		RG_rl_61_t1 = TR_73 ;
	7'h14 :
		RG_rl_61_t1 = TR_73 ;
	7'h15 :
		RG_rl_61_t1 = TR_73 ;
	7'h16 :
		RG_rl_61_t1 = TR_73 ;
	7'h17 :
		RG_rl_61_t1 = TR_73 ;
	7'h18 :
		RG_rl_61_t1 = TR_73 ;
	7'h19 :
		RG_rl_61_t1 = TR_73 ;
	7'h1a :
		RG_rl_61_t1 = TR_73 ;
	7'h1b :
		RG_rl_61_t1 = TR_73 ;
	7'h1c :
		RG_rl_61_t1 = TR_73 ;
	7'h1d :
		RG_rl_61_t1 = TR_73 ;
	7'h1e :
		RG_rl_61_t1 = TR_73 ;
	7'h1f :
		RG_rl_61_t1 = TR_73 ;
	7'h20 :
		RG_rl_61_t1 = TR_73 ;
	7'h21 :
		RG_rl_61_t1 = TR_73 ;
	7'h22 :
		RG_rl_61_t1 = TR_73 ;
	7'h23 :
		RG_rl_61_t1 = TR_73 ;
	7'h24 :
		RG_rl_61_t1 = TR_73 ;
	7'h25 :
		RG_rl_61_t1 = TR_73 ;
	7'h26 :
		RG_rl_61_t1 = TR_73 ;
	7'h27 :
		RG_rl_61_t1 = TR_73 ;
	7'h28 :
		RG_rl_61_t1 = TR_73 ;
	7'h29 :
		RG_rl_61_t1 = TR_73 ;
	7'h2a :
		RG_rl_61_t1 = TR_73 ;
	7'h2b :
		RG_rl_61_t1 = TR_73 ;
	7'h2c :
		RG_rl_61_t1 = TR_73 ;
	7'h2d :
		RG_rl_61_t1 = TR_73 ;
	7'h2e :
		RG_rl_61_t1 = TR_73 ;
	7'h2f :
		RG_rl_61_t1 = TR_73 ;
	7'h30 :
		RG_rl_61_t1 = TR_73 ;
	7'h31 :
		RG_rl_61_t1 = TR_73 ;
	7'h32 :
		RG_rl_61_t1 = TR_73 ;
	7'h33 :
		RG_rl_61_t1 = TR_73 ;
	7'h34 :
		RG_rl_61_t1 = TR_73 ;
	7'h35 :
		RG_rl_61_t1 = TR_73 ;
	7'h36 :
		RG_rl_61_t1 = TR_73 ;
	7'h37 :
		RG_rl_61_t1 = TR_73 ;
	7'h38 :
		RG_rl_61_t1 = TR_73 ;
	7'h39 :
		RG_rl_61_t1 = TR_73 ;
	7'h3a :
		RG_rl_61_t1 = TR_73 ;
	7'h3b :
		RG_rl_61_t1 = TR_73 ;
	7'h3c :
		RG_rl_61_t1 = TR_73 ;
	7'h3d :
		RG_rl_61_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3e :
		RG_rl_61_t1 = TR_73 ;
	7'h3f :
		RG_rl_61_t1 = TR_73 ;
	7'h40 :
		RG_rl_61_t1 = TR_73 ;
	7'h41 :
		RG_rl_61_t1 = TR_73 ;
	7'h42 :
		RG_rl_61_t1 = TR_73 ;
	7'h43 :
		RG_rl_61_t1 = TR_73 ;
	7'h44 :
		RG_rl_61_t1 = TR_73 ;
	7'h45 :
		RG_rl_61_t1 = TR_73 ;
	7'h46 :
		RG_rl_61_t1 = TR_73 ;
	7'h47 :
		RG_rl_61_t1 = TR_73 ;
	7'h48 :
		RG_rl_61_t1 = TR_73 ;
	7'h49 :
		RG_rl_61_t1 = TR_73 ;
	7'h4a :
		RG_rl_61_t1 = TR_73 ;
	7'h4b :
		RG_rl_61_t1 = TR_73 ;
	7'h4c :
		RG_rl_61_t1 = TR_73 ;
	7'h4d :
		RG_rl_61_t1 = TR_73 ;
	7'h4e :
		RG_rl_61_t1 = TR_73 ;
	7'h4f :
		RG_rl_61_t1 = TR_73 ;
	7'h50 :
		RG_rl_61_t1 = TR_73 ;
	7'h51 :
		RG_rl_61_t1 = TR_73 ;
	7'h52 :
		RG_rl_61_t1 = TR_73 ;
	7'h53 :
		RG_rl_61_t1 = TR_73 ;
	7'h54 :
		RG_rl_61_t1 = TR_73 ;
	7'h55 :
		RG_rl_61_t1 = TR_73 ;
	7'h56 :
		RG_rl_61_t1 = TR_73 ;
	7'h57 :
		RG_rl_61_t1 = TR_73 ;
	7'h58 :
		RG_rl_61_t1 = TR_73 ;
	7'h59 :
		RG_rl_61_t1 = TR_73 ;
	7'h5a :
		RG_rl_61_t1 = TR_73 ;
	7'h5b :
		RG_rl_61_t1 = TR_73 ;
	7'h5c :
		RG_rl_61_t1 = TR_73 ;
	7'h5d :
		RG_rl_61_t1 = TR_73 ;
	7'h5e :
		RG_rl_61_t1 = TR_73 ;
	7'h5f :
		RG_rl_61_t1 = TR_73 ;
	7'h60 :
		RG_rl_61_t1 = TR_73 ;
	7'h61 :
		RG_rl_61_t1 = TR_73 ;
	7'h62 :
		RG_rl_61_t1 = TR_73 ;
	7'h63 :
		RG_rl_61_t1 = TR_73 ;
	7'h64 :
		RG_rl_61_t1 = TR_73 ;
	7'h65 :
		RG_rl_61_t1 = TR_73 ;
	7'h66 :
		RG_rl_61_t1 = TR_73 ;
	7'h67 :
		RG_rl_61_t1 = TR_73 ;
	7'h68 :
		RG_rl_61_t1 = TR_73 ;
	7'h69 :
		RG_rl_61_t1 = TR_73 ;
	7'h6a :
		RG_rl_61_t1 = TR_73 ;
	7'h6b :
		RG_rl_61_t1 = TR_73 ;
	7'h6c :
		RG_rl_61_t1 = TR_73 ;
	7'h6d :
		RG_rl_61_t1 = TR_73 ;
	7'h6e :
		RG_rl_61_t1 = TR_73 ;
	7'h6f :
		RG_rl_61_t1 = TR_73 ;
	7'h70 :
		RG_rl_61_t1 = TR_73 ;
	7'h71 :
		RG_rl_61_t1 = TR_73 ;
	7'h72 :
		RG_rl_61_t1 = TR_73 ;
	7'h73 :
		RG_rl_61_t1 = TR_73 ;
	7'h74 :
		RG_rl_61_t1 = TR_73 ;
	7'h75 :
		RG_rl_61_t1 = TR_73 ;
	7'h76 :
		RG_rl_61_t1 = TR_73 ;
	7'h77 :
		RG_rl_61_t1 = TR_73 ;
	7'h78 :
		RG_rl_61_t1 = TR_73 ;
	7'h79 :
		RG_rl_61_t1 = TR_73 ;
	7'h7a :
		RG_rl_61_t1 = TR_73 ;
	7'h7b :
		RG_rl_61_t1 = TR_73 ;
	7'h7c :
		RG_rl_61_t1 = TR_73 ;
	7'h7d :
		RG_rl_61_t1 = TR_73 ;
	7'h7e :
		RG_rl_61_t1 = TR_73 ;
	7'h7f :
		RG_rl_61_t1 = TR_73 ;
	default :
		RG_rl_61_t1 = 9'hx ;
	endcase
always @ ( RG_rl_61_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_2 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_61_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h3d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_61_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_2 )
		| ( { 9{ U_569 } } & RG_rl_61_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_61_en = ( U_570 | RG_rl_61_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_61_en )
		RG_rl_61 <= RG_rl_61_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_74 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_62_t1 = TR_74 ;
	7'h01 :
		RG_rl_62_t1 = TR_74 ;
	7'h02 :
		RG_rl_62_t1 = TR_74 ;
	7'h03 :
		RG_rl_62_t1 = TR_74 ;
	7'h04 :
		RG_rl_62_t1 = TR_74 ;
	7'h05 :
		RG_rl_62_t1 = TR_74 ;
	7'h06 :
		RG_rl_62_t1 = TR_74 ;
	7'h07 :
		RG_rl_62_t1 = TR_74 ;
	7'h08 :
		RG_rl_62_t1 = TR_74 ;
	7'h09 :
		RG_rl_62_t1 = TR_74 ;
	7'h0a :
		RG_rl_62_t1 = TR_74 ;
	7'h0b :
		RG_rl_62_t1 = TR_74 ;
	7'h0c :
		RG_rl_62_t1 = TR_74 ;
	7'h0d :
		RG_rl_62_t1 = TR_74 ;
	7'h0e :
		RG_rl_62_t1 = TR_74 ;
	7'h0f :
		RG_rl_62_t1 = TR_74 ;
	7'h10 :
		RG_rl_62_t1 = TR_74 ;
	7'h11 :
		RG_rl_62_t1 = TR_74 ;
	7'h12 :
		RG_rl_62_t1 = TR_74 ;
	7'h13 :
		RG_rl_62_t1 = TR_74 ;
	7'h14 :
		RG_rl_62_t1 = TR_74 ;
	7'h15 :
		RG_rl_62_t1 = TR_74 ;
	7'h16 :
		RG_rl_62_t1 = TR_74 ;
	7'h17 :
		RG_rl_62_t1 = TR_74 ;
	7'h18 :
		RG_rl_62_t1 = TR_74 ;
	7'h19 :
		RG_rl_62_t1 = TR_74 ;
	7'h1a :
		RG_rl_62_t1 = TR_74 ;
	7'h1b :
		RG_rl_62_t1 = TR_74 ;
	7'h1c :
		RG_rl_62_t1 = TR_74 ;
	7'h1d :
		RG_rl_62_t1 = TR_74 ;
	7'h1e :
		RG_rl_62_t1 = TR_74 ;
	7'h1f :
		RG_rl_62_t1 = TR_74 ;
	7'h20 :
		RG_rl_62_t1 = TR_74 ;
	7'h21 :
		RG_rl_62_t1 = TR_74 ;
	7'h22 :
		RG_rl_62_t1 = TR_74 ;
	7'h23 :
		RG_rl_62_t1 = TR_74 ;
	7'h24 :
		RG_rl_62_t1 = TR_74 ;
	7'h25 :
		RG_rl_62_t1 = TR_74 ;
	7'h26 :
		RG_rl_62_t1 = TR_74 ;
	7'h27 :
		RG_rl_62_t1 = TR_74 ;
	7'h28 :
		RG_rl_62_t1 = TR_74 ;
	7'h29 :
		RG_rl_62_t1 = TR_74 ;
	7'h2a :
		RG_rl_62_t1 = TR_74 ;
	7'h2b :
		RG_rl_62_t1 = TR_74 ;
	7'h2c :
		RG_rl_62_t1 = TR_74 ;
	7'h2d :
		RG_rl_62_t1 = TR_74 ;
	7'h2e :
		RG_rl_62_t1 = TR_74 ;
	7'h2f :
		RG_rl_62_t1 = TR_74 ;
	7'h30 :
		RG_rl_62_t1 = TR_74 ;
	7'h31 :
		RG_rl_62_t1 = TR_74 ;
	7'h32 :
		RG_rl_62_t1 = TR_74 ;
	7'h33 :
		RG_rl_62_t1 = TR_74 ;
	7'h34 :
		RG_rl_62_t1 = TR_74 ;
	7'h35 :
		RG_rl_62_t1 = TR_74 ;
	7'h36 :
		RG_rl_62_t1 = TR_74 ;
	7'h37 :
		RG_rl_62_t1 = TR_74 ;
	7'h38 :
		RG_rl_62_t1 = TR_74 ;
	7'h39 :
		RG_rl_62_t1 = TR_74 ;
	7'h3a :
		RG_rl_62_t1 = TR_74 ;
	7'h3b :
		RG_rl_62_t1 = TR_74 ;
	7'h3c :
		RG_rl_62_t1 = TR_74 ;
	7'h3d :
		RG_rl_62_t1 = TR_74 ;
	7'h3e :
		RG_rl_62_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h3f :
		RG_rl_62_t1 = TR_74 ;
	7'h40 :
		RG_rl_62_t1 = TR_74 ;
	7'h41 :
		RG_rl_62_t1 = TR_74 ;
	7'h42 :
		RG_rl_62_t1 = TR_74 ;
	7'h43 :
		RG_rl_62_t1 = TR_74 ;
	7'h44 :
		RG_rl_62_t1 = TR_74 ;
	7'h45 :
		RG_rl_62_t1 = TR_74 ;
	7'h46 :
		RG_rl_62_t1 = TR_74 ;
	7'h47 :
		RG_rl_62_t1 = TR_74 ;
	7'h48 :
		RG_rl_62_t1 = TR_74 ;
	7'h49 :
		RG_rl_62_t1 = TR_74 ;
	7'h4a :
		RG_rl_62_t1 = TR_74 ;
	7'h4b :
		RG_rl_62_t1 = TR_74 ;
	7'h4c :
		RG_rl_62_t1 = TR_74 ;
	7'h4d :
		RG_rl_62_t1 = TR_74 ;
	7'h4e :
		RG_rl_62_t1 = TR_74 ;
	7'h4f :
		RG_rl_62_t1 = TR_74 ;
	7'h50 :
		RG_rl_62_t1 = TR_74 ;
	7'h51 :
		RG_rl_62_t1 = TR_74 ;
	7'h52 :
		RG_rl_62_t1 = TR_74 ;
	7'h53 :
		RG_rl_62_t1 = TR_74 ;
	7'h54 :
		RG_rl_62_t1 = TR_74 ;
	7'h55 :
		RG_rl_62_t1 = TR_74 ;
	7'h56 :
		RG_rl_62_t1 = TR_74 ;
	7'h57 :
		RG_rl_62_t1 = TR_74 ;
	7'h58 :
		RG_rl_62_t1 = TR_74 ;
	7'h59 :
		RG_rl_62_t1 = TR_74 ;
	7'h5a :
		RG_rl_62_t1 = TR_74 ;
	7'h5b :
		RG_rl_62_t1 = TR_74 ;
	7'h5c :
		RG_rl_62_t1 = TR_74 ;
	7'h5d :
		RG_rl_62_t1 = TR_74 ;
	7'h5e :
		RG_rl_62_t1 = TR_74 ;
	7'h5f :
		RG_rl_62_t1 = TR_74 ;
	7'h60 :
		RG_rl_62_t1 = TR_74 ;
	7'h61 :
		RG_rl_62_t1 = TR_74 ;
	7'h62 :
		RG_rl_62_t1 = TR_74 ;
	7'h63 :
		RG_rl_62_t1 = TR_74 ;
	7'h64 :
		RG_rl_62_t1 = TR_74 ;
	7'h65 :
		RG_rl_62_t1 = TR_74 ;
	7'h66 :
		RG_rl_62_t1 = TR_74 ;
	7'h67 :
		RG_rl_62_t1 = TR_74 ;
	7'h68 :
		RG_rl_62_t1 = TR_74 ;
	7'h69 :
		RG_rl_62_t1 = TR_74 ;
	7'h6a :
		RG_rl_62_t1 = TR_74 ;
	7'h6b :
		RG_rl_62_t1 = TR_74 ;
	7'h6c :
		RG_rl_62_t1 = TR_74 ;
	7'h6d :
		RG_rl_62_t1 = TR_74 ;
	7'h6e :
		RG_rl_62_t1 = TR_74 ;
	7'h6f :
		RG_rl_62_t1 = TR_74 ;
	7'h70 :
		RG_rl_62_t1 = TR_74 ;
	7'h71 :
		RG_rl_62_t1 = TR_74 ;
	7'h72 :
		RG_rl_62_t1 = TR_74 ;
	7'h73 :
		RG_rl_62_t1 = TR_74 ;
	7'h74 :
		RG_rl_62_t1 = TR_74 ;
	7'h75 :
		RG_rl_62_t1 = TR_74 ;
	7'h76 :
		RG_rl_62_t1 = TR_74 ;
	7'h77 :
		RG_rl_62_t1 = TR_74 ;
	7'h78 :
		RG_rl_62_t1 = TR_74 ;
	7'h79 :
		RG_rl_62_t1 = TR_74 ;
	7'h7a :
		RG_rl_62_t1 = TR_74 ;
	7'h7b :
		RG_rl_62_t1 = TR_74 ;
	7'h7c :
		RG_rl_62_t1 = TR_74 ;
	7'h7d :
		RG_rl_62_t1 = TR_74 ;
	7'h7e :
		RG_rl_62_t1 = TR_74 ;
	7'h7f :
		RG_rl_62_t1 = TR_74 ;
	default :
		RG_rl_62_t1 = 9'hx ;
	endcase
always @ ( RG_rl_62_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_3 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_62_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h3e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_62_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_3 )
		| ( { 9{ U_569 } } & RG_rl_62_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_62_en = ( U_570 | RG_rl_62_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_62_en )
		RG_rl_62 <= RG_rl_62_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_75 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_63_t1 = TR_75 ;
	7'h01 :
		RG_rl_63_t1 = TR_75 ;
	7'h02 :
		RG_rl_63_t1 = TR_75 ;
	7'h03 :
		RG_rl_63_t1 = TR_75 ;
	7'h04 :
		RG_rl_63_t1 = TR_75 ;
	7'h05 :
		RG_rl_63_t1 = TR_75 ;
	7'h06 :
		RG_rl_63_t1 = TR_75 ;
	7'h07 :
		RG_rl_63_t1 = TR_75 ;
	7'h08 :
		RG_rl_63_t1 = TR_75 ;
	7'h09 :
		RG_rl_63_t1 = TR_75 ;
	7'h0a :
		RG_rl_63_t1 = TR_75 ;
	7'h0b :
		RG_rl_63_t1 = TR_75 ;
	7'h0c :
		RG_rl_63_t1 = TR_75 ;
	7'h0d :
		RG_rl_63_t1 = TR_75 ;
	7'h0e :
		RG_rl_63_t1 = TR_75 ;
	7'h0f :
		RG_rl_63_t1 = TR_75 ;
	7'h10 :
		RG_rl_63_t1 = TR_75 ;
	7'h11 :
		RG_rl_63_t1 = TR_75 ;
	7'h12 :
		RG_rl_63_t1 = TR_75 ;
	7'h13 :
		RG_rl_63_t1 = TR_75 ;
	7'h14 :
		RG_rl_63_t1 = TR_75 ;
	7'h15 :
		RG_rl_63_t1 = TR_75 ;
	7'h16 :
		RG_rl_63_t1 = TR_75 ;
	7'h17 :
		RG_rl_63_t1 = TR_75 ;
	7'h18 :
		RG_rl_63_t1 = TR_75 ;
	7'h19 :
		RG_rl_63_t1 = TR_75 ;
	7'h1a :
		RG_rl_63_t1 = TR_75 ;
	7'h1b :
		RG_rl_63_t1 = TR_75 ;
	7'h1c :
		RG_rl_63_t1 = TR_75 ;
	7'h1d :
		RG_rl_63_t1 = TR_75 ;
	7'h1e :
		RG_rl_63_t1 = TR_75 ;
	7'h1f :
		RG_rl_63_t1 = TR_75 ;
	7'h20 :
		RG_rl_63_t1 = TR_75 ;
	7'h21 :
		RG_rl_63_t1 = TR_75 ;
	7'h22 :
		RG_rl_63_t1 = TR_75 ;
	7'h23 :
		RG_rl_63_t1 = TR_75 ;
	7'h24 :
		RG_rl_63_t1 = TR_75 ;
	7'h25 :
		RG_rl_63_t1 = TR_75 ;
	7'h26 :
		RG_rl_63_t1 = TR_75 ;
	7'h27 :
		RG_rl_63_t1 = TR_75 ;
	7'h28 :
		RG_rl_63_t1 = TR_75 ;
	7'h29 :
		RG_rl_63_t1 = TR_75 ;
	7'h2a :
		RG_rl_63_t1 = TR_75 ;
	7'h2b :
		RG_rl_63_t1 = TR_75 ;
	7'h2c :
		RG_rl_63_t1 = TR_75 ;
	7'h2d :
		RG_rl_63_t1 = TR_75 ;
	7'h2e :
		RG_rl_63_t1 = TR_75 ;
	7'h2f :
		RG_rl_63_t1 = TR_75 ;
	7'h30 :
		RG_rl_63_t1 = TR_75 ;
	7'h31 :
		RG_rl_63_t1 = TR_75 ;
	7'h32 :
		RG_rl_63_t1 = TR_75 ;
	7'h33 :
		RG_rl_63_t1 = TR_75 ;
	7'h34 :
		RG_rl_63_t1 = TR_75 ;
	7'h35 :
		RG_rl_63_t1 = TR_75 ;
	7'h36 :
		RG_rl_63_t1 = TR_75 ;
	7'h37 :
		RG_rl_63_t1 = TR_75 ;
	7'h38 :
		RG_rl_63_t1 = TR_75 ;
	7'h39 :
		RG_rl_63_t1 = TR_75 ;
	7'h3a :
		RG_rl_63_t1 = TR_75 ;
	7'h3b :
		RG_rl_63_t1 = TR_75 ;
	7'h3c :
		RG_rl_63_t1 = TR_75 ;
	7'h3d :
		RG_rl_63_t1 = TR_75 ;
	7'h3e :
		RG_rl_63_t1 = TR_75 ;
	7'h3f :
		RG_rl_63_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h40 :
		RG_rl_63_t1 = TR_75 ;
	7'h41 :
		RG_rl_63_t1 = TR_75 ;
	7'h42 :
		RG_rl_63_t1 = TR_75 ;
	7'h43 :
		RG_rl_63_t1 = TR_75 ;
	7'h44 :
		RG_rl_63_t1 = TR_75 ;
	7'h45 :
		RG_rl_63_t1 = TR_75 ;
	7'h46 :
		RG_rl_63_t1 = TR_75 ;
	7'h47 :
		RG_rl_63_t1 = TR_75 ;
	7'h48 :
		RG_rl_63_t1 = TR_75 ;
	7'h49 :
		RG_rl_63_t1 = TR_75 ;
	7'h4a :
		RG_rl_63_t1 = TR_75 ;
	7'h4b :
		RG_rl_63_t1 = TR_75 ;
	7'h4c :
		RG_rl_63_t1 = TR_75 ;
	7'h4d :
		RG_rl_63_t1 = TR_75 ;
	7'h4e :
		RG_rl_63_t1 = TR_75 ;
	7'h4f :
		RG_rl_63_t1 = TR_75 ;
	7'h50 :
		RG_rl_63_t1 = TR_75 ;
	7'h51 :
		RG_rl_63_t1 = TR_75 ;
	7'h52 :
		RG_rl_63_t1 = TR_75 ;
	7'h53 :
		RG_rl_63_t1 = TR_75 ;
	7'h54 :
		RG_rl_63_t1 = TR_75 ;
	7'h55 :
		RG_rl_63_t1 = TR_75 ;
	7'h56 :
		RG_rl_63_t1 = TR_75 ;
	7'h57 :
		RG_rl_63_t1 = TR_75 ;
	7'h58 :
		RG_rl_63_t1 = TR_75 ;
	7'h59 :
		RG_rl_63_t1 = TR_75 ;
	7'h5a :
		RG_rl_63_t1 = TR_75 ;
	7'h5b :
		RG_rl_63_t1 = TR_75 ;
	7'h5c :
		RG_rl_63_t1 = TR_75 ;
	7'h5d :
		RG_rl_63_t1 = TR_75 ;
	7'h5e :
		RG_rl_63_t1 = TR_75 ;
	7'h5f :
		RG_rl_63_t1 = TR_75 ;
	7'h60 :
		RG_rl_63_t1 = TR_75 ;
	7'h61 :
		RG_rl_63_t1 = TR_75 ;
	7'h62 :
		RG_rl_63_t1 = TR_75 ;
	7'h63 :
		RG_rl_63_t1 = TR_75 ;
	7'h64 :
		RG_rl_63_t1 = TR_75 ;
	7'h65 :
		RG_rl_63_t1 = TR_75 ;
	7'h66 :
		RG_rl_63_t1 = TR_75 ;
	7'h67 :
		RG_rl_63_t1 = TR_75 ;
	7'h68 :
		RG_rl_63_t1 = TR_75 ;
	7'h69 :
		RG_rl_63_t1 = TR_75 ;
	7'h6a :
		RG_rl_63_t1 = TR_75 ;
	7'h6b :
		RG_rl_63_t1 = TR_75 ;
	7'h6c :
		RG_rl_63_t1 = TR_75 ;
	7'h6d :
		RG_rl_63_t1 = TR_75 ;
	7'h6e :
		RG_rl_63_t1 = TR_75 ;
	7'h6f :
		RG_rl_63_t1 = TR_75 ;
	7'h70 :
		RG_rl_63_t1 = TR_75 ;
	7'h71 :
		RG_rl_63_t1 = TR_75 ;
	7'h72 :
		RG_rl_63_t1 = TR_75 ;
	7'h73 :
		RG_rl_63_t1 = TR_75 ;
	7'h74 :
		RG_rl_63_t1 = TR_75 ;
	7'h75 :
		RG_rl_63_t1 = TR_75 ;
	7'h76 :
		RG_rl_63_t1 = TR_75 ;
	7'h77 :
		RG_rl_63_t1 = TR_75 ;
	7'h78 :
		RG_rl_63_t1 = TR_75 ;
	7'h79 :
		RG_rl_63_t1 = TR_75 ;
	7'h7a :
		RG_rl_63_t1 = TR_75 ;
	7'h7b :
		RG_rl_63_t1 = TR_75 ;
	7'h7c :
		RG_rl_63_t1 = TR_75 ;
	7'h7d :
		RG_rl_63_t1 = TR_75 ;
	7'h7e :
		RG_rl_63_t1 = TR_75 ;
	7'h7f :
		RG_rl_63_t1 = TR_75 ;
	default :
		RG_rl_63_t1 = 9'hx ;
	endcase
always @ ( RG_rl_63_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_4 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_63_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h3f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_63_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_4 )
		| ( { 9{ U_569 } } & RG_rl_63_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_63_en = ( U_570 | RG_rl_63_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_63_en )
		RG_rl_63 <= RG_rl_63_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_76 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_64_t1 = TR_76 ;
	7'h01 :
		RG_rl_64_t1 = TR_76 ;
	7'h02 :
		RG_rl_64_t1 = TR_76 ;
	7'h03 :
		RG_rl_64_t1 = TR_76 ;
	7'h04 :
		RG_rl_64_t1 = TR_76 ;
	7'h05 :
		RG_rl_64_t1 = TR_76 ;
	7'h06 :
		RG_rl_64_t1 = TR_76 ;
	7'h07 :
		RG_rl_64_t1 = TR_76 ;
	7'h08 :
		RG_rl_64_t1 = TR_76 ;
	7'h09 :
		RG_rl_64_t1 = TR_76 ;
	7'h0a :
		RG_rl_64_t1 = TR_76 ;
	7'h0b :
		RG_rl_64_t1 = TR_76 ;
	7'h0c :
		RG_rl_64_t1 = TR_76 ;
	7'h0d :
		RG_rl_64_t1 = TR_76 ;
	7'h0e :
		RG_rl_64_t1 = TR_76 ;
	7'h0f :
		RG_rl_64_t1 = TR_76 ;
	7'h10 :
		RG_rl_64_t1 = TR_76 ;
	7'h11 :
		RG_rl_64_t1 = TR_76 ;
	7'h12 :
		RG_rl_64_t1 = TR_76 ;
	7'h13 :
		RG_rl_64_t1 = TR_76 ;
	7'h14 :
		RG_rl_64_t1 = TR_76 ;
	7'h15 :
		RG_rl_64_t1 = TR_76 ;
	7'h16 :
		RG_rl_64_t1 = TR_76 ;
	7'h17 :
		RG_rl_64_t1 = TR_76 ;
	7'h18 :
		RG_rl_64_t1 = TR_76 ;
	7'h19 :
		RG_rl_64_t1 = TR_76 ;
	7'h1a :
		RG_rl_64_t1 = TR_76 ;
	7'h1b :
		RG_rl_64_t1 = TR_76 ;
	7'h1c :
		RG_rl_64_t1 = TR_76 ;
	7'h1d :
		RG_rl_64_t1 = TR_76 ;
	7'h1e :
		RG_rl_64_t1 = TR_76 ;
	7'h1f :
		RG_rl_64_t1 = TR_76 ;
	7'h20 :
		RG_rl_64_t1 = TR_76 ;
	7'h21 :
		RG_rl_64_t1 = TR_76 ;
	7'h22 :
		RG_rl_64_t1 = TR_76 ;
	7'h23 :
		RG_rl_64_t1 = TR_76 ;
	7'h24 :
		RG_rl_64_t1 = TR_76 ;
	7'h25 :
		RG_rl_64_t1 = TR_76 ;
	7'h26 :
		RG_rl_64_t1 = TR_76 ;
	7'h27 :
		RG_rl_64_t1 = TR_76 ;
	7'h28 :
		RG_rl_64_t1 = TR_76 ;
	7'h29 :
		RG_rl_64_t1 = TR_76 ;
	7'h2a :
		RG_rl_64_t1 = TR_76 ;
	7'h2b :
		RG_rl_64_t1 = TR_76 ;
	7'h2c :
		RG_rl_64_t1 = TR_76 ;
	7'h2d :
		RG_rl_64_t1 = TR_76 ;
	7'h2e :
		RG_rl_64_t1 = TR_76 ;
	7'h2f :
		RG_rl_64_t1 = TR_76 ;
	7'h30 :
		RG_rl_64_t1 = TR_76 ;
	7'h31 :
		RG_rl_64_t1 = TR_76 ;
	7'h32 :
		RG_rl_64_t1 = TR_76 ;
	7'h33 :
		RG_rl_64_t1 = TR_76 ;
	7'h34 :
		RG_rl_64_t1 = TR_76 ;
	7'h35 :
		RG_rl_64_t1 = TR_76 ;
	7'h36 :
		RG_rl_64_t1 = TR_76 ;
	7'h37 :
		RG_rl_64_t1 = TR_76 ;
	7'h38 :
		RG_rl_64_t1 = TR_76 ;
	7'h39 :
		RG_rl_64_t1 = TR_76 ;
	7'h3a :
		RG_rl_64_t1 = TR_76 ;
	7'h3b :
		RG_rl_64_t1 = TR_76 ;
	7'h3c :
		RG_rl_64_t1 = TR_76 ;
	7'h3d :
		RG_rl_64_t1 = TR_76 ;
	7'h3e :
		RG_rl_64_t1 = TR_76 ;
	7'h3f :
		RG_rl_64_t1 = TR_76 ;
	7'h40 :
		RG_rl_64_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h41 :
		RG_rl_64_t1 = TR_76 ;
	7'h42 :
		RG_rl_64_t1 = TR_76 ;
	7'h43 :
		RG_rl_64_t1 = TR_76 ;
	7'h44 :
		RG_rl_64_t1 = TR_76 ;
	7'h45 :
		RG_rl_64_t1 = TR_76 ;
	7'h46 :
		RG_rl_64_t1 = TR_76 ;
	7'h47 :
		RG_rl_64_t1 = TR_76 ;
	7'h48 :
		RG_rl_64_t1 = TR_76 ;
	7'h49 :
		RG_rl_64_t1 = TR_76 ;
	7'h4a :
		RG_rl_64_t1 = TR_76 ;
	7'h4b :
		RG_rl_64_t1 = TR_76 ;
	7'h4c :
		RG_rl_64_t1 = TR_76 ;
	7'h4d :
		RG_rl_64_t1 = TR_76 ;
	7'h4e :
		RG_rl_64_t1 = TR_76 ;
	7'h4f :
		RG_rl_64_t1 = TR_76 ;
	7'h50 :
		RG_rl_64_t1 = TR_76 ;
	7'h51 :
		RG_rl_64_t1 = TR_76 ;
	7'h52 :
		RG_rl_64_t1 = TR_76 ;
	7'h53 :
		RG_rl_64_t1 = TR_76 ;
	7'h54 :
		RG_rl_64_t1 = TR_76 ;
	7'h55 :
		RG_rl_64_t1 = TR_76 ;
	7'h56 :
		RG_rl_64_t1 = TR_76 ;
	7'h57 :
		RG_rl_64_t1 = TR_76 ;
	7'h58 :
		RG_rl_64_t1 = TR_76 ;
	7'h59 :
		RG_rl_64_t1 = TR_76 ;
	7'h5a :
		RG_rl_64_t1 = TR_76 ;
	7'h5b :
		RG_rl_64_t1 = TR_76 ;
	7'h5c :
		RG_rl_64_t1 = TR_76 ;
	7'h5d :
		RG_rl_64_t1 = TR_76 ;
	7'h5e :
		RG_rl_64_t1 = TR_76 ;
	7'h5f :
		RG_rl_64_t1 = TR_76 ;
	7'h60 :
		RG_rl_64_t1 = TR_76 ;
	7'h61 :
		RG_rl_64_t1 = TR_76 ;
	7'h62 :
		RG_rl_64_t1 = TR_76 ;
	7'h63 :
		RG_rl_64_t1 = TR_76 ;
	7'h64 :
		RG_rl_64_t1 = TR_76 ;
	7'h65 :
		RG_rl_64_t1 = TR_76 ;
	7'h66 :
		RG_rl_64_t1 = TR_76 ;
	7'h67 :
		RG_rl_64_t1 = TR_76 ;
	7'h68 :
		RG_rl_64_t1 = TR_76 ;
	7'h69 :
		RG_rl_64_t1 = TR_76 ;
	7'h6a :
		RG_rl_64_t1 = TR_76 ;
	7'h6b :
		RG_rl_64_t1 = TR_76 ;
	7'h6c :
		RG_rl_64_t1 = TR_76 ;
	7'h6d :
		RG_rl_64_t1 = TR_76 ;
	7'h6e :
		RG_rl_64_t1 = TR_76 ;
	7'h6f :
		RG_rl_64_t1 = TR_76 ;
	7'h70 :
		RG_rl_64_t1 = TR_76 ;
	7'h71 :
		RG_rl_64_t1 = TR_76 ;
	7'h72 :
		RG_rl_64_t1 = TR_76 ;
	7'h73 :
		RG_rl_64_t1 = TR_76 ;
	7'h74 :
		RG_rl_64_t1 = TR_76 ;
	7'h75 :
		RG_rl_64_t1 = TR_76 ;
	7'h76 :
		RG_rl_64_t1 = TR_76 ;
	7'h77 :
		RG_rl_64_t1 = TR_76 ;
	7'h78 :
		RG_rl_64_t1 = TR_76 ;
	7'h79 :
		RG_rl_64_t1 = TR_76 ;
	7'h7a :
		RG_rl_64_t1 = TR_76 ;
	7'h7b :
		RG_rl_64_t1 = TR_76 ;
	7'h7c :
		RG_rl_64_t1 = TR_76 ;
	7'h7d :
		RG_rl_64_t1 = TR_76 ;
	7'h7e :
		RG_rl_64_t1 = TR_76 ;
	7'h7f :
		RG_rl_64_t1 = TR_76 ;
	default :
		RG_rl_64_t1 = 9'hx ;
	endcase
always @ ( RG_rl_64_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_5 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_64_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h40 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_64_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_5 )
		| ( { 9{ U_569 } } & RG_rl_64_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_64_en = ( U_570 | RG_rl_64_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_64_en )
		RG_rl_64 <= RG_rl_64_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_77 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_65_t1 = TR_77 ;
	7'h01 :
		RG_rl_65_t1 = TR_77 ;
	7'h02 :
		RG_rl_65_t1 = TR_77 ;
	7'h03 :
		RG_rl_65_t1 = TR_77 ;
	7'h04 :
		RG_rl_65_t1 = TR_77 ;
	7'h05 :
		RG_rl_65_t1 = TR_77 ;
	7'h06 :
		RG_rl_65_t1 = TR_77 ;
	7'h07 :
		RG_rl_65_t1 = TR_77 ;
	7'h08 :
		RG_rl_65_t1 = TR_77 ;
	7'h09 :
		RG_rl_65_t1 = TR_77 ;
	7'h0a :
		RG_rl_65_t1 = TR_77 ;
	7'h0b :
		RG_rl_65_t1 = TR_77 ;
	7'h0c :
		RG_rl_65_t1 = TR_77 ;
	7'h0d :
		RG_rl_65_t1 = TR_77 ;
	7'h0e :
		RG_rl_65_t1 = TR_77 ;
	7'h0f :
		RG_rl_65_t1 = TR_77 ;
	7'h10 :
		RG_rl_65_t1 = TR_77 ;
	7'h11 :
		RG_rl_65_t1 = TR_77 ;
	7'h12 :
		RG_rl_65_t1 = TR_77 ;
	7'h13 :
		RG_rl_65_t1 = TR_77 ;
	7'h14 :
		RG_rl_65_t1 = TR_77 ;
	7'h15 :
		RG_rl_65_t1 = TR_77 ;
	7'h16 :
		RG_rl_65_t1 = TR_77 ;
	7'h17 :
		RG_rl_65_t1 = TR_77 ;
	7'h18 :
		RG_rl_65_t1 = TR_77 ;
	7'h19 :
		RG_rl_65_t1 = TR_77 ;
	7'h1a :
		RG_rl_65_t1 = TR_77 ;
	7'h1b :
		RG_rl_65_t1 = TR_77 ;
	7'h1c :
		RG_rl_65_t1 = TR_77 ;
	7'h1d :
		RG_rl_65_t1 = TR_77 ;
	7'h1e :
		RG_rl_65_t1 = TR_77 ;
	7'h1f :
		RG_rl_65_t1 = TR_77 ;
	7'h20 :
		RG_rl_65_t1 = TR_77 ;
	7'h21 :
		RG_rl_65_t1 = TR_77 ;
	7'h22 :
		RG_rl_65_t1 = TR_77 ;
	7'h23 :
		RG_rl_65_t1 = TR_77 ;
	7'h24 :
		RG_rl_65_t1 = TR_77 ;
	7'h25 :
		RG_rl_65_t1 = TR_77 ;
	7'h26 :
		RG_rl_65_t1 = TR_77 ;
	7'h27 :
		RG_rl_65_t1 = TR_77 ;
	7'h28 :
		RG_rl_65_t1 = TR_77 ;
	7'h29 :
		RG_rl_65_t1 = TR_77 ;
	7'h2a :
		RG_rl_65_t1 = TR_77 ;
	7'h2b :
		RG_rl_65_t1 = TR_77 ;
	7'h2c :
		RG_rl_65_t1 = TR_77 ;
	7'h2d :
		RG_rl_65_t1 = TR_77 ;
	7'h2e :
		RG_rl_65_t1 = TR_77 ;
	7'h2f :
		RG_rl_65_t1 = TR_77 ;
	7'h30 :
		RG_rl_65_t1 = TR_77 ;
	7'h31 :
		RG_rl_65_t1 = TR_77 ;
	7'h32 :
		RG_rl_65_t1 = TR_77 ;
	7'h33 :
		RG_rl_65_t1 = TR_77 ;
	7'h34 :
		RG_rl_65_t1 = TR_77 ;
	7'h35 :
		RG_rl_65_t1 = TR_77 ;
	7'h36 :
		RG_rl_65_t1 = TR_77 ;
	7'h37 :
		RG_rl_65_t1 = TR_77 ;
	7'h38 :
		RG_rl_65_t1 = TR_77 ;
	7'h39 :
		RG_rl_65_t1 = TR_77 ;
	7'h3a :
		RG_rl_65_t1 = TR_77 ;
	7'h3b :
		RG_rl_65_t1 = TR_77 ;
	7'h3c :
		RG_rl_65_t1 = TR_77 ;
	7'h3d :
		RG_rl_65_t1 = TR_77 ;
	7'h3e :
		RG_rl_65_t1 = TR_77 ;
	7'h3f :
		RG_rl_65_t1 = TR_77 ;
	7'h40 :
		RG_rl_65_t1 = TR_77 ;
	7'h41 :
		RG_rl_65_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h42 :
		RG_rl_65_t1 = TR_77 ;
	7'h43 :
		RG_rl_65_t1 = TR_77 ;
	7'h44 :
		RG_rl_65_t1 = TR_77 ;
	7'h45 :
		RG_rl_65_t1 = TR_77 ;
	7'h46 :
		RG_rl_65_t1 = TR_77 ;
	7'h47 :
		RG_rl_65_t1 = TR_77 ;
	7'h48 :
		RG_rl_65_t1 = TR_77 ;
	7'h49 :
		RG_rl_65_t1 = TR_77 ;
	7'h4a :
		RG_rl_65_t1 = TR_77 ;
	7'h4b :
		RG_rl_65_t1 = TR_77 ;
	7'h4c :
		RG_rl_65_t1 = TR_77 ;
	7'h4d :
		RG_rl_65_t1 = TR_77 ;
	7'h4e :
		RG_rl_65_t1 = TR_77 ;
	7'h4f :
		RG_rl_65_t1 = TR_77 ;
	7'h50 :
		RG_rl_65_t1 = TR_77 ;
	7'h51 :
		RG_rl_65_t1 = TR_77 ;
	7'h52 :
		RG_rl_65_t1 = TR_77 ;
	7'h53 :
		RG_rl_65_t1 = TR_77 ;
	7'h54 :
		RG_rl_65_t1 = TR_77 ;
	7'h55 :
		RG_rl_65_t1 = TR_77 ;
	7'h56 :
		RG_rl_65_t1 = TR_77 ;
	7'h57 :
		RG_rl_65_t1 = TR_77 ;
	7'h58 :
		RG_rl_65_t1 = TR_77 ;
	7'h59 :
		RG_rl_65_t1 = TR_77 ;
	7'h5a :
		RG_rl_65_t1 = TR_77 ;
	7'h5b :
		RG_rl_65_t1 = TR_77 ;
	7'h5c :
		RG_rl_65_t1 = TR_77 ;
	7'h5d :
		RG_rl_65_t1 = TR_77 ;
	7'h5e :
		RG_rl_65_t1 = TR_77 ;
	7'h5f :
		RG_rl_65_t1 = TR_77 ;
	7'h60 :
		RG_rl_65_t1 = TR_77 ;
	7'h61 :
		RG_rl_65_t1 = TR_77 ;
	7'h62 :
		RG_rl_65_t1 = TR_77 ;
	7'h63 :
		RG_rl_65_t1 = TR_77 ;
	7'h64 :
		RG_rl_65_t1 = TR_77 ;
	7'h65 :
		RG_rl_65_t1 = TR_77 ;
	7'h66 :
		RG_rl_65_t1 = TR_77 ;
	7'h67 :
		RG_rl_65_t1 = TR_77 ;
	7'h68 :
		RG_rl_65_t1 = TR_77 ;
	7'h69 :
		RG_rl_65_t1 = TR_77 ;
	7'h6a :
		RG_rl_65_t1 = TR_77 ;
	7'h6b :
		RG_rl_65_t1 = TR_77 ;
	7'h6c :
		RG_rl_65_t1 = TR_77 ;
	7'h6d :
		RG_rl_65_t1 = TR_77 ;
	7'h6e :
		RG_rl_65_t1 = TR_77 ;
	7'h6f :
		RG_rl_65_t1 = TR_77 ;
	7'h70 :
		RG_rl_65_t1 = TR_77 ;
	7'h71 :
		RG_rl_65_t1 = TR_77 ;
	7'h72 :
		RG_rl_65_t1 = TR_77 ;
	7'h73 :
		RG_rl_65_t1 = TR_77 ;
	7'h74 :
		RG_rl_65_t1 = TR_77 ;
	7'h75 :
		RG_rl_65_t1 = TR_77 ;
	7'h76 :
		RG_rl_65_t1 = TR_77 ;
	7'h77 :
		RG_rl_65_t1 = TR_77 ;
	7'h78 :
		RG_rl_65_t1 = TR_77 ;
	7'h79 :
		RG_rl_65_t1 = TR_77 ;
	7'h7a :
		RG_rl_65_t1 = TR_77 ;
	7'h7b :
		RG_rl_65_t1 = TR_77 ;
	7'h7c :
		RG_rl_65_t1 = TR_77 ;
	7'h7d :
		RG_rl_65_t1 = TR_77 ;
	7'h7e :
		RG_rl_65_t1 = TR_77 ;
	7'h7f :
		RG_rl_65_t1 = TR_77 ;
	default :
		RG_rl_65_t1 = 9'hx ;
	endcase
always @ ( RG_rl_65_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_6 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_65_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h41 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_65_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_6 )
		| ( { 9{ U_569 } } & RG_rl_65_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_65_en = ( U_570 | RG_rl_65_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_65_en )
		RG_rl_65 <= RG_rl_65_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_78 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_66_t1 = TR_78 ;
	7'h01 :
		RG_rl_66_t1 = TR_78 ;
	7'h02 :
		RG_rl_66_t1 = TR_78 ;
	7'h03 :
		RG_rl_66_t1 = TR_78 ;
	7'h04 :
		RG_rl_66_t1 = TR_78 ;
	7'h05 :
		RG_rl_66_t1 = TR_78 ;
	7'h06 :
		RG_rl_66_t1 = TR_78 ;
	7'h07 :
		RG_rl_66_t1 = TR_78 ;
	7'h08 :
		RG_rl_66_t1 = TR_78 ;
	7'h09 :
		RG_rl_66_t1 = TR_78 ;
	7'h0a :
		RG_rl_66_t1 = TR_78 ;
	7'h0b :
		RG_rl_66_t1 = TR_78 ;
	7'h0c :
		RG_rl_66_t1 = TR_78 ;
	7'h0d :
		RG_rl_66_t1 = TR_78 ;
	7'h0e :
		RG_rl_66_t1 = TR_78 ;
	7'h0f :
		RG_rl_66_t1 = TR_78 ;
	7'h10 :
		RG_rl_66_t1 = TR_78 ;
	7'h11 :
		RG_rl_66_t1 = TR_78 ;
	7'h12 :
		RG_rl_66_t1 = TR_78 ;
	7'h13 :
		RG_rl_66_t1 = TR_78 ;
	7'h14 :
		RG_rl_66_t1 = TR_78 ;
	7'h15 :
		RG_rl_66_t1 = TR_78 ;
	7'h16 :
		RG_rl_66_t1 = TR_78 ;
	7'h17 :
		RG_rl_66_t1 = TR_78 ;
	7'h18 :
		RG_rl_66_t1 = TR_78 ;
	7'h19 :
		RG_rl_66_t1 = TR_78 ;
	7'h1a :
		RG_rl_66_t1 = TR_78 ;
	7'h1b :
		RG_rl_66_t1 = TR_78 ;
	7'h1c :
		RG_rl_66_t1 = TR_78 ;
	7'h1d :
		RG_rl_66_t1 = TR_78 ;
	7'h1e :
		RG_rl_66_t1 = TR_78 ;
	7'h1f :
		RG_rl_66_t1 = TR_78 ;
	7'h20 :
		RG_rl_66_t1 = TR_78 ;
	7'h21 :
		RG_rl_66_t1 = TR_78 ;
	7'h22 :
		RG_rl_66_t1 = TR_78 ;
	7'h23 :
		RG_rl_66_t1 = TR_78 ;
	7'h24 :
		RG_rl_66_t1 = TR_78 ;
	7'h25 :
		RG_rl_66_t1 = TR_78 ;
	7'h26 :
		RG_rl_66_t1 = TR_78 ;
	7'h27 :
		RG_rl_66_t1 = TR_78 ;
	7'h28 :
		RG_rl_66_t1 = TR_78 ;
	7'h29 :
		RG_rl_66_t1 = TR_78 ;
	7'h2a :
		RG_rl_66_t1 = TR_78 ;
	7'h2b :
		RG_rl_66_t1 = TR_78 ;
	7'h2c :
		RG_rl_66_t1 = TR_78 ;
	7'h2d :
		RG_rl_66_t1 = TR_78 ;
	7'h2e :
		RG_rl_66_t1 = TR_78 ;
	7'h2f :
		RG_rl_66_t1 = TR_78 ;
	7'h30 :
		RG_rl_66_t1 = TR_78 ;
	7'h31 :
		RG_rl_66_t1 = TR_78 ;
	7'h32 :
		RG_rl_66_t1 = TR_78 ;
	7'h33 :
		RG_rl_66_t1 = TR_78 ;
	7'h34 :
		RG_rl_66_t1 = TR_78 ;
	7'h35 :
		RG_rl_66_t1 = TR_78 ;
	7'h36 :
		RG_rl_66_t1 = TR_78 ;
	7'h37 :
		RG_rl_66_t1 = TR_78 ;
	7'h38 :
		RG_rl_66_t1 = TR_78 ;
	7'h39 :
		RG_rl_66_t1 = TR_78 ;
	7'h3a :
		RG_rl_66_t1 = TR_78 ;
	7'h3b :
		RG_rl_66_t1 = TR_78 ;
	7'h3c :
		RG_rl_66_t1 = TR_78 ;
	7'h3d :
		RG_rl_66_t1 = TR_78 ;
	7'h3e :
		RG_rl_66_t1 = TR_78 ;
	7'h3f :
		RG_rl_66_t1 = TR_78 ;
	7'h40 :
		RG_rl_66_t1 = TR_78 ;
	7'h41 :
		RG_rl_66_t1 = TR_78 ;
	7'h42 :
		RG_rl_66_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h43 :
		RG_rl_66_t1 = TR_78 ;
	7'h44 :
		RG_rl_66_t1 = TR_78 ;
	7'h45 :
		RG_rl_66_t1 = TR_78 ;
	7'h46 :
		RG_rl_66_t1 = TR_78 ;
	7'h47 :
		RG_rl_66_t1 = TR_78 ;
	7'h48 :
		RG_rl_66_t1 = TR_78 ;
	7'h49 :
		RG_rl_66_t1 = TR_78 ;
	7'h4a :
		RG_rl_66_t1 = TR_78 ;
	7'h4b :
		RG_rl_66_t1 = TR_78 ;
	7'h4c :
		RG_rl_66_t1 = TR_78 ;
	7'h4d :
		RG_rl_66_t1 = TR_78 ;
	7'h4e :
		RG_rl_66_t1 = TR_78 ;
	7'h4f :
		RG_rl_66_t1 = TR_78 ;
	7'h50 :
		RG_rl_66_t1 = TR_78 ;
	7'h51 :
		RG_rl_66_t1 = TR_78 ;
	7'h52 :
		RG_rl_66_t1 = TR_78 ;
	7'h53 :
		RG_rl_66_t1 = TR_78 ;
	7'h54 :
		RG_rl_66_t1 = TR_78 ;
	7'h55 :
		RG_rl_66_t1 = TR_78 ;
	7'h56 :
		RG_rl_66_t1 = TR_78 ;
	7'h57 :
		RG_rl_66_t1 = TR_78 ;
	7'h58 :
		RG_rl_66_t1 = TR_78 ;
	7'h59 :
		RG_rl_66_t1 = TR_78 ;
	7'h5a :
		RG_rl_66_t1 = TR_78 ;
	7'h5b :
		RG_rl_66_t1 = TR_78 ;
	7'h5c :
		RG_rl_66_t1 = TR_78 ;
	7'h5d :
		RG_rl_66_t1 = TR_78 ;
	7'h5e :
		RG_rl_66_t1 = TR_78 ;
	7'h5f :
		RG_rl_66_t1 = TR_78 ;
	7'h60 :
		RG_rl_66_t1 = TR_78 ;
	7'h61 :
		RG_rl_66_t1 = TR_78 ;
	7'h62 :
		RG_rl_66_t1 = TR_78 ;
	7'h63 :
		RG_rl_66_t1 = TR_78 ;
	7'h64 :
		RG_rl_66_t1 = TR_78 ;
	7'h65 :
		RG_rl_66_t1 = TR_78 ;
	7'h66 :
		RG_rl_66_t1 = TR_78 ;
	7'h67 :
		RG_rl_66_t1 = TR_78 ;
	7'h68 :
		RG_rl_66_t1 = TR_78 ;
	7'h69 :
		RG_rl_66_t1 = TR_78 ;
	7'h6a :
		RG_rl_66_t1 = TR_78 ;
	7'h6b :
		RG_rl_66_t1 = TR_78 ;
	7'h6c :
		RG_rl_66_t1 = TR_78 ;
	7'h6d :
		RG_rl_66_t1 = TR_78 ;
	7'h6e :
		RG_rl_66_t1 = TR_78 ;
	7'h6f :
		RG_rl_66_t1 = TR_78 ;
	7'h70 :
		RG_rl_66_t1 = TR_78 ;
	7'h71 :
		RG_rl_66_t1 = TR_78 ;
	7'h72 :
		RG_rl_66_t1 = TR_78 ;
	7'h73 :
		RG_rl_66_t1 = TR_78 ;
	7'h74 :
		RG_rl_66_t1 = TR_78 ;
	7'h75 :
		RG_rl_66_t1 = TR_78 ;
	7'h76 :
		RG_rl_66_t1 = TR_78 ;
	7'h77 :
		RG_rl_66_t1 = TR_78 ;
	7'h78 :
		RG_rl_66_t1 = TR_78 ;
	7'h79 :
		RG_rl_66_t1 = TR_78 ;
	7'h7a :
		RG_rl_66_t1 = TR_78 ;
	7'h7b :
		RG_rl_66_t1 = TR_78 ;
	7'h7c :
		RG_rl_66_t1 = TR_78 ;
	7'h7d :
		RG_rl_66_t1 = TR_78 ;
	7'h7e :
		RG_rl_66_t1 = TR_78 ;
	7'h7f :
		RG_rl_66_t1 = TR_78 ;
	default :
		RG_rl_66_t1 = 9'hx ;
	endcase
always @ ( RG_rl_66_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_7 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_66_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h42 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_66_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_7 )
		| ( { 9{ U_569 } } & RG_rl_66_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_66_en = ( U_570 | RG_rl_66_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_66_en )
		RG_rl_66 <= RG_rl_66_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_79 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_67_t1 = TR_79 ;
	7'h01 :
		RG_rl_67_t1 = TR_79 ;
	7'h02 :
		RG_rl_67_t1 = TR_79 ;
	7'h03 :
		RG_rl_67_t1 = TR_79 ;
	7'h04 :
		RG_rl_67_t1 = TR_79 ;
	7'h05 :
		RG_rl_67_t1 = TR_79 ;
	7'h06 :
		RG_rl_67_t1 = TR_79 ;
	7'h07 :
		RG_rl_67_t1 = TR_79 ;
	7'h08 :
		RG_rl_67_t1 = TR_79 ;
	7'h09 :
		RG_rl_67_t1 = TR_79 ;
	7'h0a :
		RG_rl_67_t1 = TR_79 ;
	7'h0b :
		RG_rl_67_t1 = TR_79 ;
	7'h0c :
		RG_rl_67_t1 = TR_79 ;
	7'h0d :
		RG_rl_67_t1 = TR_79 ;
	7'h0e :
		RG_rl_67_t1 = TR_79 ;
	7'h0f :
		RG_rl_67_t1 = TR_79 ;
	7'h10 :
		RG_rl_67_t1 = TR_79 ;
	7'h11 :
		RG_rl_67_t1 = TR_79 ;
	7'h12 :
		RG_rl_67_t1 = TR_79 ;
	7'h13 :
		RG_rl_67_t1 = TR_79 ;
	7'h14 :
		RG_rl_67_t1 = TR_79 ;
	7'h15 :
		RG_rl_67_t1 = TR_79 ;
	7'h16 :
		RG_rl_67_t1 = TR_79 ;
	7'h17 :
		RG_rl_67_t1 = TR_79 ;
	7'h18 :
		RG_rl_67_t1 = TR_79 ;
	7'h19 :
		RG_rl_67_t1 = TR_79 ;
	7'h1a :
		RG_rl_67_t1 = TR_79 ;
	7'h1b :
		RG_rl_67_t1 = TR_79 ;
	7'h1c :
		RG_rl_67_t1 = TR_79 ;
	7'h1d :
		RG_rl_67_t1 = TR_79 ;
	7'h1e :
		RG_rl_67_t1 = TR_79 ;
	7'h1f :
		RG_rl_67_t1 = TR_79 ;
	7'h20 :
		RG_rl_67_t1 = TR_79 ;
	7'h21 :
		RG_rl_67_t1 = TR_79 ;
	7'h22 :
		RG_rl_67_t1 = TR_79 ;
	7'h23 :
		RG_rl_67_t1 = TR_79 ;
	7'h24 :
		RG_rl_67_t1 = TR_79 ;
	7'h25 :
		RG_rl_67_t1 = TR_79 ;
	7'h26 :
		RG_rl_67_t1 = TR_79 ;
	7'h27 :
		RG_rl_67_t1 = TR_79 ;
	7'h28 :
		RG_rl_67_t1 = TR_79 ;
	7'h29 :
		RG_rl_67_t1 = TR_79 ;
	7'h2a :
		RG_rl_67_t1 = TR_79 ;
	7'h2b :
		RG_rl_67_t1 = TR_79 ;
	7'h2c :
		RG_rl_67_t1 = TR_79 ;
	7'h2d :
		RG_rl_67_t1 = TR_79 ;
	7'h2e :
		RG_rl_67_t1 = TR_79 ;
	7'h2f :
		RG_rl_67_t1 = TR_79 ;
	7'h30 :
		RG_rl_67_t1 = TR_79 ;
	7'h31 :
		RG_rl_67_t1 = TR_79 ;
	7'h32 :
		RG_rl_67_t1 = TR_79 ;
	7'h33 :
		RG_rl_67_t1 = TR_79 ;
	7'h34 :
		RG_rl_67_t1 = TR_79 ;
	7'h35 :
		RG_rl_67_t1 = TR_79 ;
	7'h36 :
		RG_rl_67_t1 = TR_79 ;
	7'h37 :
		RG_rl_67_t1 = TR_79 ;
	7'h38 :
		RG_rl_67_t1 = TR_79 ;
	7'h39 :
		RG_rl_67_t1 = TR_79 ;
	7'h3a :
		RG_rl_67_t1 = TR_79 ;
	7'h3b :
		RG_rl_67_t1 = TR_79 ;
	7'h3c :
		RG_rl_67_t1 = TR_79 ;
	7'h3d :
		RG_rl_67_t1 = TR_79 ;
	7'h3e :
		RG_rl_67_t1 = TR_79 ;
	7'h3f :
		RG_rl_67_t1 = TR_79 ;
	7'h40 :
		RG_rl_67_t1 = TR_79 ;
	7'h41 :
		RG_rl_67_t1 = TR_79 ;
	7'h42 :
		RG_rl_67_t1 = TR_79 ;
	7'h43 :
		RG_rl_67_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h44 :
		RG_rl_67_t1 = TR_79 ;
	7'h45 :
		RG_rl_67_t1 = TR_79 ;
	7'h46 :
		RG_rl_67_t1 = TR_79 ;
	7'h47 :
		RG_rl_67_t1 = TR_79 ;
	7'h48 :
		RG_rl_67_t1 = TR_79 ;
	7'h49 :
		RG_rl_67_t1 = TR_79 ;
	7'h4a :
		RG_rl_67_t1 = TR_79 ;
	7'h4b :
		RG_rl_67_t1 = TR_79 ;
	7'h4c :
		RG_rl_67_t1 = TR_79 ;
	7'h4d :
		RG_rl_67_t1 = TR_79 ;
	7'h4e :
		RG_rl_67_t1 = TR_79 ;
	7'h4f :
		RG_rl_67_t1 = TR_79 ;
	7'h50 :
		RG_rl_67_t1 = TR_79 ;
	7'h51 :
		RG_rl_67_t1 = TR_79 ;
	7'h52 :
		RG_rl_67_t1 = TR_79 ;
	7'h53 :
		RG_rl_67_t1 = TR_79 ;
	7'h54 :
		RG_rl_67_t1 = TR_79 ;
	7'h55 :
		RG_rl_67_t1 = TR_79 ;
	7'h56 :
		RG_rl_67_t1 = TR_79 ;
	7'h57 :
		RG_rl_67_t1 = TR_79 ;
	7'h58 :
		RG_rl_67_t1 = TR_79 ;
	7'h59 :
		RG_rl_67_t1 = TR_79 ;
	7'h5a :
		RG_rl_67_t1 = TR_79 ;
	7'h5b :
		RG_rl_67_t1 = TR_79 ;
	7'h5c :
		RG_rl_67_t1 = TR_79 ;
	7'h5d :
		RG_rl_67_t1 = TR_79 ;
	7'h5e :
		RG_rl_67_t1 = TR_79 ;
	7'h5f :
		RG_rl_67_t1 = TR_79 ;
	7'h60 :
		RG_rl_67_t1 = TR_79 ;
	7'h61 :
		RG_rl_67_t1 = TR_79 ;
	7'h62 :
		RG_rl_67_t1 = TR_79 ;
	7'h63 :
		RG_rl_67_t1 = TR_79 ;
	7'h64 :
		RG_rl_67_t1 = TR_79 ;
	7'h65 :
		RG_rl_67_t1 = TR_79 ;
	7'h66 :
		RG_rl_67_t1 = TR_79 ;
	7'h67 :
		RG_rl_67_t1 = TR_79 ;
	7'h68 :
		RG_rl_67_t1 = TR_79 ;
	7'h69 :
		RG_rl_67_t1 = TR_79 ;
	7'h6a :
		RG_rl_67_t1 = TR_79 ;
	7'h6b :
		RG_rl_67_t1 = TR_79 ;
	7'h6c :
		RG_rl_67_t1 = TR_79 ;
	7'h6d :
		RG_rl_67_t1 = TR_79 ;
	7'h6e :
		RG_rl_67_t1 = TR_79 ;
	7'h6f :
		RG_rl_67_t1 = TR_79 ;
	7'h70 :
		RG_rl_67_t1 = TR_79 ;
	7'h71 :
		RG_rl_67_t1 = TR_79 ;
	7'h72 :
		RG_rl_67_t1 = TR_79 ;
	7'h73 :
		RG_rl_67_t1 = TR_79 ;
	7'h74 :
		RG_rl_67_t1 = TR_79 ;
	7'h75 :
		RG_rl_67_t1 = TR_79 ;
	7'h76 :
		RG_rl_67_t1 = TR_79 ;
	7'h77 :
		RG_rl_67_t1 = TR_79 ;
	7'h78 :
		RG_rl_67_t1 = TR_79 ;
	7'h79 :
		RG_rl_67_t1 = TR_79 ;
	7'h7a :
		RG_rl_67_t1 = TR_79 ;
	7'h7b :
		RG_rl_67_t1 = TR_79 ;
	7'h7c :
		RG_rl_67_t1 = TR_79 ;
	7'h7d :
		RG_rl_67_t1 = TR_79 ;
	7'h7e :
		RG_rl_67_t1 = TR_79 ;
	7'h7f :
		RG_rl_67_t1 = TR_79 ;
	default :
		RG_rl_67_t1 = 9'hx ;
	endcase
always @ ( RG_rl_67_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_8 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_67_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h43 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_67_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_8 )
		| ( { 9{ U_569 } } & RG_rl_67_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_67_en = ( U_570 | RG_rl_67_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_67_en )
		RG_rl_67 <= RG_rl_67_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_80 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_68_t1 = TR_80 ;
	7'h01 :
		RG_rl_68_t1 = TR_80 ;
	7'h02 :
		RG_rl_68_t1 = TR_80 ;
	7'h03 :
		RG_rl_68_t1 = TR_80 ;
	7'h04 :
		RG_rl_68_t1 = TR_80 ;
	7'h05 :
		RG_rl_68_t1 = TR_80 ;
	7'h06 :
		RG_rl_68_t1 = TR_80 ;
	7'h07 :
		RG_rl_68_t1 = TR_80 ;
	7'h08 :
		RG_rl_68_t1 = TR_80 ;
	7'h09 :
		RG_rl_68_t1 = TR_80 ;
	7'h0a :
		RG_rl_68_t1 = TR_80 ;
	7'h0b :
		RG_rl_68_t1 = TR_80 ;
	7'h0c :
		RG_rl_68_t1 = TR_80 ;
	7'h0d :
		RG_rl_68_t1 = TR_80 ;
	7'h0e :
		RG_rl_68_t1 = TR_80 ;
	7'h0f :
		RG_rl_68_t1 = TR_80 ;
	7'h10 :
		RG_rl_68_t1 = TR_80 ;
	7'h11 :
		RG_rl_68_t1 = TR_80 ;
	7'h12 :
		RG_rl_68_t1 = TR_80 ;
	7'h13 :
		RG_rl_68_t1 = TR_80 ;
	7'h14 :
		RG_rl_68_t1 = TR_80 ;
	7'h15 :
		RG_rl_68_t1 = TR_80 ;
	7'h16 :
		RG_rl_68_t1 = TR_80 ;
	7'h17 :
		RG_rl_68_t1 = TR_80 ;
	7'h18 :
		RG_rl_68_t1 = TR_80 ;
	7'h19 :
		RG_rl_68_t1 = TR_80 ;
	7'h1a :
		RG_rl_68_t1 = TR_80 ;
	7'h1b :
		RG_rl_68_t1 = TR_80 ;
	7'h1c :
		RG_rl_68_t1 = TR_80 ;
	7'h1d :
		RG_rl_68_t1 = TR_80 ;
	7'h1e :
		RG_rl_68_t1 = TR_80 ;
	7'h1f :
		RG_rl_68_t1 = TR_80 ;
	7'h20 :
		RG_rl_68_t1 = TR_80 ;
	7'h21 :
		RG_rl_68_t1 = TR_80 ;
	7'h22 :
		RG_rl_68_t1 = TR_80 ;
	7'h23 :
		RG_rl_68_t1 = TR_80 ;
	7'h24 :
		RG_rl_68_t1 = TR_80 ;
	7'h25 :
		RG_rl_68_t1 = TR_80 ;
	7'h26 :
		RG_rl_68_t1 = TR_80 ;
	7'h27 :
		RG_rl_68_t1 = TR_80 ;
	7'h28 :
		RG_rl_68_t1 = TR_80 ;
	7'h29 :
		RG_rl_68_t1 = TR_80 ;
	7'h2a :
		RG_rl_68_t1 = TR_80 ;
	7'h2b :
		RG_rl_68_t1 = TR_80 ;
	7'h2c :
		RG_rl_68_t1 = TR_80 ;
	7'h2d :
		RG_rl_68_t1 = TR_80 ;
	7'h2e :
		RG_rl_68_t1 = TR_80 ;
	7'h2f :
		RG_rl_68_t1 = TR_80 ;
	7'h30 :
		RG_rl_68_t1 = TR_80 ;
	7'h31 :
		RG_rl_68_t1 = TR_80 ;
	7'h32 :
		RG_rl_68_t1 = TR_80 ;
	7'h33 :
		RG_rl_68_t1 = TR_80 ;
	7'h34 :
		RG_rl_68_t1 = TR_80 ;
	7'h35 :
		RG_rl_68_t1 = TR_80 ;
	7'h36 :
		RG_rl_68_t1 = TR_80 ;
	7'h37 :
		RG_rl_68_t1 = TR_80 ;
	7'h38 :
		RG_rl_68_t1 = TR_80 ;
	7'h39 :
		RG_rl_68_t1 = TR_80 ;
	7'h3a :
		RG_rl_68_t1 = TR_80 ;
	7'h3b :
		RG_rl_68_t1 = TR_80 ;
	7'h3c :
		RG_rl_68_t1 = TR_80 ;
	7'h3d :
		RG_rl_68_t1 = TR_80 ;
	7'h3e :
		RG_rl_68_t1 = TR_80 ;
	7'h3f :
		RG_rl_68_t1 = TR_80 ;
	7'h40 :
		RG_rl_68_t1 = TR_80 ;
	7'h41 :
		RG_rl_68_t1 = TR_80 ;
	7'h42 :
		RG_rl_68_t1 = TR_80 ;
	7'h43 :
		RG_rl_68_t1 = TR_80 ;
	7'h44 :
		RG_rl_68_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h45 :
		RG_rl_68_t1 = TR_80 ;
	7'h46 :
		RG_rl_68_t1 = TR_80 ;
	7'h47 :
		RG_rl_68_t1 = TR_80 ;
	7'h48 :
		RG_rl_68_t1 = TR_80 ;
	7'h49 :
		RG_rl_68_t1 = TR_80 ;
	7'h4a :
		RG_rl_68_t1 = TR_80 ;
	7'h4b :
		RG_rl_68_t1 = TR_80 ;
	7'h4c :
		RG_rl_68_t1 = TR_80 ;
	7'h4d :
		RG_rl_68_t1 = TR_80 ;
	7'h4e :
		RG_rl_68_t1 = TR_80 ;
	7'h4f :
		RG_rl_68_t1 = TR_80 ;
	7'h50 :
		RG_rl_68_t1 = TR_80 ;
	7'h51 :
		RG_rl_68_t1 = TR_80 ;
	7'h52 :
		RG_rl_68_t1 = TR_80 ;
	7'h53 :
		RG_rl_68_t1 = TR_80 ;
	7'h54 :
		RG_rl_68_t1 = TR_80 ;
	7'h55 :
		RG_rl_68_t1 = TR_80 ;
	7'h56 :
		RG_rl_68_t1 = TR_80 ;
	7'h57 :
		RG_rl_68_t1 = TR_80 ;
	7'h58 :
		RG_rl_68_t1 = TR_80 ;
	7'h59 :
		RG_rl_68_t1 = TR_80 ;
	7'h5a :
		RG_rl_68_t1 = TR_80 ;
	7'h5b :
		RG_rl_68_t1 = TR_80 ;
	7'h5c :
		RG_rl_68_t1 = TR_80 ;
	7'h5d :
		RG_rl_68_t1 = TR_80 ;
	7'h5e :
		RG_rl_68_t1 = TR_80 ;
	7'h5f :
		RG_rl_68_t1 = TR_80 ;
	7'h60 :
		RG_rl_68_t1 = TR_80 ;
	7'h61 :
		RG_rl_68_t1 = TR_80 ;
	7'h62 :
		RG_rl_68_t1 = TR_80 ;
	7'h63 :
		RG_rl_68_t1 = TR_80 ;
	7'h64 :
		RG_rl_68_t1 = TR_80 ;
	7'h65 :
		RG_rl_68_t1 = TR_80 ;
	7'h66 :
		RG_rl_68_t1 = TR_80 ;
	7'h67 :
		RG_rl_68_t1 = TR_80 ;
	7'h68 :
		RG_rl_68_t1 = TR_80 ;
	7'h69 :
		RG_rl_68_t1 = TR_80 ;
	7'h6a :
		RG_rl_68_t1 = TR_80 ;
	7'h6b :
		RG_rl_68_t1 = TR_80 ;
	7'h6c :
		RG_rl_68_t1 = TR_80 ;
	7'h6d :
		RG_rl_68_t1 = TR_80 ;
	7'h6e :
		RG_rl_68_t1 = TR_80 ;
	7'h6f :
		RG_rl_68_t1 = TR_80 ;
	7'h70 :
		RG_rl_68_t1 = TR_80 ;
	7'h71 :
		RG_rl_68_t1 = TR_80 ;
	7'h72 :
		RG_rl_68_t1 = TR_80 ;
	7'h73 :
		RG_rl_68_t1 = TR_80 ;
	7'h74 :
		RG_rl_68_t1 = TR_80 ;
	7'h75 :
		RG_rl_68_t1 = TR_80 ;
	7'h76 :
		RG_rl_68_t1 = TR_80 ;
	7'h77 :
		RG_rl_68_t1 = TR_80 ;
	7'h78 :
		RG_rl_68_t1 = TR_80 ;
	7'h79 :
		RG_rl_68_t1 = TR_80 ;
	7'h7a :
		RG_rl_68_t1 = TR_80 ;
	7'h7b :
		RG_rl_68_t1 = TR_80 ;
	7'h7c :
		RG_rl_68_t1 = TR_80 ;
	7'h7d :
		RG_rl_68_t1 = TR_80 ;
	7'h7e :
		RG_rl_68_t1 = TR_80 ;
	7'h7f :
		RG_rl_68_t1 = TR_80 ;
	default :
		RG_rl_68_t1 = 9'hx ;
	endcase
always @ ( RG_rl_68_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_9 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_68_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h44 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_68_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_9 )
		| ( { 9{ U_569 } } & RG_rl_68_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_68_en = ( U_570 | RG_rl_68_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_68_en )
		RG_rl_68 <= RG_rl_68_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_81 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_69_t1 = TR_81 ;
	7'h01 :
		RG_rl_69_t1 = TR_81 ;
	7'h02 :
		RG_rl_69_t1 = TR_81 ;
	7'h03 :
		RG_rl_69_t1 = TR_81 ;
	7'h04 :
		RG_rl_69_t1 = TR_81 ;
	7'h05 :
		RG_rl_69_t1 = TR_81 ;
	7'h06 :
		RG_rl_69_t1 = TR_81 ;
	7'h07 :
		RG_rl_69_t1 = TR_81 ;
	7'h08 :
		RG_rl_69_t1 = TR_81 ;
	7'h09 :
		RG_rl_69_t1 = TR_81 ;
	7'h0a :
		RG_rl_69_t1 = TR_81 ;
	7'h0b :
		RG_rl_69_t1 = TR_81 ;
	7'h0c :
		RG_rl_69_t1 = TR_81 ;
	7'h0d :
		RG_rl_69_t1 = TR_81 ;
	7'h0e :
		RG_rl_69_t1 = TR_81 ;
	7'h0f :
		RG_rl_69_t1 = TR_81 ;
	7'h10 :
		RG_rl_69_t1 = TR_81 ;
	7'h11 :
		RG_rl_69_t1 = TR_81 ;
	7'h12 :
		RG_rl_69_t1 = TR_81 ;
	7'h13 :
		RG_rl_69_t1 = TR_81 ;
	7'h14 :
		RG_rl_69_t1 = TR_81 ;
	7'h15 :
		RG_rl_69_t1 = TR_81 ;
	7'h16 :
		RG_rl_69_t1 = TR_81 ;
	7'h17 :
		RG_rl_69_t1 = TR_81 ;
	7'h18 :
		RG_rl_69_t1 = TR_81 ;
	7'h19 :
		RG_rl_69_t1 = TR_81 ;
	7'h1a :
		RG_rl_69_t1 = TR_81 ;
	7'h1b :
		RG_rl_69_t1 = TR_81 ;
	7'h1c :
		RG_rl_69_t1 = TR_81 ;
	7'h1d :
		RG_rl_69_t1 = TR_81 ;
	7'h1e :
		RG_rl_69_t1 = TR_81 ;
	7'h1f :
		RG_rl_69_t1 = TR_81 ;
	7'h20 :
		RG_rl_69_t1 = TR_81 ;
	7'h21 :
		RG_rl_69_t1 = TR_81 ;
	7'h22 :
		RG_rl_69_t1 = TR_81 ;
	7'h23 :
		RG_rl_69_t1 = TR_81 ;
	7'h24 :
		RG_rl_69_t1 = TR_81 ;
	7'h25 :
		RG_rl_69_t1 = TR_81 ;
	7'h26 :
		RG_rl_69_t1 = TR_81 ;
	7'h27 :
		RG_rl_69_t1 = TR_81 ;
	7'h28 :
		RG_rl_69_t1 = TR_81 ;
	7'h29 :
		RG_rl_69_t1 = TR_81 ;
	7'h2a :
		RG_rl_69_t1 = TR_81 ;
	7'h2b :
		RG_rl_69_t1 = TR_81 ;
	7'h2c :
		RG_rl_69_t1 = TR_81 ;
	7'h2d :
		RG_rl_69_t1 = TR_81 ;
	7'h2e :
		RG_rl_69_t1 = TR_81 ;
	7'h2f :
		RG_rl_69_t1 = TR_81 ;
	7'h30 :
		RG_rl_69_t1 = TR_81 ;
	7'h31 :
		RG_rl_69_t1 = TR_81 ;
	7'h32 :
		RG_rl_69_t1 = TR_81 ;
	7'h33 :
		RG_rl_69_t1 = TR_81 ;
	7'h34 :
		RG_rl_69_t1 = TR_81 ;
	7'h35 :
		RG_rl_69_t1 = TR_81 ;
	7'h36 :
		RG_rl_69_t1 = TR_81 ;
	7'h37 :
		RG_rl_69_t1 = TR_81 ;
	7'h38 :
		RG_rl_69_t1 = TR_81 ;
	7'h39 :
		RG_rl_69_t1 = TR_81 ;
	7'h3a :
		RG_rl_69_t1 = TR_81 ;
	7'h3b :
		RG_rl_69_t1 = TR_81 ;
	7'h3c :
		RG_rl_69_t1 = TR_81 ;
	7'h3d :
		RG_rl_69_t1 = TR_81 ;
	7'h3e :
		RG_rl_69_t1 = TR_81 ;
	7'h3f :
		RG_rl_69_t1 = TR_81 ;
	7'h40 :
		RG_rl_69_t1 = TR_81 ;
	7'h41 :
		RG_rl_69_t1 = TR_81 ;
	7'h42 :
		RG_rl_69_t1 = TR_81 ;
	7'h43 :
		RG_rl_69_t1 = TR_81 ;
	7'h44 :
		RG_rl_69_t1 = TR_81 ;
	7'h45 :
		RG_rl_69_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h46 :
		RG_rl_69_t1 = TR_81 ;
	7'h47 :
		RG_rl_69_t1 = TR_81 ;
	7'h48 :
		RG_rl_69_t1 = TR_81 ;
	7'h49 :
		RG_rl_69_t1 = TR_81 ;
	7'h4a :
		RG_rl_69_t1 = TR_81 ;
	7'h4b :
		RG_rl_69_t1 = TR_81 ;
	7'h4c :
		RG_rl_69_t1 = TR_81 ;
	7'h4d :
		RG_rl_69_t1 = TR_81 ;
	7'h4e :
		RG_rl_69_t1 = TR_81 ;
	7'h4f :
		RG_rl_69_t1 = TR_81 ;
	7'h50 :
		RG_rl_69_t1 = TR_81 ;
	7'h51 :
		RG_rl_69_t1 = TR_81 ;
	7'h52 :
		RG_rl_69_t1 = TR_81 ;
	7'h53 :
		RG_rl_69_t1 = TR_81 ;
	7'h54 :
		RG_rl_69_t1 = TR_81 ;
	7'h55 :
		RG_rl_69_t1 = TR_81 ;
	7'h56 :
		RG_rl_69_t1 = TR_81 ;
	7'h57 :
		RG_rl_69_t1 = TR_81 ;
	7'h58 :
		RG_rl_69_t1 = TR_81 ;
	7'h59 :
		RG_rl_69_t1 = TR_81 ;
	7'h5a :
		RG_rl_69_t1 = TR_81 ;
	7'h5b :
		RG_rl_69_t1 = TR_81 ;
	7'h5c :
		RG_rl_69_t1 = TR_81 ;
	7'h5d :
		RG_rl_69_t1 = TR_81 ;
	7'h5e :
		RG_rl_69_t1 = TR_81 ;
	7'h5f :
		RG_rl_69_t1 = TR_81 ;
	7'h60 :
		RG_rl_69_t1 = TR_81 ;
	7'h61 :
		RG_rl_69_t1 = TR_81 ;
	7'h62 :
		RG_rl_69_t1 = TR_81 ;
	7'h63 :
		RG_rl_69_t1 = TR_81 ;
	7'h64 :
		RG_rl_69_t1 = TR_81 ;
	7'h65 :
		RG_rl_69_t1 = TR_81 ;
	7'h66 :
		RG_rl_69_t1 = TR_81 ;
	7'h67 :
		RG_rl_69_t1 = TR_81 ;
	7'h68 :
		RG_rl_69_t1 = TR_81 ;
	7'h69 :
		RG_rl_69_t1 = TR_81 ;
	7'h6a :
		RG_rl_69_t1 = TR_81 ;
	7'h6b :
		RG_rl_69_t1 = TR_81 ;
	7'h6c :
		RG_rl_69_t1 = TR_81 ;
	7'h6d :
		RG_rl_69_t1 = TR_81 ;
	7'h6e :
		RG_rl_69_t1 = TR_81 ;
	7'h6f :
		RG_rl_69_t1 = TR_81 ;
	7'h70 :
		RG_rl_69_t1 = TR_81 ;
	7'h71 :
		RG_rl_69_t1 = TR_81 ;
	7'h72 :
		RG_rl_69_t1 = TR_81 ;
	7'h73 :
		RG_rl_69_t1 = TR_81 ;
	7'h74 :
		RG_rl_69_t1 = TR_81 ;
	7'h75 :
		RG_rl_69_t1 = TR_81 ;
	7'h76 :
		RG_rl_69_t1 = TR_81 ;
	7'h77 :
		RG_rl_69_t1 = TR_81 ;
	7'h78 :
		RG_rl_69_t1 = TR_81 ;
	7'h79 :
		RG_rl_69_t1 = TR_81 ;
	7'h7a :
		RG_rl_69_t1 = TR_81 ;
	7'h7b :
		RG_rl_69_t1 = TR_81 ;
	7'h7c :
		RG_rl_69_t1 = TR_81 ;
	7'h7d :
		RG_rl_69_t1 = TR_81 ;
	7'h7e :
		RG_rl_69_t1 = TR_81 ;
	7'h7f :
		RG_rl_69_t1 = TR_81 ;
	default :
		RG_rl_69_t1 = 9'hx ;
	endcase
always @ ( RG_rl_69_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_10 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_69_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h45 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_69_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_10 )
		| ( { 9{ U_569 } } & RG_rl_69_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_69_en = ( U_570 | RG_rl_69_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_69_en )
		RG_rl_69 <= RG_rl_69_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_82 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_70_t1 = TR_82 ;
	7'h01 :
		RG_rl_70_t1 = TR_82 ;
	7'h02 :
		RG_rl_70_t1 = TR_82 ;
	7'h03 :
		RG_rl_70_t1 = TR_82 ;
	7'h04 :
		RG_rl_70_t1 = TR_82 ;
	7'h05 :
		RG_rl_70_t1 = TR_82 ;
	7'h06 :
		RG_rl_70_t1 = TR_82 ;
	7'h07 :
		RG_rl_70_t1 = TR_82 ;
	7'h08 :
		RG_rl_70_t1 = TR_82 ;
	7'h09 :
		RG_rl_70_t1 = TR_82 ;
	7'h0a :
		RG_rl_70_t1 = TR_82 ;
	7'h0b :
		RG_rl_70_t1 = TR_82 ;
	7'h0c :
		RG_rl_70_t1 = TR_82 ;
	7'h0d :
		RG_rl_70_t1 = TR_82 ;
	7'h0e :
		RG_rl_70_t1 = TR_82 ;
	7'h0f :
		RG_rl_70_t1 = TR_82 ;
	7'h10 :
		RG_rl_70_t1 = TR_82 ;
	7'h11 :
		RG_rl_70_t1 = TR_82 ;
	7'h12 :
		RG_rl_70_t1 = TR_82 ;
	7'h13 :
		RG_rl_70_t1 = TR_82 ;
	7'h14 :
		RG_rl_70_t1 = TR_82 ;
	7'h15 :
		RG_rl_70_t1 = TR_82 ;
	7'h16 :
		RG_rl_70_t1 = TR_82 ;
	7'h17 :
		RG_rl_70_t1 = TR_82 ;
	7'h18 :
		RG_rl_70_t1 = TR_82 ;
	7'h19 :
		RG_rl_70_t1 = TR_82 ;
	7'h1a :
		RG_rl_70_t1 = TR_82 ;
	7'h1b :
		RG_rl_70_t1 = TR_82 ;
	7'h1c :
		RG_rl_70_t1 = TR_82 ;
	7'h1d :
		RG_rl_70_t1 = TR_82 ;
	7'h1e :
		RG_rl_70_t1 = TR_82 ;
	7'h1f :
		RG_rl_70_t1 = TR_82 ;
	7'h20 :
		RG_rl_70_t1 = TR_82 ;
	7'h21 :
		RG_rl_70_t1 = TR_82 ;
	7'h22 :
		RG_rl_70_t1 = TR_82 ;
	7'h23 :
		RG_rl_70_t1 = TR_82 ;
	7'h24 :
		RG_rl_70_t1 = TR_82 ;
	7'h25 :
		RG_rl_70_t1 = TR_82 ;
	7'h26 :
		RG_rl_70_t1 = TR_82 ;
	7'h27 :
		RG_rl_70_t1 = TR_82 ;
	7'h28 :
		RG_rl_70_t1 = TR_82 ;
	7'h29 :
		RG_rl_70_t1 = TR_82 ;
	7'h2a :
		RG_rl_70_t1 = TR_82 ;
	7'h2b :
		RG_rl_70_t1 = TR_82 ;
	7'h2c :
		RG_rl_70_t1 = TR_82 ;
	7'h2d :
		RG_rl_70_t1 = TR_82 ;
	7'h2e :
		RG_rl_70_t1 = TR_82 ;
	7'h2f :
		RG_rl_70_t1 = TR_82 ;
	7'h30 :
		RG_rl_70_t1 = TR_82 ;
	7'h31 :
		RG_rl_70_t1 = TR_82 ;
	7'h32 :
		RG_rl_70_t1 = TR_82 ;
	7'h33 :
		RG_rl_70_t1 = TR_82 ;
	7'h34 :
		RG_rl_70_t1 = TR_82 ;
	7'h35 :
		RG_rl_70_t1 = TR_82 ;
	7'h36 :
		RG_rl_70_t1 = TR_82 ;
	7'h37 :
		RG_rl_70_t1 = TR_82 ;
	7'h38 :
		RG_rl_70_t1 = TR_82 ;
	7'h39 :
		RG_rl_70_t1 = TR_82 ;
	7'h3a :
		RG_rl_70_t1 = TR_82 ;
	7'h3b :
		RG_rl_70_t1 = TR_82 ;
	7'h3c :
		RG_rl_70_t1 = TR_82 ;
	7'h3d :
		RG_rl_70_t1 = TR_82 ;
	7'h3e :
		RG_rl_70_t1 = TR_82 ;
	7'h3f :
		RG_rl_70_t1 = TR_82 ;
	7'h40 :
		RG_rl_70_t1 = TR_82 ;
	7'h41 :
		RG_rl_70_t1 = TR_82 ;
	7'h42 :
		RG_rl_70_t1 = TR_82 ;
	7'h43 :
		RG_rl_70_t1 = TR_82 ;
	7'h44 :
		RG_rl_70_t1 = TR_82 ;
	7'h45 :
		RG_rl_70_t1 = TR_82 ;
	7'h46 :
		RG_rl_70_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h47 :
		RG_rl_70_t1 = TR_82 ;
	7'h48 :
		RG_rl_70_t1 = TR_82 ;
	7'h49 :
		RG_rl_70_t1 = TR_82 ;
	7'h4a :
		RG_rl_70_t1 = TR_82 ;
	7'h4b :
		RG_rl_70_t1 = TR_82 ;
	7'h4c :
		RG_rl_70_t1 = TR_82 ;
	7'h4d :
		RG_rl_70_t1 = TR_82 ;
	7'h4e :
		RG_rl_70_t1 = TR_82 ;
	7'h4f :
		RG_rl_70_t1 = TR_82 ;
	7'h50 :
		RG_rl_70_t1 = TR_82 ;
	7'h51 :
		RG_rl_70_t1 = TR_82 ;
	7'h52 :
		RG_rl_70_t1 = TR_82 ;
	7'h53 :
		RG_rl_70_t1 = TR_82 ;
	7'h54 :
		RG_rl_70_t1 = TR_82 ;
	7'h55 :
		RG_rl_70_t1 = TR_82 ;
	7'h56 :
		RG_rl_70_t1 = TR_82 ;
	7'h57 :
		RG_rl_70_t1 = TR_82 ;
	7'h58 :
		RG_rl_70_t1 = TR_82 ;
	7'h59 :
		RG_rl_70_t1 = TR_82 ;
	7'h5a :
		RG_rl_70_t1 = TR_82 ;
	7'h5b :
		RG_rl_70_t1 = TR_82 ;
	7'h5c :
		RG_rl_70_t1 = TR_82 ;
	7'h5d :
		RG_rl_70_t1 = TR_82 ;
	7'h5e :
		RG_rl_70_t1 = TR_82 ;
	7'h5f :
		RG_rl_70_t1 = TR_82 ;
	7'h60 :
		RG_rl_70_t1 = TR_82 ;
	7'h61 :
		RG_rl_70_t1 = TR_82 ;
	7'h62 :
		RG_rl_70_t1 = TR_82 ;
	7'h63 :
		RG_rl_70_t1 = TR_82 ;
	7'h64 :
		RG_rl_70_t1 = TR_82 ;
	7'h65 :
		RG_rl_70_t1 = TR_82 ;
	7'h66 :
		RG_rl_70_t1 = TR_82 ;
	7'h67 :
		RG_rl_70_t1 = TR_82 ;
	7'h68 :
		RG_rl_70_t1 = TR_82 ;
	7'h69 :
		RG_rl_70_t1 = TR_82 ;
	7'h6a :
		RG_rl_70_t1 = TR_82 ;
	7'h6b :
		RG_rl_70_t1 = TR_82 ;
	7'h6c :
		RG_rl_70_t1 = TR_82 ;
	7'h6d :
		RG_rl_70_t1 = TR_82 ;
	7'h6e :
		RG_rl_70_t1 = TR_82 ;
	7'h6f :
		RG_rl_70_t1 = TR_82 ;
	7'h70 :
		RG_rl_70_t1 = TR_82 ;
	7'h71 :
		RG_rl_70_t1 = TR_82 ;
	7'h72 :
		RG_rl_70_t1 = TR_82 ;
	7'h73 :
		RG_rl_70_t1 = TR_82 ;
	7'h74 :
		RG_rl_70_t1 = TR_82 ;
	7'h75 :
		RG_rl_70_t1 = TR_82 ;
	7'h76 :
		RG_rl_70_t1 = TR_82 ;
	7'h77 :
		RG_rl_70_t1 = TR_82 ;
	7'h78 :
		RG_rl_70_t1 = TR_82 ;
	7'h79 :
		RG_rl_70_t1 = TR_82 ;
	7'h7a :
		RG_rl_70_t1 = TR_82 ;
	7'h7b :
		RG_rl_70_t1 = TR_82 ;
	7'h7c :
		RG_rl_70_t1 = TR_82 ;
	7'h7d :
		RG_rl_70_t1 = TR_82 ;
	7'h7e :
		RG_rl_70_t1 = TR_82 ;
	7'h7f :
		RG_rl_70_t1 = TR_82 ;
	default :
		RG_rl_70_t1 = 9'hx ;
	endcase
always @ ( RG_rl_70_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_11 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_70_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h46 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_70_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_11 )
		| ( { 9{ U_569 } } & RG_rl_70_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_70_en = ( U_570 | RG_rl_70_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_70_en )
		RG_rl_70 <= RG_rl_70_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_83 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_71_t1 = TR_83 ;
	7'h01 :
		RG_rl_71_t1 = TR_83 ;
	7'h02 :
		RG_rl_71_t1 = TR_83 ;
	7'h03 :
		RG_rl_71_t1 = TR_83 ;
	7'h04 :
		RG_rl_71_t1 = TR_83 ;
	7'h05 :
		RG_rl_71_t1 = TR_83 ;
	7'h06 :
		RG_rl_71_t1 = TR_83 ;
	7'h07 :
		RG_rl_71_t1 = TR_83 ;
	7'h08 :
		RG_rl_71_t1 = TR_83 ;
	7'h09 :
		RG_rl_71_t1 = TR_83 ;
	7'h0a :
		RG_rl_71_t1 = TR_83 ;
	7'h0b :
		RG_rl_71_t1 = TR_83 ;
	7'h0c :
		RG_rl_71_t1 = TR_83 ;
	7'h0d :
		RG_rl_71_t1 = TR_83 ;
	7'h0e :
		RG_rl_71_t1 = TR_83 ;
	7'h0f :
		RG_rl_71_t1 = TR_83 ;
	7'h10 :
		RG_rl_71_t1 = TR_83 ;
	7'h11 :
		RG_rl_71_t1 = TR_83 ;
	7'h12 :
		RG_rl_71_t1 = TR_83 ;
	7'h13 :
		RG_rl_71_t1 = TR_83 ;
	7'h14 :
		RG_rl_71_t1 = TR_83 ;
	7'h15 :
		RG_rl_71_t1 = TR_83 ;
	7'h16 :
		RG_rl_71_t1 = TR_83 ;
	7'h17 :
		RG_rl_71_t1 = TR_83 ;
	7'h18 :
		RG_rl_71_t1 = TR_83 ;
	7'h19 :
		RG_rl_71_t1 = TR_83 ;
	7'h1a :
		RG_rl_71_t1 = TR_83 ;
	7'h1b :
		RG_rl_71_t1 = TR_83 ;
	7'h1c :
		RG_rl_71_t1 = TR_83 ;
	7'h1d :
		RG_rl_71_t1 = TR_83 ;
	7'h1e :
		RG_rl_71_t1 = TR_83 ;
	7'h1f :
		RG_rl_71_t1 = TR_83 ;
	7'h20 :
		RG_rl_71_t1 = TR_83 ;
	7'h21 :
		RG_rl_71_t1 = TR_83 ;
	7'h22 :
		RG_rl_71_t1 = TR_83 ;
	7'h23 :
		RG_rl_71_t1 = TR_83 ;
	7'h24 :
		RG_rl_71_t1 = TR_83 ;
	7'h25 :
		RG_rl_71_t1 = TR_83 ;
	7'h26 :
		RG_rl_71_t1 = TR_83 ;
	7'h27 :
		RG_rl_71_t1 = TR_83 ;
	7'h28 :
		RG_rl_71_t1 = TR_83 ;
	7'h29 :
		RG_rl_71_t1 = TR_83 ;
	7'h2a :
		RG_rl_71_t1 = TR_83 ;
	7'h2b :
		RG_rl_71_t1 = TR_83 ;
	7'h2c :
		RG_rl_71_t1 = TR_83 ;
	7'h2d :
		RG_rl_71_t1 = TR_83 ;
	7'h2e :
		RG_rl_71_t1 = TR_83 ;
	7'h2f :
		RG_rl_71_t1 = TR_83 ;
	7'h30 :
		RG_rl_71_t1 = TR_83 ;
	7'h31 :
		RG_rl_71_t1 = TR_83 ;
	7'h32 :
		RG_rl_71_t1 = TR_83 ;
	7'h33 :
		RG_rl_71_t1 = TR_83 ;
	7'h34 :
		RG_rl_71_t1 = TR_83 ;
	7'h35 :
		RG_rl_71_t1 = TR_83 ;
	7'h36 :
		RG_rl_71_t1 = TR_83 ;
	7'h37 :
		RG_rl_71_t1 = TR_83 ;
	7'h38 :
		RG_rl_71_t1 = TR_83 ;
	7'h39 :
		RG_rl_71_t1 = TR_83 ;
	7'h3a :
		RG_rl_71_t1 = TR_83 ;
	7'h3b :
		RG_rl_71_t1 = TR_83 ;
	7'h3c :
		RG_rl_71_t1 = TR_83 ;
	7'h3d :
		RG_rl_71_t1 = TR_83 ;
	7'h3e :
		RG_rl_71_t1 = TR_83 ;
	7'h3f :
		RG_rl_71_t1 = TR_83 ;
	7'h40 :
		RG_rl_71_t1 = TR_83 ;
	7'h41 :
		RG_rl_71_t1 = TR_83 ;
	7'h42 :
		RG_rl_71_t1 = TR_83 ;
	7'h43 :
		RG_rl_71_t1 = TR_83 ;
	7'h44 :
		RG_rl_71_t1 = TR_83 ;
	7'h45 :
		RG_rl_71_t1 = TR_83 ;
	7'h46 :
		RG_rl_71_t1 = TR_83 ;
	7'h47 :
		RG_rl_71_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h48 :
		RG_rl_71_t1 = TR_83 ;
	7'h49 :
		RG_rl_71_t1 = TR_83 ;
	7'h4a :
		RG_rl_71_t1 = TR_83 ;
	7'h4b :
		RG_rl_71_t1 = TR_83 ;
	7'h4c :
		RG_rl_71_t1 = TR_83 ;
	7'h4d :
		RG_rl_71_t1 = TR_83 ;
	7'h4e :
		RG_rl_71_t1 = TR_83 ;
	7'h4f :
		RG_rl_71_t1 = TR_83 ;
	7'h50 :
		RG_rl_71_t1 = TR_83 ;
	7'h51 :
		RG_rl_71_t1 = TR_83 ;
	7'h52 :
		RG_rl_71_t1 = TR_83 ;
	7'h53 :
		RG_rl_71_t1 = TR_83 ;
	7'h54 :
		RG_rl_71_t1 = TR_83 ;
	7'h55 :
		RG_rl_71_t1 = TR_83 ;
	7'h56 :
		RG_rl_71_t1 = TR_83 ;
	7'h57 :
		RG_rl_71_t1 = TR_83 ;
	7'h58 :
		RG_rl_71_t1 = TR_83 ;
	7'h59 :
		RG_rl_71_t1 = TR_83 ;
	7'h5a :
		RG_rl_71_t1 = TR_83 ;
	7'h5b :
		RG_rl_71_t1 = TR_83 ;
	7'h5c :
		RG_rl_71_t1 = TR_83 ;
	7'h5d :
		RG_rl_71_t1 = TR_83 ;
	7'h5e :
		RG_rl_71_t1 = TR_83 ;
	7'h5f :
		RG_rl_71_t1 = TR_83 ;
	7'h60 :
		RG_rl_71_t1 = TR_83 ;
	7'h61 :
		RG_rl_71_t1 = TR_83 ;
	7'h62 :
		RG_rl_71_t1 = TR_83 ;
	7'h63 :
		RG_rl_71_t1 = TR_83 ;
	7'h64 :
		RG_rl_71_t1 = TR_83 ;
	7'h65 :
		RG_rl_71_t1 = TR_83 ;
	7'h66 :
		RG_rl_71_t1 = TR_83 ;
	7'h67 :
		RG_rl_71_t1 = TR_83 ;
	7'h68 :
		RG_rl_71_t1 = TR_83 ;
	7'h69 :
		RG_rl_71_t1 = TR_83 ;
	7'h6a :
		RG_rl_71_t1 = TR_83 ;
	7'h6b :
		RG_rl_71_t1 = TR_83 ;
	7'h6c :
		RG_rl_71_t1 = TR_83 ;
	7'h6d :
		RG_rl_71_t1 = TR_83 ;
	7'h6e :
		RG_rl_71_t1 = TR_83 ;
	7'h6f :
		RG_rl_71_t1 = TR_83 ;
	7'h70 :
		RG_rl_71_t1 = TR_83 ;
	7'h71 :
		RG_rl_71_t1 = TR_83 ;
	7'h72 :
		RG_rl_71_t1 = TR_83 ;
	7'h73 :
		RG_rl_71_t1 = TR_83 ;
	7'h74 :
		RG_rl_71_t1 = TR_83 ;
	7'h75 :
		RG_rl_71_t1 = TR_83 ;
	7'h76 :
		RG_rl_71_t1 = TR_83 ;
	7'h77 :
		RG_rl_71_t1 = TR_83 ;
	7'h78 :
		RG_rl_71_t1 = TR_83 ;
	7'h79 :
		RG_rl_71_t1 = TR_83 ;
	7'h7a :
		RG_rl_71_t1 = TR_83 ;
	7'h7b :
		RG_rl_71_t1 = TR_83 ;
	7'h7c :
		RG_rl_71_t1 = TR_83 ;
	7'h7d :
		RG_rl_71_t1 = TR_83 ;
	7'h7e :
		RG_rl_71_t1 = TR_83 ;
	7'h7f :
		RG_rl_71_t1 = TR_83 ;
	default :
		RG_rl_71_t1 = 9'hx ;
	endcase
always @ ( RG_rl_71_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_12 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_71_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h47 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_71_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_12 )
		| ( { 9{ U_569 } } & RG_rl_71_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_71_en = ( U_570 | RG_rl_71_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_71_en )
		RG_rl_71 <= RG_rl_71_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_84 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_72_t1 = TR_84 ;
	7'h01 :
		RG_rl_72_t1 = TR_84 ;
	7'h02 :
		RG_rl_72_t1 = TR_84 ;
	7'h03 :
		RG_rl_72_t1 = TR_84 ;
	7'h04 :
		RG_rl_72_t1 = TR_84 ;
	7'h05 :
		RG_rl_72_t1 = TR_84 ;
	7'h06 :
		RG_rl_72_t1 = TR_84 ;
	7'h07 :
		RG_rl_72_t1 = TR_84 ;
	7'h08 :
		RG_rl_72_t1 = TR_84 ;
	7'h09 :
		RG_rl_72_t1 = TR_84 ;
	7'h0a :
		RG_rl_72_t1 = TR_84 ;
	7'h0b :
		RG_rl_72_t1 = TR_84 ;
	7'h0c :
		RG_rl_72_t1 = TR_84 ;
	7'h0d :
		RG_rl_72_t1 = TR_84 ;
	7'h0e :
		RG_rl_72_t1 = TR_84 ;
	7'h0f :
		RG_rl_72_t1 = TR_84 ;
	7'h10 :
		RG_rl_72_t1 = TR_84 ;
	7'h11 :
		RG_rl_72_t1 = TR_84 ;
	7'h12 :
		RG_rl_72_t1 = TR_84 ;
	7'h13 :
		RG_rl_72_t1 = TR_84 ;
	7'h14 :
		RG_rl_72_t1 = TR_84 ;
	7'h15 :
		RG_rl_72_t1 = TR_84 ;
	7'h16 :
		RG_rl_72_t1 = TR_84 ;
	7'h17 :
		RG_rl_72_t1 = TR_84 ;
	7'h18 :
		RG_rl_72_t1 = TR_84 ;
	7'h19 :
		RG_rl_72_t1 = TR_84 ;
	7'h1a :
		RG_rl_72_t1 = TR_84 ;
	7'h1b :
		RG_rl_72_t1 = TR_84 ;
	7'h1c :
		RG_rl_72_t1 = TR_84 ;
	7'h1d :
		RG_rl_72_t1 = TR_84 ;
	7'h1e :
		RG_rl_72_t1 = TR_84 ;
	7'h1f :
		RG_rl_72_t1 = TR_84 ;
	7'h20 :
		RG_rl_72_t1 = TR_84 ;
	7'h21 :
		RG_rl_72_t1 = TR_84 ;
	7'h22 :
		RG_rl_72_t1 = TR_84 ;
	7'h23 :
		RG_rl_72_t1 = TR_84 ;
	7'h24 :
		RG_rl_72_t1 = TR_84 ;
	7'h25 :
		RG_rl_72_t1 = TR_84 ;
	7'h26 :
		RG_rl_72_t1 = TR_84 ;
	7'h27 :
		RG_rl_72_t1 = TR_84 ;
	7'h28 :
		RG_rl_72_t1 = TR_84 ;
	7'h29 :
		RG_rl_72_t1 = TR_84 ;
	7'h2a :
		RG_rl_72_t1 = TR_84 ;
	7'h2b :
		RG_rl_72_t1 = TR_84 ;
	7'h2c :
		RG_rl_72_t1 = TR_84 ;
	7'h2d :
		RG_rl_72_t1 = TR_84 ;
	7'h2e :
		RG_rl_72_t1 = TR_84 ;
	7'h2f :
		RG_rl_72_t1 = TR_84 ;
	7'h30 :
		RG_rl_72_t1 = TR_84 ;
	7'h31 :
		RG_rl_72_t1 = TR_84 ;
	7'h32 :
		RG_rl_72_t1 = TR_84 ;
	7'h33 :
		RG_rl_72_t1 = TR_84 ;
	7'h34 :
		RG_rl_72_t1 = TR_84 ;
	7'h35 :
		RG_rl_72_t1 = TR_84 ;
	7'h36 :
		RG_rl_72_t1 = TR_84 ;
	7'h37 :
		RG_rl_72_t1 = TR_84 ;
	7'h38 :
		RG_rl_72_t1 = TR_84 ;
	7'h39 :
		RG_rl_72_t1 = TR_84 ;
	7'h3a :
		RG_rl_72_t1 = TR_84 ;
	7'h3b :
		RG_rl_72_t1 = TR_84 ;
	7'h3c :
		RG_rl_72_t1 = TR_84 ;
	7'h3d :
		RG_rl_72_t1 = TR_84 ;
	7'h3e :
		RG_rl_72_t1 = TR_84 ;
	7'h3f :
		RG_rl_72_t1 = TR_84 ;
	7'h40 :
		RG_rl_72_t1 = TR_84 ;
	7'h41 :
		RG_rl_72_t1 = TR_84 ;
	7'h42 :
		RG_rl_72_t1 = TR_84 ;
	7'h43 :
		RG_rl_72_t1 = TR_84 ;
	7'h44 :
		RG_rl_72_t1 = TR_84 ;
	7'h45 :
		RG_rl_72_t1 = TR_84 ;
	7'h46 :
		RG_rl_72_t1 = TR_84 ;
	7'h47 :
		RG_rl_72_t1 = TR_84 ;
	7'h48 :
		RG_rl_72_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h49 :
		RG_rl_72_t1 = TR_84 ;
	7'h4a :
		RG_rl_72_t1 = TR_84 ;
	7'h4b :
		RG_rl_72_t1 = TR_84 ;
	7'h4c :
		RG_rl_72_t1 = TR_84 ;
	7'h4d :
		RG_rl_72_t1 = TR_84 ;
	7'h4e :
		RG_rl_72_t1 = TR_84 ;
	7'h4f :
		RG_rl_72_t1 = TR_84 ;
	7'h50 :
		RG_rl_72_t1 = TR_84 ;
	7'h51 :
		RG_rl_72_t1 = TR_84 ;
	7'h52 :
		RG_rl_72_t1 = TR_84 ;
	7'h53 :
		RG_rl_72_t1 = TR_84 ;
	7'h54 :
		RG_rl_72_t1 = TR_84 ;
	7'h55 :
		RG_rl_72_t1 = TR_84 ;
	7'h56 :
		RG_rl_72_t1 = TR_84 ;
	7'h57 :
		RG_rl_72_t1 = TR_84 ;
	7'h58 :
		RG_rl_72_t1 = TR_84 ;
	7'h59 :
		RG_rl_72_t1 = TR_84 ;
	7'h5a :
		RG_rl_72_t1 = TR_84 ;
	7'h5b :
		RG_rl_72_t1 = TR_84 ;
	7'h5c :
		RG_rl_72_t1 = TR_84 ;
	7'h5d :
		RG_rl_72_t1 = TR_84 ;
	7'h5e :
		RG_rl_72_t1 = TR_84 ;
	7'h5f :
		RG_rl_72_t1 = TR_84 ;
	7'h60 :
		RG_rl_72_t1 = TR_84 ;
	7'h61 :
		RG_rl_72_t1 = TR_84 ;
	7'h62 :
		RG_rl_72_t1 = TR_84 ;
	7'h63 :
		RG_rl_72_t1 = TR_84 ;
	7'h64 :
		RG_rl_72_t1 = TR_84 ;
	7'h65 :
		RG_rl_72_t1 = TR_84 ;
	7'h66 :
		RG_rl_72_t1 = TR_84 ;
	7'h67 :
		RG_rl_72_t1 = TR_84 ;
	7'h68 :
		RG_rl_72_t1 = TR_84 ;
	7'h69 :
		RG_rl_72_t1 = TR_84 ;
	7'h6a :
		RG_rl_72_t1 = TR_84 ;
	7'h6b :
		RG_rl_72_t1 = TR_84 ;
	7'h6c :
		RG_rl_72_t1 = TR_84 ;
	7'h6d :
		RG_rl_72_t1 = TR_84 ;
	7'h6e :
		RG_rl_72_t1 = TR_84 ;
	7'h6f :
		RG_rl_72_t1 = TR_84 ;
	7'h70 :
		RG_rl_72_t1 = TR_84 ;
	7'h71 :
		RG_rl_72_t1 = TR_84 ;
	7'h72 :
		RG_rl_72_t1 = TR_84 ;
	7'h73 :
		RG_rl_72_t1 = TR_84 ;
	7'h74 :
		RG_rl_72_t1 = TR_84 ;
	7'h75 :
		RG_rl_72_t1 = TR_84 ;
	7'h76 :
		RG_rl_72_t1 = TR_84 ;
	7'h77 :
		RG_rl_72_t1 = TR_84 ;
	7'h78 :
		RG_rl_72_t1 = TR_84 ;
	7'h79 :
		RG_rl_72_t1 = TR_84 ;
	7'h7a :
		RG_rl_72_t1 = TR_84 ;
	7'h7b :
		RG_rl_72_t1 = TR_84 ;
	7'h7c :
		RG_rl_72_t1 = TR_84 ;
	7'h7d :
		RG_rl_72_t1 = TR_84 ;
	7'h7e :
		RG_rl_72_t1 = TR_84 ;
	7'h7f :
		RG_rl_72_t1 = TR_84 ;
	default :
		RG_rl_72_t1 = 9'hx ;
	endcase
always @ ( RG_rl_72_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_13 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_72_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h48 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_72_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_13 )
		| ( { 9{ U_569 } } & RG_rl_72_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_72_en = ( U_570 | RG_rl_72_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_72_en )
		RG_rl_72 <= RG_rl_72_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_85 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_73_t1 = TR_85 ;
	7'h01 :
		RG_rl_73_t1 = TR_85 ;
	7'h02 :
		RG_rl_73_t1 = TR_85 ;
	7'h03 :
		RG_rl_73_t1 = TR_85 ;
	7'h04 :
		RG_rl_73_t1 = TR_85 ;
	7'h05 :
		RG_rl_73_t1 = TR_85 ;
	7'h06 :
		RG_rl_73_t1 = TR_85 ;
	7'h07 :
		RG_rl_73_t1 = TR_85 ;
	7'h08 :
		RG_rl_73_t1 = TR_85 ;
	7'h09 :
		RG_rl_73_t1 = TR_85 ;
	7'h0a :
		RG_rl_73_t1 = TR_85 ;
	7'h0b :
		RG_rl_73_t1 = TR_85 ;
	7'h0c :
		RG_rl_73_t1 = TR_85 ;
	7'h0d :
		RG_rl_73_t1 = TR_85 ;
	7'h0e :
		RG_rl_73_t1 = TR_85 ;
	7'h0f :
		RG_rl_73_t1 = TR_85 ;
	7'h10 :
		RG_rl_73_t1 = TR_85 ;
	7'h11 :
		RG_rl_73_t1 = TR_85 ;
	7'h12 :
		RG_rl_73_t1 = TR_85 ;
	7'h13 :
		RG_rl_73_t1 = TR_85 ;
	7'h14 :
		RG_rl_73_t1 = TR_85 ;
	7'h15 :
		RG_rl_73_t1 = TR_85 ;
	7'h16 :
		RG_rl_73_t1 = TR_85 ;
	7'h17 :
		RG_rl_73_t1 = TR_85 ;
	7'h18 :
		RG_rl_73_t1 = TR_85 ;
	7'h19 :
		RG_rl_73_t1 = TR_85 ;
	7'h1a :
		RG_rl_73_t1 = TR_85 ;
	7'h1b :
		RG_rl_73_t1 = TR_85 ;
	7'h1c :
		RG_rl_73_t1 = TR_85 ;
	7'h1d :
		RG_rl_73_t1 = TR_85 ;
	7'h1e :
		RG_rl_73_t1 = TR_85 ;
	7'h1f :
		RG_rl_73_t1 = TR_85 ;
	7'h20 :
		RG_rl_73_t1 = TR_85 ;
	7'h21 :
		RG_rl_73_t1 = TR_85 ;
	7'h22 :
		RG_rl_73_t1 = TR_85 ;
	7'h23 :
		RG_rl_73_t1 = TR_85 ;
	7'h24 :
		RG_rl_73_t1 = TR_85 ;
	7'h25 :
		RG_rl_73_t1 = TR_85 ;
	7'h26 :
		RG_rl_73_t1 = TR_85 ;
	7'h27 :
		RG_rl_73_t1 = TR_85 ;
	7'h28 :
		RG_rl_73_t1 = TR_85 ;
	7'h29 :
		RG_rl_73_t1 = TR_85 ;
	7'h2a :
		RG_rl_73_t1 = TR_85 ;
	7'h2b :
		RG_rl_73_t1 = TR_85 ;
	7'h2c :
		RG_rl_73_t1 = TR_85 ;
	7'h2d :
		RG_rl_73_t1 = TR_85 ;
	7'h2e :
		RG_rl_73_t1 = TR_85 ;
	7'h2f :
		RG_rl_73_t1 = TR_85 ;
	7'h30 :
		RG_rl_73_t1 = TR_85 ;
	7'h31 :
		RG_rl_73_t1 = TR_85 ;
	7'h32 :
		RG_rl_73_t1 = TR_85 ;
	7'h33 :
		RG_rl_73_t1 = TR_85 ;
	7'h34 :
		RG_rl_73_t1 = TR_85 ;
	7'h35 :
		RG_rl_73_t1 = TR_85 ;
	7'h36 :
		RG_rl_73_t1 = TR_85 ;
	7'h37 :
		RG_rl_73_t1 = TR_85 ;
	7'h38 :
		RG_rl_73_t1 = TR_85 ;
	7'h39 :
		RG_rl_73_t1 = TR_85 ;
	7'h3a :
		RG_rl_73_t1 = TR_85 ;
	7'h3b :
		RG_rl_73_t1 = TR_85 ;
	7'h3c :
		RG_rl_73_t1 = TR_85 ;
	7'h3d :
		RG_rl_73_t1 = TR_85 ;
	7'h3e :
		RG_rl_73_t1 = TR_85 ;
	7'h3f :
		RG_rl_73_t1 = TR_85 ;
	7'h40 :
		RG_rl_73_t1 = TR_85 ;
	7'h41 :
		RG_rl_73_t1 = TR_85 ;
	7'h42 :
		RG_rl_73_t1 = TR_85 ;
	7'h43 :
		RG_rl_73_t1 = TR_85 ;
	7'h44 :
		RG_rl_73_t1 = TR_85 ;
	7'h45 :
		RG_rl_73_t1 = TR_85 ;
	7'h46 :
		RG_rl_73_t1 = TR_85 ;
	7'h47 :
		RG_rl_73_t1 = TR_85 ;
	7'h48 :
		RG_rl_73_t1 = TR_85 ;
	7'h49 :
		RG_rl_73_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4a :
		RG_rl_73_t1 = TR_85 ;
	7'h4b :
		RG_rl_73_t1 = TR_85 ;
	7'h4c :
		RG_rl_73_t1 = TR_85 ;
	7'h4d :
		RG_rl_73_t1 = TR_85 ;
	7'h4e :
		RG_rl_73_t1 = TR_85 ;
	7'h4f :
		RG_rl_73_t1 = TR_85 ;
	7'h50 :
		RG_rl_73_t1 = TR_85 ;
	7'h51 :
		RG_rl_73_t1 = TR_85 ;
	7'h52 :
		RG_rl_73_t1 = TR_85 ;
	7'h53 :
		RG_rl_73_t1 = TR_85 ;
	7'h54 :
		RG_rl_73_t1 = TR_85 ;
	7'h55 :
		RG_rl_73_t1 = TR_85 ;
	7'h56 :
		RG_rl_73_t1 = TR_85 ;
	7'h57 :
		RG_rl_73_t1 = TR_85 ;
	7'h58 :
		RG_rl_73_t1 = TR_85 ;
	7'h59 :
		RG_rl_73_t1 = TR_85 ;
	7'h5a :
		RG_rl_73_t1 = TR_85 ;
	7'h5b :
		RG_rl_73_t1 = TR_85 ;
	7'h5c :
		RG_rl_73_t1 = TR_85 ;
	7'h5d :
		RG_rl_73_t1 = TR_85 ;
	7'h5e :
		RG_rl_73_t1 = TR_85 ;
	7'h5f :
		RG_rl_73_t1 = TR_85 ;
	7'h60 :
		RG_rl_73_t1 = TR_85 ;
	7'h61 :
		RG_rl_73_t1 = TR_85 ;
	7'h62 :
		RG_rl_73_t1 = TR_85 ;
	7'h63 :
		RG_rl_73_t1 = TR_85 ;
	7'h64 :
		RG_rl_73_t1 = TR_85 ;
	7'h65 :
		RG_rl_73_t1 = TR_85 ;
	7'h66 :
		RG_rl_73_t1 = TR_85 ;
	7'h67 :
		RG_rl_73_t1 = TR_85 ;
	7'h68 :
		RG_rl_73_t1 = TR_85 ;
	7'h69 :
		RG_rl_73_t1 = TR_85 ;
	7'h6a :
		RG_rl_73_t1 = TR_85 ;
	7'h6b :
		RG_rl_73_t1 = TR_85 ;
	7'h6c :
		RG_rl_73_t1 = TR_85 ;
	7'h6d :
		RG_rl_73_t1 = TR_85 ;
	7'h6e :
		RG_rl_73_t1 = TR_85 ;
	7'h6f :
		RG_rl_73_t1 = TR_85 ;
	7'h70 :
		RG_rl_73_t1 = TR_85 ;
	7'h71 :
		RG_rl_73_t1 = TR_85 ;
	7'h72 :
		RG_rl_73_t1 = TR_85 ;
	7'h73 :
		RG_rl_73_t1 = TR_85 ;
	7'h74 :
		RG_rl_73_t1 = TR_85 ;
	7'h75 :
		RG_rl_73_t1 = TR_85 ;
	7'h76 :
		RG_rl_73_t1 = TR_85 ;
	7'h77 :
		RG_rl_73_t1 = TR_85 ;
	7'h78 :
		RG_rl_73_t1 = TR_85 ;
	7'h79 :
		RG_rl_73_t1 = TR_85 ;
	7'h7a :
		RG_rl_73_t1 = TR_85 ;
	7'h7b :
		RG_rl_73_t1 = TR_85 ;
	7'h7c :
		RG_rl_73_t1 = TR_85 ;
	7'h7d :
		RG_rl_73_t1 = TR_85 ;
	7'h7e :
		RG_rl_73_t1 = TR_85 ;
	7'h7f :
		RG_rl_73_t1 = TR_85 ;
	default :
		RG_rl_73_t1 = 9'hx ;
	endcase
always @ ( RG_rl_73_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_14 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_73_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h49 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_73_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_14 )
		| ( { 9{ U_569 } } & RG_rl_73_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_73_en = ( U_570 | RG_rl_73_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_73_en )
		RG_rl_73 <= RG_rl_73_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_86 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_74_t1 = TR_86 ;
	7'h01 :
		RG_rl_74_t1 = TR_86 ;
	7'h02 :
		RG_rl_74_t1 = TR_86 ;
	7'h03 :
		RG_rl_74_t1 = TR_86 ;
	7'h04 :
		RG_rl_74_t1 = TR_86 ;
	7'h05 :
		RG_rl_74_t1 = TR_86 ;
	7'h06 :
		RG_rl_74_t1 = TR_86 ;
	7'h07 :
		RG_rl_74_t1 = TR_86 ;
	7'h08 :
		RG_rl_74_t1 = TR_86 ;
	7'h09 :
		RG_rl_74_t1 = TR_86 ;
	7'h0a :
		RG_rl_74_t1 = TR_86 ;
	7'h0b :
		RG_rl_74_t1 = TR_86 ;
	7'h0c :
		RG_rl_74_t1 = TR_86 ;
	7'h0d :
		RG_rl_74_t1 = TR_86 ;
	7'h0e :
		RG_rl_74_t1 = TR_86 ;
	7'h0f :
		RG_rl_74_t1 = TR_86 ;
	7'h10 :
		RG_rl_74_t1 = TR_86 ;
	7'h11 :
		RG_rl_74_t1 = TR_86 ;
	7'h12 :
		RG_rl_74_t1 = TR_86 ;
	7'h13 :
		RG_rl_74_t1 = TR_86 ;
	7'h14 :
		RG_rl_74_t1 = TR_86 ;
	7'h15 :
		RG_rl_74_t1 = TR_86 ;
	7'h16 :
		RG_rl_74_t1 = TR_86 ;
	7'h17 :
		RG_rl_74_t1 = TR_86 ;
	7'h18 :
		RG_rl_74_t1 = TR_86 ;
	7'h19 :
		RG_rl_74_t1 = TR_86 ;
	7'h1a :
		RG_rl_74_t1 = TR_86 ;
	7'h1b :
		RG_rl_74_t1 = TR_86 ;
	7'h1c :
		RG_rl_74_t1 = TR_86 ;
	7'h1d :
		RG_rl_74_t1 = TR_86 ;
	7'h1e :
		RG_rl_74_t1 = TR_86 ;
	7'h1f :
		RG_rl_74_t1 = TR_86 ;
	7'h20 :
		RG_rl_74_t1 = TR_86 ;
	7'h21 :
		RG_rl_74_t1 = TR_86 ;
	7'h22 :
		RG_rl_74_t1 = TR_86 ;
	7'h23 :
		RG_rl_74_t1 = TR_86 ;
	7'h24 :
		RG_rl_74_t1 = TR_86 ;
	7'h25 :
		RG_rl_74_t1 = TR_86 ;
	7'h26 :
		RG_rl_74_t1 = TR_86 ;
	7'h27 :
		RG_rl_74_t1 = TR_86 ;
	7'h28 :
		RG_rl_74_t1 = TR_86 ;
	7'h29 :
		RG_rl_74_t1 = TR_86 ;
	7'h2a :
		RG_rl_74_t1 = TR_86 ;
	7'h2b :
		RG_rl_74_t1 = TR_86 ;
	7'h2c :
		RG_rl_74_t1 = TR_86 ;
	7'h2d :
		RG_rl_74_t1 = TR_86 ;
	7'h2e :
		RG_rl_74_t1 = TR_86 ;
	7'h2f :
		RG_rl_74_t1 = TR_86 ;
	7'h30 :
		RG_rl_74_t1 = TR_86 ;
	7'h31 :
		RG_rl_74_t1 = TR_86 ;
	7'h32 :
		RG_rl_74_t1 = TR_86 ;
	7'h33 :
		RG_rl_74_t1 = TR_86 ;
	7'h34 :
		RG_rl_74_t1 = TR_86 ;
	7'h35 :
		RG_rl_74_t1 = TR_86 ;
	7'h36 :
		RG_rl_74_t1 = TR_86 ;
	7'h37 :
		RG_rl_74_t1 = TR_86 ;
	7'h38 :
		RG_rl_74_t1 = TR_86 ;
	7'h39 :
		RG_rl_74_t1 = TR_86 ;
	7'h3a :
		RG_rl_74_t1 = TR_86 ;
	7'h3b :
		RG_rl_74_t1 = TR_86 ;
	7'h3c :
		RG_rl_74_t1 = TR_86 ;
	7'h3d :
		RG_rl_74_t1 = TR_86 ;
	7'h3e :
		RG_rl_74_t1 = TR_86 ;
	7'h3f :
		RG_rl_74_t1 = TR_86 ;
	7'h40 :
		RG_rl_74_t1 = TR_86 ;
	7'h41 :
		RG_rl_74_t1 = TR_86 ;
	7'h42 :
		RG_rl_74_t1 = TR_86 ;
	7'h43 :
		RG_rl_74_t1 = TR_86 ;
	7'h44 :
		RG_rl_74_t1 = TR_86 ;
	7'h45 :
		RG_rl_74_t1 = TR_86 ;
	7'h46 :
		RG_rl_74_t1 = TR_86 ;
	7'h47 :
		RG_rl_74_t1 = TR_86 ;
	7'h48 :
		RG_rl_74_t1 = TR_86 ;
	7'h49 :
		RG_rl_74_t1 = TR_86 ;
	7'h4a :
		RG_rl_74_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4b :
		RG_rl_74_t1 = TR_86 ;
	7'h4c :
		RG_rl_74_t1 = TR_86 ;
	7'h4d :
		RG_rl_74_t1 = TR_86 ;
	7'h4e :
		RG_rl_74_t1 = TR_86 ;
	7'h4f :
		RG_rl_74_t1 = TR_86 ;
	7'h50 :
		RG_rl_74_t1 = TR_86 ;
	7'h51 :
		RG_rl_74_t1 = TR_86 ;
	7'h52 :
		RG_rl_74_t1 = TR_86 ;
	7'h53 :
		RG_rl_74_t1 = TR_86 ;
	7'h54 :
		RG_rl_74_t1 = TR_86 ;
	7'h55 :
		RG_rl_74_t1 = TR_86 ;
	7'h56 :
		RG_rl_74_t1 = TR_86 ;
	7'h57 :
		RG_rl_74_t1 = TR_86 ;
	7'h58 :
		RG_rl_74_t1 = TR_86 ;
	7'h59 :
		RG_rl_74_t1 = TR_86 ;
	7'h5a :
		RG_rl_74_t1 = TR_86 ;
	7'h5b :
		RG_rl_74_t1 = TR_86 ;
	7'h5c :
		RG_rl_74_t1 = TR_86 ;
	7'h5d :
		RG_rl_74_t1 = TR_86 ;
	7'h5e :
		RG_rl_74_t1 = TR_86 ;
	7'h5f :
		RG_rl_74_t1 = TR_86 ;
	7'h60 :
		RG_rl_74_t1 = TR_86 ;
	7'h61 :
		RG_rl_74_t1 = TR_86 ;
	7'h62 :
		RG_rl_74_t1 = TR_86 ;
	7'h63 :
		RG_rl_74_t1 = TR_86 ;
	7'h64 :
		RG_rl_74_t1 = TR_86 ;
	7'h65 :
		RG_rl_74_t1 = TR_86 ;
	7'h66 :
		RG_rl_74_t1 = TR_86 ;
	7'h67 :
		RG_rl_74_t1 = TR_86 ;
	7'h68 :
		RG_rl_74_t1 = TR_86 ;
	7'h69 :
		RG_rl_74_t1 = TR_86 ;
	7'h6a :
		RG_rl_74_t1 = TR_86 ;
	7'h6b :
		RG_rl_74_t1 = TR_86 ;
	7'h6c :
		RG_rl_74_t1 = TR_86 ;
	7'h6d :
		RG_rl_74_t1 = TR_86 ;
	7'h6e :
		RG_rl_74_t1 = TR_86 ;
	7'h6f :
		RG_rl_74_t1 = TR_86 ;
	7'h70 :
		RG_rl_74_t1 = TR_86 ;
	7'h71 :
		RG_rl_74_t1 = TR_86 ;
	7'h72 :
		RG_rl_74_t1 = TR_86 ;
	7'h73 :
		RG_rl_74_t1 = TR_86 ;
	7'h74 :
		RG_rl_74_t1 = TR_86 ;
	7'h75 :
		RG_rl_74_t1 = TR_86 ;
	7'h76 :
		RG_rl_74_t1 = TR_86 ;
	7'h77 :
		RG_rl_74_t1 = TR_86 ;
	7'h78 :
		RG_rl_74_t1 = TR_86 ;
	7'h79 :
		RG_rl_74_t1 = TR_86 ;
	7'h7a :
		RG_rl_74_t1 = TR_86 ;
	7'h7b :
		RG_rl_74_t1 = TR_86 ;
	7'h7c :
		RG_rl_74_t1 = TR_86 ;
	7'h7d :
		RG_rl_74_t1 = TR_86 ;
	7'h7e :
		RG_rl_74_t1 = TR_86 ;
	7'h7f :
		RG_rl_74_t1 = TR_86 ;
	default :
		RG_rl_74_t1 = 9'hx ;
	endcase
always @ ( RG_rl_74_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_15 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_74_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h4a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_74_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_15 )
		| ( { 9{ U_569 } } & RG_rl_74_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_74_en = ( U_570 | RG_rl_74_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_74_en )
		RG_rl_74 <= RG_rl_74_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_87 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_75_t1 = TR_87 ;
	7'h01 :
		RG_rl_75_t1 = TR_87 ;
	7'h02 :
		RG_rl_75_t1 = TR_87 ;
	7'h03 :
		RG_rl_75_t1 = TR_87 ;
	7'h04 :
		RG_rl_75_t1 = TR_87 ;
	7'h05 :
		RG_rl_75_t1 = TR_87 ;
	7'h06 :
		RG_rl_75_t1 = TR_87 ;
	7'h07 :
		RG_rl_75_t1 = TR_87 ;
	7'h08 :
		RG_rl_75_t1 = TR_87 ;
	7'h09 :
		RG_rl_75_t1 = TR_87 ;
	7'h0a :
		RG_rl_75_t1 = TR_87 ;
	7'h0b :
		RG_rl_75_t1 = TR_87 ;
	7'h0c :
		RG_rl_75_t1 = TR_87 ;
	7'h0d :
		RG_rl_75_t1 = TR_87 ;
	7'h0e :
		RG_rl_75_t1 = TR_87 ;
	7'h0f :
		RG_rl_75_t1 = TR_87 ;
	7'h10 :
		RG_rl_75_t1 = TR_87 ;
	7'h11 :
		RG_rl_75_t1 = TR_87 ;
	7'h12 :
		RG_rl_75_t1 = TR_87 ;
	7'h13 :
		RG_rl_75_t1 = TR_87 ;
	7'h14 :
		RG_rl_75_t1 = TR_87 ;
	7'h15 :
		RG_rl_75_t1 = TR_87 ;
	7'h16 :
		RG_rl_75_t1 = TR_87 ;
	7'h17 :
		RG_rl_75_t1 = TR_87 ;
	7'h18 :
		RG_rl_75_t1 = TR_87 ;
	7'h19 :
		RG_rl_75_t1 = TR_87 ;
	7'h1a :
		RG_rl_75_t1 = TR_87 ;
	7'h1b :
		RG_rl_75_t1 = TR_87 ;
	7'h1c :
		RG_rl_75_t1 = TR_87 ;
	7'h1d :
		RG_rl_75_t1 = TR_87 ;
	7'h1e :
		RG_rl_75_t1 = TR_87 ;
	7'h1f :
		RG_rl_75_t1 = TR_87 ;
	7'h20 :
		RG_rl_75_t1 = TR_87 ;
	7'h21 :
		RG_rl_75_t1 = TR_87 ;
	7'h22 :
		RG_rl_75_t1 = TR_87 ;
	7'h23 :
		RG_rl_75_t1 = TR_87 ;
	7'h24 :
		RG_rl_75_t1 = TR_87 ;
	7'h25 :
		RG_rl_75_t1 = TR_87 ;
	7'h26 :
		RG_rl_75_t1 = TR_87 ;
	7'h27 :
		RG_rl_75_t1 = TR_87 ;
	7'h28 :
		RG_rl_75_t1 = TR_87 ;
	7'h29 :
		RG_rl_75_t1 = TR_87 ;
	7'h2a :
		RG_rl_75_t1 = TR_87 ;
	7'h2b :
		RG_rl_75_t1 = TR_87 ;
	7'h2c :
		RG_rl_75_t1 = TR_87 ;
	7'h2d :
		RG_rl_75_t1 = TR_87 ;
	7'h2e :
		RG_rl_75_t1 = TR_87 ;
	7'h2f :
		RG_rl_75_t1 = TR_87 ;
	7'h30 :
		RG_rl_75_t1 = TR_87 ;
	7'h31 :
		RG_rl_75_t1 = TR_87 ;
	7'h32 :
		RG_rl_75_t1 = TR_87 ;
	7'h33 :
		RG_rl_75_t1 = TR_87 ;
	7'h34 :
		RG_rl_75_t1 = TR_87 ;
	7'h35 :
		RG_rl_75_t1 = TR_87 ;
	7'h36 :
		RG_rl_75_t1 = TR_87 ;
	7'h37 :
		RG_rl_75_t1 = TR_87 ;
	7'h38 :
		RG_rl_75_t1 = TR_87 ;
	7'h39 :
		RG_rl_75_t1 = TR_87 ;
	7'h3a :
		RG_rl_75_t1 = TR_87 ;
	7'h3b :
		RG_rl_75_t1 = TR_87 ;
	7'h3c :
		RG_rl_75_t1 = TR_87 ;
	7'h3d :
		RG_rl_75_t1 = TR_87 ;
	7'h3e :
		RG_rl_75_t1 = TR_87 ;
	7'h3f :
		RG_rl_75_t1 = TR_87 ;
	7'h40 :
		RG_rl_75_t1 = TR_87 ;
	7'h41 :
		RG_rl_75_t1 = TR_87 ;
	7'h42 :
		RG_rl_75_t1 = TR_87 ;
	7'h43 :
		RG_rl_75_t1 = TR_87 ;
	7'h44 :
		RG_rl_75_t1 = TR_87 ;
	7'h45 :
		RG_rl_75_t1 = TR_87 ;
	7'h46 :
		RG_rl_75_t1 = TR_87 ;
	7'h47 :
		RG_rl_75_t1 = TR_87 ;
	7'h48 :
		RG_rl_75_t1 = TR_87 ;
	7'h49 :
		RG_rl_75_t1 = TR_87 ;
	7'h4a :
		RG_rl_75_t1 = TR_87 ;
	7'h4b :
		RG_rl_75_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4c :
		RG_rl_75_t1 = TR_87 ;
	7'h4d :
		RG_rl_75_t1 = TR_87 ;
	7'h4e :
		RG_rl_75_t1 = TR_87 ;
	7'h4f :
		RG_rl_75_t1 = TR_87 ;
	7'h50 :
		RG_rl_75_t1 = TR_87 ;
	7'h51 :
		RG_rl_75_t1 = TR_87 ;
	7'h52 :
		RG_rl_75_t1 = TR_87 ;
	7'h53 :
		RG_rl_75_t1 = TR_87 ;
	7'h54 :
		RG_rl_75_t1 = TR_87 ;
	7'h55 :
		RG_rl_75_t1 = TR_87 ;
	7'h56 :
		RG_rl_75_t1 = TR_87 ;
	7'h57 :
		RG_rl_75_t1 = TR_87 ;
	7'h58 :
		RG_rl_75_t1 = TR_87 ;
	7'h59 :
		RG_rl_75_t1 = TR_87 ;
	7'h5a :
		RG_rl_75_t1 = TR_87 ;
	7'h5b :
		RG_rl_75_t1 = TR_87 ;
	7'h5c :
		RG_rl_75_t1 = TR_87 ;
	7'h5d :
		RG_rl_75_t1 = TR_87 ;
	7'h5e :
		RG_rl_75_t1 = TR_87 ;
	7'h5f :
		RG_rl_75_t1 = TR_87 ;
	7'h60 :
		RG_rl_75_t1 = TR_87 ;
	7'h61 :
		RG_rl_75_t1 = TR_87 ;
	7'h62 :
		RG_rl_75_t1 = TR_87 ;
	7'h63 :
		RG_rl_75_t1 = TR_87 ;
	7'h64 :
		RG_rl_75_t1 = TR_87 ;
	7'h65 :
		RG_rl_75_t1 = TR_87 ;
	7'h66 :
		RG_rl_75_t1 = TR_87 ;
	7'h67 :
		RG_rl_75_t1 = TR_87 ;
	7'h68 :
		RG_rl_75_t1 = TR_87 ;
	7'h69 :
		RG_rl_75_t1 = TR_87 ;
	7'h6a :
		RG_rl_75_t1 = TR_87 ;
	7'h6b :
		RG_rl_75_t1 = TR_87 ;
	7'h6c :
		RG_rl_75_t1 = TR_87 ;
	7'h6d :
		RG_rl_75_t1 = TR_87 ;
	7'h6e :
		RG_rl_75_t1 = TR_87 ;
	7'h6f :
		RG_rl_75_t1 = TR_87 ;
	7'h70 :
		RG_rl_75_t1 = TR_87 ;
	7'h71 :
		RG_rl_75_t1 = TR_87 ;
	7'h72 :
		RG_rl_75_t1 = TR_87 ;
	7'h73 :
		RG_rl_75_t1 = TR_87 ;
	7'h74 :
		RG_rl_75_t1 = TR_87 ;
	7'h75 :
		RG_rl_75_t1 = TR_87 ;
	7'h76 :
		RG_rl_75_t1 = TR_87 ;
	7'h77 :
		RG_rl_75_t1 = TR_87 ;
	7'h78 :
		RG_rl_75_t1 = TR_87 ;
	7'h79 :
		RG_rl_75_t1 = TR_87 ;
	7'h7a :
		RG_rl_75_t1 = TR_87 ;
	7'h7b :
		RG_rl_75_t1 = TR_87 ;
	7'h7c :
		RG_rl_75_t1 = TR_87 ;
	7'h7d :
		RG_rl_75_t1 = TR_87 ;
	7'h7e :
		RG_rl_75_t1 = TR_87 ;
	7'h7f :
		RG_rl_75_t1 = TR_87 ;
	default :
		RG_rl_75_t1 = 9'hx ;
	endcase
always @ ( RG_rl_75_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_16 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_75_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h4b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_75_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_16 )
		| ( { 9{ U_569 } } & RG_rl_75_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_75_en = ( U_570 | RG_rl_75_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_75_en )
		RG_rl_75 <= RG_rl_75_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_88 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_76_t1 = TR_88 ;
	7'h01 :
		RG_rl_76_t1 = TR_88 ;
	7'h02 :
		RG_rl_76_t1 = TR_88 ;
	7'h03 :
		RG_rl_76_t1 = TR_88 ;
	7'h04 :
		RG_rl_76_t1 = TR_88 ;
	7'h05 :
		RG_rl_76_t1 = TR_88 ;
	7'h06 :
		RG_rl_76_t1 = TR_88 ;
	7'h07 :
		RG_rl_76_t1 = TR_88 ;
	7'h08 :
		RG_rl_76_t1 = TR_88 ;
	7'h09 :
		RG_rl_76_t1 = TR_88 ;
	7'h0a :
		RG_rl_76_t1 = TR_88 ;
	7'h0b :
		RG_rl_76_t1 = TR_88 ;
	7'h0c :
		RG_rl_76_t1 = TR_88 ;
	7'h0d :
		RG_rl_76_t1 = TR_88 ;
	7'h0e :
		RG_rl_76_t1 = TR_88 ;
	7'h0f :
		RG_rl_76_t1 = TR_88 ;
	7'h10 :
		RG_rl_76_t1 = TR_88 ;
	7'h11 :
		RG_rl_76_t1 = TR_88 ;
	7'h12 :
		RG_rl_76_t1 = TR_88 ;
	7'h13 :
		RG_rl_76_t1 = TR_88 ;
	7'h14 :
		RG_rl_76_t1 = TR_88 ;
	7'h15 :
		RG_rl_76_t1 = TR_88 ;
	7'h16 :
		RG_rl_76_t1 = TR_88 ;
	7'h17 :
		RG_rl_76_t1 = TR_88 ;
	7'h18 :
		RG_rl_76_t1 = TR_88 ;
	7'h19 :
		RG_rl_76_t1 = TR_88 ;
	7'h1a :
		RG_rl_76_t1 = TR_88 ;
	7'h1b :
		RG_rl_76_t1 = TR_88 ;
	7'h1c :
		RG_rl_76_t1 = TR_88 ;
	7'h1d :
		RG_rl_76_t1 = TR_88 ;
	7'h1e :
		RG_rl_76_t1 = TR_88 ;
	7'h1f :
		RG_rl_76_t1 = TR_88 ;
	7'h20 :
		RG_rl_76_t1 = TR_88 ;
	7'h21 :
		RG_rl_76_t1 = TR_88 ;
	7'h22 :
		RG_rl_76_t1 = TR_88 ;
	7'h23 :
		RG_rl_76_t1 = TR_88 ;
	7'h24 :
		RG_rl_76_t1 = TR_88 ;
	7'h25 :
		RG_rl_76_t1 = TR_88 ;
	7'h26 :
		RG_rl_76_t1 = TR_88 ;
	7'h27 :
		RG_rl_76_t1 = TR_88 ;
	7'h28 :
		RG_rl_76_t1 = TR_88 ;
	7'h29 :
		RG_rl_76_t1 = TR_88 ;
	7'h2a :
		RG_rl_76_t1 = TR_88 ;
	7'h2b :
		RG_rl_76_t1 = TR_88 ;
	7'h2c :
		RG_rl_76_t1 = TR_88 ;
	7'h2d :
		RG_rl_76_t1 = TR_88 ;
	7'h2e :
		RG_rl_76_t1 = TR_88 ;
	7'h2f :
		RG_rl_76_t1 = TR_88 ;
	7'h30 :
		RG_rl_76_t1 = TR_88 ;
	7'h31 :
		RG_rl_76_t1 = TR_88 ;
	7'h32 :
		RG_rl_76_t1 = TR_88 ;
	7'h33 :
		RG_rl_76_t1 = TR_88 ;
	7'h34 :
		RG_rl_76_t1 = TR_88 ;
	7'h35 :
		RG_rl_76_t1 = TR_88 ;
	7'h36 :
		RG_rl_76_t1 = TR_88 ;
	7'h37 :
		RG_rl_76_t1 = TR_88 ;
	7'h38 :
		RG_rl_76_t1 = TR_88 ;
	7'h39 :
		RG_rl_76_t1 = TR_88 ;
	7'h3a :
		RG_rl_76_t1 = TR_88 ;
	7'h3b :
		RG_rl_76_t1 = TR_88 ;
	7'h3c :
		RG_rl_76_t1 = TR_88 ;
	7'h3d :
		RG_rl_76_t1 = TR_88 ;
	7'h3e :
		RG_rl_76_t1 = TR_88 ;
	7'h3f :
		RG_rl_76_t1 = TR_88 ;
	7'h40 :
		RG_rl_76_t1 = TR_88 ;
	7'h41 :
		RG_rl_76_t1 = TR_88 ;
	7'h42 :
		RG_rl_76_t1 = TR_88 ;
	7'h43 :
		RG_rl_76_t1 = TR_88 ;
	7'h44 :
		RG_rl_76_t1 = TR_88 ;
	7'h45 :
		RG_rl_76_t1 = TR_88 ;
	7'h46 :
		RG_rl_76_t1 = TR_88 ;
	7'h47 :
		RG_rl_76_t1 = TR_88 ;
	7'h48 :
		RG_rl_76_t1 = TR_88 ;
	7'h49 :
		RG_rl_76_t1 = TR_88 ;
	7'h4a :
		RG_rl_76_t1 = TR_88 ;
	7'h4b :
		RG_rl_76_t1 = TR_88 ;
	7'h4c :
		RG_rl_76_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4d :
		RG_rl_76_t1 = TR_88 ;
	7'h4e :
		RG_rl_76_t1 = TR_88 ;
	7'h4f :
		RG_rl_76_t1 = TR_88 ;
	7'h50 :
		RG_rl_76_t1 = TR_88 ;
	7'h51 :
		RG_rl_76_t1 = TR_88 ;
	7'h52 :
		RG_rl_76_t1 = TR_88 ;
	7'h53 :
		RG_rl_76_t1 = TR_88 ;
	7'h54 :
		RG_rl_76_t1 = TR_88 ;
	7'h55 :
		RG_rl_76_t1 = TR_88 ;
	7'h56 :
		RG_rl_76_t1 = TR_88 ;
	7'h57 :
		RG_rl_76_t1 = TR_88 ;
	7'h58 :
		RG_rl_76_t1 = TR_88 ;
	7'h59 :
		RG_rl_76_t1 = TR_88 ;
	7'h5a :
		RG_rl_76_t1 = TR_88 ;
	7'h5b :
		RG_rl_76_t1 = TR_88 ;
	7'h5c :
		RG_rl_76_t1 = TR_88 ;
	7'h5d :
		RG_rl_76_t1 = TR_88 ;
	7'h5e :
		RG_rl_76_t1 = TR_88 ;
	7'h5f :
		RG_rl_76_t1 = TR_88 ;
	7'h60 :
		RG_rl_76_t1 = TR_88 ;
	7'h61 :
		RG_rl_76_t1 = TR_88 ;
	7'h62 :
		RG_rl_76_t1 = TR_88 ;
	7'h63 :
		RG_rl_76_t1 = TR_88 ;
	7'h64 :
		RG_rl_76_t1 = TR_88 ;
	7'h65 :
		RG_rl_76_t1 = TR_88 ;
	7'h66 :
		RG_rl_76_t1 = TR_88 ;
	7'h67 :
		RG_rl_76_t1 = TR_88 ;
	7'h68 :
		RG_rl_76_t1 = TR_88 ;
	7'h69 :
		RG_rl_76_t1 = TR_88 ;
	7'h6a :
		RG_rl_76_t1 = TR_88 ;
	7'h6b :
		RG_rl_76_t1 = TR_88 ;
	7'h6c :
		RG_rl_76_t1 = TR_88 ;
	7'h6d :
		RG_rl_76_t1 = TR_88 ;
	7'h6e :
		RG_rl_76_t1 = TR_88 ;
	7'h6f :
		RG_rl_76_t1 = TR_88 ;
	7'h70 :
		RG_rl_76_t1 = TR_88 ;
	7'h71 :
		RG_rl_76_t1 = TR_88 ;
	7'h72 :
		RG_rl_76_t1 = TR_88 ;
	7'h73 :
		RG_rl_76_t1 = TR_88 ;
	7'h74 :
		RG_rl_76_t1 = TR_88 ;
	7'h75 :
		RG_rl_76_t1 = TR_88 ;
	7'h76 :
		RG_rl_76_t1 = TR_88 ;
	7'h77 :
		RG_rl_76_t1 = TR_88 ;
	7'h78 :
		RG_rl_76_t1 = TR_88 ;
	7'h79 :
		RG_rl_76_t1 = TR_88 ;
	7'h7a :
		RG_rl_76_t1 = TR_88 ;
	7'h7b :
		RG_rl_76_t1 = TR_88 ;
	7'h7c :
		RG_rl_76_t1 = TR_88 ;
	7'h7d :
		RG_rl_76_t1 = TR_88 ;
	7'h7e :
		RG_rl_76_t1 = TR_88 ;
	7'h7f :
		RG_rl_76_t1 = TR_88 ;
	default :
		RG_rl_76_t1 = 9'hx ;
	endcase
always @ ( RG_rl_76_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_17 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_76_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h4c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_76_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_17 )
		| ( { 9{ U_569 } } & RG_rl_76_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_76_en = ( U_570 | RG_rl_76_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_76_en )
		RG_rl_76 <= RG_rl_76_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_89 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_77_t1 = TR_89 ;
	7'h01 :
		RG_rl_77_t1 = TR_89 ;
	7'h02 :
		RG_rl_77_t1 = TR_89 ;
	7'h03 :
		RG_rl_77_t1 = TR_89 ;
	7'h04 :
		RG_rl_77_t1 = TR_89 ;
	7'h05 :
		RG_rl_77_t1 = TR_89 ;
	7'h06 :
		RG_rl_77_t1 = TR_89 ;
	7'h07 :
		RG_rl_77_t1 = TR_89 ;
	7'h08 :
		RG_rl_77_t1 = TR_89 ;
	7'h09 :
		RG_rl_77_t1 = TR_89 ;
	7'h0a :
		RG_rl_77_t1 = TR_89 ;
	7'h0b :
		RG_rl_77_t1 = TR_89 ;
	7'h0c :
		RG_rl_77_t1 = TR_89 ;
	7'h0d :
		RG_rl_77_t1 = TR_89 ;
	7'h0e :
		RG_rl_77_t1 = TR_89 ;
	7'h0f :
		RG_rl_77_t1 = TR_89 ;
	7'h10 :
		RG_rl_77_t1 = TR_89 ;
	7'h11 :
		RG_rl_77_t1 = TR_89 ;
	7'h12 :
		RG_rl_77_t1 = TR_89 ;
	7'h13 :
		RG_rl_77_t1 = TR_89 ;
	7'h14 :
		RG_rl_77_t1 = TR_89 ;
	7'h15 :
		RG_rl_77_t1 = TR_89 ;
	7'h16 :
		RG_rl_77_t1 = TR_89 ;
	7'h17 :
		RG_rl_77_t1 = TR_89 ;
	7'h18 :
		RG_rl_77_t1 = TR_89 ;
	7'h19 :
		RG_rl_77_t1 = TR_89 ;
	7'h1a :
		RG_rl_77_t1 = TR_89 ;
	7'h1b :
		RG_rl_77_t1 = TR_89 ;
	7'h1c :
		RG_rl_77_t1 = TR_89 ;
	7'h1d :
		RG_rl_77_t1 = TR_89 ;
	7'h1e :
		RG_rl_77_t1 = TR_89 ;
	7'h1f :
		RG_rl_77_t1 = TR_89 ;
	7'h20 :
		RG_rl_77_t1 = TR_89 ;
	7'h21 :
		RG_rl_77_t1 = TR_89 ;
	7'h22 :
		RG_rl_77_t1 = TR_89 ;
	7'h23 :
		RG_rl_77_t1 = TR_89 ;
	7'h24 :
		RG_rl_77_t1 = TR_89 ;
	7'h25 :
		RG_rl_77_t1 = TR_89 ;
	7'h26 :
		RG_rl_77_t1 = TR_89 ;
	7'h27 :
		RG_rl_77_t1 = TR_89 ;
	7'h28 :
		RG_rl_77_t1 = TR_89 ;
	7'h29 :
		RG_rl_77_t1 = TR_89 ;
	7'h2a :
		RG_rl_77_t1 = TR_89 ;
	7'h2b :
		RG_rl_77_t1 = TR_89 ;
	7'h2c :
		RG_rl_77_t1 = TR_89 ;
	7'h2d :
		RG_rl_77_t1 = TR_89 ;
	7'h2e :
		RG_rl_77_t1 = TR_89 ;
	7'h2f :
		RG_rl_77_t1 = TR_89 ;
	7'h30 :
		RG_rl_77_t1 = TR_89 ;
	7'h31 :
		RG_rl_77_t1 = TR_89 ;
	7'h32 :
		RG_rl_77_t1 = TR_89 ;
	7'h33 :
		RG_rl_77_t1 = TR_89 ;
	7'h34 :
		RG_rl_77_t1 = TR_89 ;
	7'h35 :
		RG_rl_77_t1 = TR_89 ;
	7'h36 :
		RG_rl_77_t1 = TR_89 ;
	7'h37 :
		RG_rl_77_t1 = TR_89 ;
	7'h38 :
		RG_rl_77_t1 = TR_89 ;
	7'h39 :
		RG_rl_77_t1 = TR_89 ;
	7'h3a :
		RG_rl_77_t1 = TR_89 ;
	7'h3b :
		RG_rl_77_t1 = TR_89 ;
	7'h3c :
		RG_rl_77_t1 = TR_89 ;
	7'h3d :
		RG_rl_77_t1 = TR_89 ;
	7'h3e :
		RG_rl_77_t1 = TR_89 ;
	7'h3f :
		RG_rl_77_t1 = TR_89 ;
	7'h40 :
		RG_rl_77_t1 = TR_89 ;
	7'h41 :
		RG_rl_77_t1 = TR_89 ;
	7'h42 :
		RG_rl_77_t1 = TR_89 ;
	7'h43 :
		RG_rl_77_t1 = TR_89 ;
	7'h44 :
		RG_rl_77_t1 = TR_89 ;
	7'h45 :
		RG_rl_77_t1 = TR_89 ;
	7'h46 :
		RG_rl_77_t1 = TR_89 ;
	7'h47 :
		RG_rl_77_t1 = TR_89 ;
	7'h48 :
		RG_rl_77_t1 = TR_89 ;
	7'h49 :
		RG_rl_77_t1 = TR_89 ;
	7'h4a :
		RG_rl_77_t1 = TR_89 ;
	7'h4b :
		RG_rl_77_t1 = TR_89 ;
	7'h4c :
		RG_rl_77_t1 = TR_89 ;
	7'h4d :
		RG_rl_77_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4e :
		RG_rl_77_t1 = TR_89 ;
	7'h4f :
		RG_rl_77_t1 = TR_89 ;
	7'h50 :
		RG_rl_77_t1 = TR_89 ;
	7'h51 :
		RG_rl_77_t1 = TR_89 ;
	7'h52 :
		RG_rl_77_t1 = TR_89 ;
	7'h53 :
		RG_rl_77_t1 = TR_89 ;
	7'h54 :
		RG_rl_77_t1 = TR_89 ;
	7'h55 :
		RG_rl_77_t1 = TR_89 ;
	7'h56 :
		RG_rl_77_t1 = TR_89 ;
	7'h57 :
		RG_rl_77_t1 = TR_89 ;
	7'h58 :
		RG_rl_77_t1 = TR_89 ;
	7'h59 :
		RG_rl_77_t1 = TR_89 ;
	7'h5a :
		RG_rl_77_t1 = TR_89 ;
	7'h5b :
		RG_rl_77_t1 = TR_89 ;
	7'h5c :
		RG_rl_77_t1 = TR_89 ;
	7'h5d :
		RG_rl_77_t1 = TR_89 ;
	7'h5e :
		RG_rl_77_t1 = TR_89 ;
	7'h5f :
		RG_rl_77_t1 = TR_89 ;
	7'h60 :
		RG_rl_77_t1 = TR_89 ;
	7'h61 :
		RG_rl_77_t1 = TR_89 ;
	7'h62 :
		RG_rl_77_t1 = TR_89 ;
	7'h63 :
		RG_rl_77_t1 = TR_89 ;
	7'h64 :
		RG_rl_77_t1 = TR_89 ;
	7'h65 :
		RG_rl_77_t1 = TR_89 ;
	7'h66 :
		RG_rl_77_t1 = TR_89 ;
	7'h67 :
		RG_rl_77_t1 = TR_89 ;
	7'h68 :
		RG_rl_77_t1 = TR_89 ;
	7'h69 :
		RG_rl_77_t1 = TR_89 ;
	7'h6a :
		RG_rl_77_t1 = TR_89 ;
	7'h6b :
		RG_rl_77_t1 = TR_89 ;
	7'h6c :
		RG_rl_77_t1 = TR_89 ;
	7'h6d :
		RG_rl_77_t1 = TR_89 ;
	7'h6e :
		RG_rl_77_t1 = TR_89 ;
	7'h6f :
		RG_rl_77_t1 = TR_89 ;
	7'h70 :
		RG_rl_77_t1 = TR_89 ;
	7'h71 :
		RG_rl_77_t1 = TR_89 ;
	7'h72 :
		RG_rl_77_t1 = TR_89 ;
	7'h73 :
		RG_rl_77_t1 = TR_89 ;
	7'h74 :
		RG_rl_77_t1 = TR_89 ;
	7'h75 :
		RG_rl_77_t1 = TR_89 ;
	7'h76 :
		RG_rl_77_t1 = TR_89 ;
	7'h77 :
		RG_rl_77_t1 = TR_89 ;
	7'h78 :
		RG_rl_77_t1 = TR_89 ;
	7'h79 :
		RG_rl_77_t1 = TR_89 ;
	7'h7a :
		RG_rl_77_t1 = TR_89 ;
	7'h7b :
		RG_rl_77_t1 = TR_89 ;
	7'h7c :
		RG_rl_77_t1 = TR_89 ;
	7'h7d :
		RG_rl_77_t1 = TR_89 ;
	7'h7e :
		RG_rl_77_t1 = TR_89 ;
	7'h7f :
		RG_rl_77_t1 = TR_89 ;
	default :
		RG_rl_77_t1 = 9'hx ;
	endcase
always @ ( RG_rl_77_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_18 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_77_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h4d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_77_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_18 )
		| ( { 9{ U_569 } } & RG_rl_77_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_77_en = ( U_570 | RG_rl_77_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_77_en )
		RG_rl_77 <= RG_rl_77_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_90 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_78_t1 = TR_90 ;
	7'h01 :
		RG_rl_78_t1 = TR_90 ;
	7'h02 :
		RG_rl_78_t1 = TR_90 ;
	7'h03 :
		RG_rl_78_t1 = TR_90 ;
	7'h04 :
		RG_rl_78_t1 = TR_90 ;
	7'h05 :
		RG_rl_78_t1 = TR_90 ;
	7'h06 :
		RG_rl_78_t1 = TR_90 ;
	7'h07 :
		RG_rl_78_t1 = TR_90 ;
	7'h08 :
		RG_rl_78_t1 = TR_90 ;
	7'h09 :
		RG_rl_78_t1 = TR_90 ;
	7'h0a :
		RG_rl_78_t1 = TR_90 ;
	7'h0b :
		RG_rl_78_t1 = TR_90 ;
	7'h0c :
		RG_rl_78_t1 = TR_90 ;
	7'h0d :
		RG_rl_78_t1 = TR_90 ;
	7'h0e :
		RG_rl_78_t1 = TR_90 ;
	7'h0f :
		RG_rl_78_t1 = TR_90 ;
	7'h10 :
		RG_rl_78_t1 = TR_90 ;
	7'h11 :
		RG_rl_78_t1 = TR_90 ;
	7'h12 :
		RG_rl_78_t1 = TR_90 ;
	7'h13 :
		RG_rl_78_t1 = TR_90 ;
	7'h14 :
		RG_rl_78_t1 = TR_90 ;
	7'h15 :
		RG_rl_78_t1 = TR_90 ;
	7'h16 :
		RG_rl_78_t1 = TR_90 ;
	7'h17 :
		RG_rl_78_t1 = TR_90 ;
	7'h18 :
		RG_rl_78_t1 = TR_90 ;
	7'h19 :
		RG_rl_78_t1 = TR_90 ;
	7'h1a :
		RG_rl_78_t1 = TR_90 ;
	7'h1b :
		RG_rl_78_t1 = TR_90 ;
	7'h1c :
		RG_rl_78_t1 = TR_90 ;
	7'h1d :
		RG_rl_78_t1 = TR_90 ;
	7'h1e :
		RG_rl_78_t1 = TR_90 ;
	7'h1f :
		RG_rl_78_t1 = TR_90 ;
	7'h20 :
		RG_rl_78_t1 = TR_90 ;
	7'h21 :
		RG_rl_78_t1 = TR_90 ;
	7'h22 :
		RG_rl_78_t1 = TR_90 ;
	7'h23 :
		RG_rl_78_t1 = TR_90 ;
	7'h24 :
		RG_rl_78_t1 = TR_90 ;
	7'h25 :
		RG_rl_78_t1 = TR_90 ;
	7'h26 :
		RG_rl_78_t1 = TR_90 ;
	7'h27 :
		RG_rl_78_t1 = TR_90 ;
	7'h28 :
		RG_rl_78_t1 = TR_90 ;
	7'h29 :
		RG_rl_78_t1 = TR_90 ;
	7'h2a :
		RG_rl_78_t1 = TR_90 ;
	7'h2b :
		RG_rl_78_t1 = TR_90 ;
	7'h2c :
		RG_rl_78_t1 = TR_90 ;
	7'h2d :
		RG_rl_78_t1 = TR_90 ;
	7'h2e :
		RG_rl_78_t1 = TR_90 ;
	7'h2f :
		RG_rl_78_t1 = TR_90 ;
	7'h30 :
		RG_rl_78_t1 = TR_90 ;
	7'h31 :
		RG_rl_78_t1 = TR_90 ;
	7'h32 :
		RG_rl_78_t1 = TR_90 ;
	7'h33 :
		RG_rl_78_t1 = TR_90 ;
	7'h34 :
		RG_rl_78_t1 = TR_90 ;
	7'h35 :
		RG_rl_78_t1 = TR_90 ;
	7'h36 :
		RG_rl_78_t1 = TR_90 ;
	7'h37 :
		RG_rl_78_t1 = TR_90 ;
	7'h38 :
		RG_rl_78_t1 = TR_90 ;
	7'h39 :
		RG_rl_78_t1 = TR_90 ;
	7'h3a :
		RG_rl_78_t1 = TR_90 ;
	7'h3b :
		RG_rl_78_t1 = TR_90 ;
	7'h3c :
		RG_rl_78_t1 = TR_90 ;
	7'h3d :
		RG_rl_78_t1 = TR_90 ;
	7'h3e :
		RG_rl_78_t1 = TR_90 ;
	7'h3f :
		RG_rl_78_t1 = TR_90 ;
	7'h40 :
		RG_rl_78_t1 = TR_90 ;
	7'h41 :
		RG_rl_78_t1 = TR_90 ;
	7'h42 :
		RG_rl_78_t1 = TR_90 ;
	7'h43 :
		RG_rl_78_t1 = TR_90 ;
	7'h44 :
		RG_rl_78_t1 = TR_90 ;
	7'h45 :
		RG_rl_78_t1 = TR_90 ;
	7'h46 :
		RG_rl_78_t1 = TR_90 ;
	7'h47 :
		RG_rl_78_t1 = TR_90 ;
	7'h48 :
		RG_rl_78_t1 = TR_90 ;
	7'h49 :
		RG_rl_78_t1 = TR_90 ;
	7'h4a :
		RG_rl_78_t1 = TR_90 ;
	7'h4b :
		RG_rl_78_t1 = TR_90 ;
	7'h4c :
		RG_rl_78_t1 = TR_90 ;
	7'h4d :
		RG_rl_78_t1 = TR_90 ;
	7'h4e :
		RG_rl_78_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h4f :
		RG_rl_78_t1 = TR_90 ;
	7'h50 :
		RG_rl_78_t1 = TR_90 ;
	7'h51 :
		RG_rl_78_t1 = TR_90 ;
	7'h52 :
		RG_rl_78_t1 = TR_90 ;
	7'h53 :
		RG_rl_78_t1 = TR_90 ;
	7'h54 :
		RG_rl_78_t1 = TR_90 ;
	7'h55 :
		RG_rl_78_t1 = TR_90 ;
	7'h56 :
		RG_rl_78_t1 = TR_90 ;
	7'h57 :
		RG_rl_78_t1 = TR_90 ;
	7'h58 :
		RG_rl_78_t1 = TR_90 ;
	7'h59 :
		RG_rl_78_t1 = TR_90 ;
	7'h5a :
		RG_rl_78_t1 = TR_90 ;
	7'h5b :
		RG_rl_78_t1 = TR_90 ;
	7'h5c :
		RG_rl_78_t1 = TR_90 ;
	7'h5d :
		RG_rl_78_t1 = TR_90 ;
	7'h5e :
		RG_rl_78_t1 = TR_90 ;
	7'h5f :
		RG_rl_78_t1 = TR_90 ;
	7'h60 :
		RG_rl_78_t1 = TR_90 ;
	7'h61 :
		RG_rl_78_t1 = TR_90 ;
	7'h62 :
		RG_rl_78_t1 = TR_90 ;
	7'h63 :
		RG_rl_78_t1 = TR_90 ;
	7'h64 :
		RG_rl_78_t1 = TR_90 ;
	7'h65 :
		RG_rl_78_t1 = TR_90 ;
	7'h66 :
		RG_rl_78_t1 = TR_90 ;
	7'h67 :
		RG_rl_78_t1 = TR_90 ;
	7'h68 :
		RG_rl_78_t1 = TR_90 ;
	7'h69 :
		RG_rl_78_t1 = TR_90 ;
	7'h6a :
		RG_rl_78_t1 = TR_90 ;
	7'h6b :
		RG_rl_78_t1 = TR_90 ;
	7'h6c :
		RG_rl_78_t1 = TR_90 ;
	7'h6d :
		RG_rl_78_t1 = TR_90 ;
	7'h6e :
		RG_rl_78_t1 = TR_90 ;
	7'h6f :
		RG_rl_78_t1 = TR_90 ;
	7'h70 :
		RG_rl_78_t1 = TR_90 ;
	7'h71 :
		RG_rl_78_t1 = TR_90 ;
	7'h72 :
		RG_rl_78_t1 = TR_90 ;
	7'h73 :
		RG_rl_78_t1 = TR_90 ;
	7'h74 :
		RG_rl_78_t1 = TR_90 ;
	7'h75 :
		RG_rl_78_t1 = TR_90 ;
	7'h76 :
		RG_rl_78_t1 = TR_90 ;
	7'h77 :
		RG_rl_78_t1 = TR_90 ;
	7'h78 :
		RG_rl_78_t1 = TR_90 ;
	7'h79 :
		RG_rl_78_t1 = TR_90 ;
	7'h7a :
		RG_rl_78_t1 = TR_90 ;
	7'h7b :
		RG_rl_78_t1 = TR_90 ;
	7'h7c :
		RG_rl_78_t1 = TR_90 ;
	7'h7d :
		RG_rl_78_t1 = TR_90 ;
	7'h7e :
		RG_rl_78_t1 = TR_90 ;
	7'h7f :
		RG_rl_78_t1 = TR_90 ;
	default :
		RG_rl_78_t1 = 9'hx ;
	endcase
always @ ( RG_rl_78_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_19 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_78_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h4e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_78_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_19 )
		| ( { 9{ U_569 } } & RG_rl_78_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_78_en = ( U_570 | RG_rl_78_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_78_en )
		RG_rl_78 <= RG_rl_78_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_91 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_79_t1 = TR_91 ;
	7'h01 :
		RG_rl_79_t1 = TR_91 ;
	7'h02 :
		RG_rl_79_t1 = TR_91 ;
	7'h03 :
		RG_rl_79_t1 = TR_91 ;
	7'h04 :
		RG_rl_79_t1 = TR_91 ;
	7'h05 :
		RG_rl_79_t1 = TR_91 ;
	7'h06 :
		RG_rl_79_t1 = TR_91 ;
	7'h07 :
		RG_rl_79_t1 = TR_91 ;
	7'h08 :
		RG_rl_79_t1 = TR_91 ;
	7'h09 :
		RG_rl_79_t1 = TR_91 ;
	7'h0a :
		RG_rl_79_t1 = TR_91 ;
	7'h0b :
		RG_rl_79_t1 = TR_91 ;
	7'h0c :
		RG_rl_79_t1 = TR_91 ;
	7'h0d :
		RG_rl_79_t1 = TR_91 ;
	7'h0e :
		RG_rl_79_t1 = TR_91 ;
	7'h0f :
		RG_rl_79_t1 = TR_91 ;
	7'h10 :
		RG_rl_79_t1 = TR_91 ;
	7'h11 :
		RG_rl_79_t1 = TR_91 ;
	7'h12 :
		RG_rl_79_t1 = TR_91 ;
	7'h13 :
		RG_rl_79_t1 = TR_91 ;
	7'h14 :
		RG_rl_79_t1 = TR_91 ;
	7'h15 :
		RG_rl_79_t1 = TR_91 ;
	7'h16 :
		RG_rl_79_t1 = TR_91 ;
	7'h17 :
		RG_rl_79_t1 = TR_91 ;
	7'h18 :
		RG_rl_79_t1 = TR_91 ;
	7'h19 :
		RG_rl_79_t1 = TR_91 ;
	7'h1a :
		RG_rl_79_t1 = TR_91 ;
	7'h1b :
		RG_rl_79_t1 = TR_91 ;
	7'h1c :
		RG_rl_79_t1 = TR_91 ;
	7'h1d :
		RG_rl_79_t1 = TR_91 ;
	7'h1e :
		RG_rl_79_t1 = TR_91 ;
	7'h1f :
		RG_rl_79_t1 = TR_91 ;
	7'h20 :
		RG_rl_79_t1 = TR_91 ;
	7'h21 :
		RG_rl_79_t1 = TR_91 ;
	7'h22 :
		RG_rl_79_t1 = TR_91 ;
	7'h23 :
		RG_rl_79_t1 = TR_91 ;
	7'h24 :
		RG_rl_79_t1 = TR_91 ;
	7'h25 :
		RG_rl_79_t1 = TR_91 ;
	7'h26 :
		RG_rl_79_t1 = TR_91 ;
	7'h27 :
		RG_rl_79_t1 = TR_91 ;
	7'h28 :
		RG_rl_79_t1 = TR_91 ;
	7'h29 :
		RG_rl_79_t1 = TR_91 ;
	7'h2a :
		RG_rl_79_t1 = TR_91 ;
	7'h2b :
		RG_rl_79_t1 = TR_91 ;
	7'h2c :
		RG_rl_79_t1 = TR_91 ;
	7'h2d :
		RG_rl_79_t1 = TR_91 ;
	7'h2e :
		RG_rl_79_t1 = TR_91 ;
	7'h2f :
		RG_rl_79_t1 = TR_91 ;
	7'h30 :
		RG_rl_79_t1 = TR_91 ;
	7'h31 :
		RG_rl_79_t1 = TR_91 ;
	7'h32 :
		RG_rl_79_t1 = TR_91 ;
	7'h33 :
		RG_rl_79_t1 = TR_91 ;
	7'h34 :
		RG_rl_79_t1 = TR_91 ;
	7'h35 :
		RG_rl_79_t1 = TR_91 ;
	7'h36 :
		RG_rl_79_t1 = TR_91 ;
	7'h37 :
		RG_rl_79_t1 = TR_91 ;
	7'h38 :
		RG_rl_79_t1 = TR_91 ;
	7'h39 :
		RG_rl_79_t1 = TR_91 ;
	7'h3a :
		RG_rl_79_t1 = TR_91 ;
	7'h3b :
		RG_rl_79_t1 = TR_91 ;
	7'h3c :
		RG_rl_79_t1 = TR_91 ;
	7'h3d :
		RG_rl_79_t1 = TR_91 ;
	7'h3e :
		RG_rl_79_t1 = TR_91 ;
	7'h3f :
		RG_rl_79_t1 = TR_91 ;
	7'h40 :
		RG_rl_79_t1 = TR_91 ;
	7'h41 :
		RG_rl_79_t1 = TR_91 ;
	7'h42 :
		RG_rl_79_t1 = TR_91 ;
	7'h43 :
		RG_rl_79_t1 = TR_91 ;
	7'h44 :
		RG_rl_79_t1 = TR_91 ;
	7'h45 :
		RG_rl_79_t1 = TR_91 ;
	7'h46 :
		RG_rl_79_t1 = TR_91 ;
	7'h47 :
		RG_rl_79_t1 = TR_91 ;
	7'h48 :
		RG_rl_79_t1 = TR_91 ;
	7'h49 :
		RG_rl_79_t1 = TR_91 ;
	7'h4a :
		RG_rl_79_t1 = TR_91 ;
	7'h4b :
		RG_rl_79_t1 = TR_91 ;
	7'h4c :
		RG_rl_79_t1 = TR_91 ;
	7'h4d :
		RG_rl_79_t1 = TR_91 ;
	7'h4e :
		RG_rl_79_t1 = TR_91 ;
	7'h4f :
		RG_rl_79_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h50 :
		RG_rl_79_t1 = TR_91 ;
	7'h51 :
		RG_rl_79_t1 = TR_91 ;
	7'h52 :
		RG_rl_79_t1 = TR_91 ;
	7'h53 :
		RG_rl_79_t1 = TR_91 ;
	7'h54 :
		RG_rl_79_t1 = TR_91 ;
	7'h55 :
		RG_rl_79_t1 = TR_91 ;
	7'h56 :
		RG_rl_79_t1 = TR_91 ;
	7'h57 :
		RG_rl_79_t1 = TR_91 ;
	7'h58 :
		RG_rl_79_t1 = TR_91 ;
	7'h59 :
		RG_rl_79_t1 = TR_91 ;
	7'h5a :
		RG_rl_79_t1 = TR_91 ;
	7'h5b :
		RG_rl_79_t1 = TR_91 ;
	7'h5c :
		RG_rl_79_t1 = TR_91 ;
	7'h5d :
		RG_rl_79_t1 = TR_91 ;
	7'h5e :
		RG_rl_79_t1 = TR_91 ;
	7'h5f :
		RG_rl_79_t1 = TR_91 ;
	7'h60 :
		RG_rl_79_t1 = TR_91 ;
	7'h61 :
		RG_rl_79_t1 = TR_91 ;
	7'h62 :
		RG_rl_79_t1 = TR_91 ;
	7'h63 :
		RG_rl_79_t1 = TR_91 ;
	7'h64 :
		RG_rl_79_t1 = TR_91 ;
	7'h65 :
		RG_rl_79_t1 = TR_91 ;
	7'h66 :
		RG_rl_79_t1 = TR_91 ;
	7'h67 :
		RG_rl_79_t1 = TR_91 ;
	7'h68 :
		RG_rl_79_t1 = TR_91 ;
	7'h69 :
		RG_rl_79_t1 = TR_91 ;
	7'h6a :
		RG_rl_79_t1 = TR_91 ;
	7'h6b :
		RG_rl_79_t1 = TR_91 ;
	7'h6c :
		RG_rl_79_t1 = TR_91 ;
	7'h6d :
		RG_rl_79_t1 = TR_91 ;
	7'h6e :
		RG_rl_79_t1 = TR_91 ;
	7'h6f :
		RG_rl_79_t1 = TR_91 ;
	7'h70 :
		RG_rl_79_t1 = TR_91 ;
	7'h71 :
		RG_rl_79_t1 = TR_91 ;
	7'h72 :
		RG_rl_79_t1 = TR_91 ;
	7'h73 :
		RG_rl_79_t1 = TR_91 ;
	7'h74 :
		RG_rl_79_t1 = TR_91 ;
	7'h75 :
		RG_rl_79_t1 = TR_91 ;
	7'h76 :
		RG_rl_79_t1 = TR_91 ;
	7'h77 :
		RG_rl_79_t1 = TR_91 ;
	7'h78 :
		RG_rl_79_t1 = TR_91 ;
	7'h79 :
		RG_rl_79_t1 = TR_91 ;
	7'h7a :
		RG_rl_79_t1 = TR_91 ;
	7'h7b :
		RG_rl_79_t1 = TR_91 ;
	7'h7c :
		RG_rl_79_t1 = TR_91 ;
	7'h7d :
		RG_rl_79_t1 = TR_91 ;
	7'h7e :
		RG_rl_79_t1 = TR_91 ;
	7'h7f :
		RG_rl_79_t1 = TR_91 ;
	default :
		RG_rl_79_t1 = 9'hx ;
	endcase
always @ ( RG_rl_79_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_20 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_79_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h4f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_79_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_20 )
		| ( { 9{ U_569 } } & RG_rl_79_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_79_en = ( U_570 | RG_rl_79_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_79_en )
		RG_rl_79 <= RG_rl_79_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_92 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_80_t1 = TR_92 ;
	7'h01 :
		RG_rl_80_t1 = TR_92 ;
	7'h02 :
		RG_rl_80_t1 = TR_92 ;
	7'h03 :
		RG_rl_80_t1 = TR_92 ;
	7'h04 :
		RG_rl_80_t1 = TR_92 ;
	7'h05 :
		RG_rl_80_t1 = TR_92 ;
	7'h06 :
		RG_rl_80_t1 = TR_92 ;
	7'h07 :
		RG_rl_80_t1 = TR_92 ;
	7'h08 :
		RG_rl_80_t1 = TR_92 ;
	7'h09 :
		RG_rl_80_t1 = TR_92 ;
	7'h0a :
		RG_rl_80_t1 = TR_92 ;
	7'h0b :
		RG_rl_80_t1 = TR_92 ;
	7'h0c :
		RG_rl_80_t1 = TR_92 ;
	7'h0d :
		RG_rl_80_t1 = TR_92 ;
	7'h0e :
		RG_rl_80_t1 = TR_92 ;
	7'h0f :
		RG_rl_80_t1 = TR_92 ;
	7'h10 :
		RG_rl_80_t1 = TR_92 ;
	7'h11 :
		RG_rl_80_t1 = TR_92 ;
	7'h12 :
		RG_rl_80_t1 = TR_92 ;
	7'h13 :
		RG_rl_80_t1 = TR_92 ;
	7'h14 :
		RG_rl_80_t1 = TR_92 ;
	7'h15 :
		RG_rl_80_t1 = TR_92 ;
	7'h16 :
		RG_rl_80_t1 = TR_92 ;
	7'h17 :
		RG_rl_80_t1 = TR_92 ;
	7'h18 :
		RG_rl_80_t1 = TR_92 ;
	7'h19 :
		RG_rl_80_t1 = TR_92 ;
	7'h1a :
		RG_rl_80_t1 = TR_92 ;
	7'h1b :
		RG_rl_80_t1 = TR_92 ;
	7'h1c :
		RG_rl_80_t1 = TR_92 ;
	7'h1d :
		RG_rl_80_t1 = TR_92 ;
	7'h1e :
		RG_rl_80_t1 = TR_92 ;
	7'h1f :
		RG_rl_80_t1 = TR_92 ;
	7'h20 :
		RG_rl_80_t1 = TR_92 ;
	7'h21 :
		RG_rl_80_t1 = TR_92 ;
	7'h22 :
		RG_rl_80_t1 = TR_92 ;
	7'h23 :
		RG_rl_80_t1 = TR_92 ;
	7'h24 :
		RG_rl_80_t1 = TR_92 ;
	7'h25 :
		RG_rl_80_t1 = TR_92 ;
	7'h26 :
		RG_rl_80_t1 = TR_92 ;
	7'h27 :
		RG_rl_80_t1 = TR_92 ;
	7'h28 :
		RG_rl_80_t1 = TR_92 ;
	7'h29 :
		RG_rl_80_t1 = TR_92 ;
	7'h2a :
		RG_rl_80_t1 = TR_92 ;
	7'h2b :
		RG_rl_80_t1 = TR_92 ;
	7'h2c :
		RG_rl_80_t1 = TR_92 ;
	7'h2d :
		RG_rl_80_t1 = TR_92 ;
	7'h2e :
		RG_rl_80_t1 = TR_92 ;
	7'h2f :
		RG_rl_80_t1 = TR_92 ;
	7'h30 :
		RG_rl_80_t1 = TR_92 ;
	7'h31 :
		RG_rl_80_t1 = TR_92 ;
	7'h32 :
		RG_rl_80_t1 = TR_92 ;
	7'h33 :
		RG_rl_80_t1 = TR_92 ;
	7'h34 :
		RG_rl_80_t1 = TR_92 ;
	7'h35 :
		RG_rl_80_t1 = TR_92 ;
	7'h36 :
		RG_rl_80_t1 = TR_92 ;
	7'h37 :
		RG_rl_80_t1 = TR_92 ;
	7'h38 :
		RG_rl_80_t1 = TR_92 ;
	7'h39 :
		RG_rl_80_t1 = TR_92 ;
	7'h3a :
		RG_rl_80_t1 = TR_92 ;
	7'h3b :
		RG_rl_80_t1 = TR_92 ;
	7'h3c :
		RG_rl_80_t1 = TR_92 ;
	7'h3d :
		RG_rl_80_t1 = TR_92 ;
	7'h3e :
		RG_rl_80_t1 = TR_92 ;
	7'h3f :
		RG_rl_80_t1 = TR_92 ;
	7'h40 :
		RG_rl_80_t1 = TR_92 ;
	7'h41 :
		RG_rl_80_t1 = TR_92 ;
	7'h42 :
		RG_rl_80_t1 = TR_92 ;
	7'h43 :
		RG_rl_80_t1 = TR_92 ;
	7'h44 :
		RG_rl_80_t1 = TR_92 ;
	7'h45 :
		RG_rl_80_t1 = TR_92 ;
	7'h46 :
		RG_rl_80_t1 = TR_92 ;
	7'h47 :
		RG_rl_80_t1 = TR_92 ;
	7'h48 :
		RG_rl_80_t1 = TR_92 ;
	7'h49 :
		RG_rl_80_t1 = TR_92 ;
	7'h4a :
		RG_rl_80_t1 = TR_92 ;
	7'h4b :
		RG_rl_80_t1 = TR_92 ;
	7'h4c :
		RG_rl_80_t1 = TR_92 ;
	7'h4d :
		RG_rl_80_t1 = TR_92 ;
	7'h4e :
		RG_rl_80_t1 = TR_92 ;
	7'h4f :
		RG_rl_80_t1 = TR_92 ;
	7'h50 :
		RG_rl_80_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h51 :
		RG_rl_80_t1 = TR_92 ;
	7'h52 :
		RG_rl_80_t1 = TR_92 ;
	7'h53 :
		RG_rl_80_t1 = TR_92 ;
	7'h54 :
		RG_rl_80_t1 = TR_92 ;
	7'h55 :
		RG_rl_80_t1 = TR_92 ;
	7'h56 :
		RG_rl_80_t1 = TR_92 ;
	7'h57 :
		RG_rl_80_t1 = TR_92 ;
	7'h58 :
		RG_rl_80_t1 = TR_92 ;
	7'h59 :
		RG_rl_80_t1 = TR_92 ;
	7'h5a :
		RG_rl_80_t1 = TR_92 ;
	7'h5b :
		RG_rl_80_t1 = TR_92 ;
	7'h5c :
		RG_rl_80_t1 = TR_92 ;
	7'h5d :
		RG_rl_80_t1 = TR_92 ;
	7'h5e :
		RG_rl_80_t1 = TR_92 ;
	7'h5f :
		RG_rl_80_t1 = TR_92 ;
	7'h60 :
		RG_rl_80_t1 = TR_92 ;
	7'h61 :
		RG_rl_80_t1 = TR_92 ;
	7'h62 :
		RG_rl_80_t1 = TR_92 ;
	7'h63 :
		RG_rl_80_t1 = TR_92 ;
	7'h64 :
		RG_rl_80_t1 = TR_92 ;
	7'h65 :
		RG_rl_80_t1 = TR_92 ;
	7'h66 :
		RG_rl_80_t1 = TR_92 ;
	7'h67 :
		RG_rl_80_t1 = TR_92 ;
	7'h68 :
		RG_rl_80_t1 = TR_92 ;
	7'h69 :
		RG_rl_80_t1 = TR_92 ;
	7'h6a :
		RG_rl_80_t1 = TR_92 ;
	7'h6b :
		RG_rl_80_t1 = TR_92 ;
	7'h6c :
		RG_rl_80_t1 = TR_92 ;
	7'h6d :
		RG_rl_80_t1 = TR_92 ;
	7'h6e :
		RG_rl_80_t1 = TR_92 ;
	7'h6f :
		RG_rl_80_t1 = TR_92 ;
	7'h70 :
		RG_rl_80_t1 = TR_92 ;
	7'h71 :
		RG_rl_80_t1 = TR_92 ;
	7'h72 :
		RG_rl_80_t1 = TR_92 ;
	7'h73 :
		RG_rl_80_t1 = TR_92 ;
	7'h74 :
		RG_rl_80_t1 = TR_92 ;
	7'h75 :
		RG_rl_80_t1 = TR_92 ;
	7'h76 :
		RG_rl_80_t1 = TR_92 ;
	7'h77 :
		RG_rl_80_t1 = TR_92 ;
	7'h78 :
		RG_rl_80_t1 = TR_92 ;
	7'h79 :
		RG_rl_80_t1 = TR_92 ;
	7'h7a :
		RG_rl_80_t1 = TR_92 ;
	7'h7b :
		RG_rl_80_t1 = TR_92 ;
	7'h7c :
		RG_rl_80_t1 = TR_92 ;
	7'h7d :
		RG_rl_80_t1 = TR_92 ;
	7'h7e :
		RG_rl_80_t1 = TR_92 ;
	7'h7f :
		RG_rl_80_t1 = TR_92 ;
	default :
		RG_rl_80_t1 = 9'hx ;
	endcase
always @ ( RG_rl_80_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_21 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_80_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h50 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_80_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_21 )
		| ( { 9{ U_569 } } & RG_rl_80_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_80_en = ( U_570 | RG_rl_80_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_80_en )
		RG_rl_80 <= RG_rl_80_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_93 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_81_t1 = TR_93 ;
	7'h01 :
		RG_rl_81_t1 = TR_93 ;
	7'h02 :
		RG_rl_81_t1 = TR_93 ;
	7'h03 :
		RG_rl_81_t1 = TR_93 ;
	7'h04 :
		RG_rl_81_t1 = TR_93 ;
	7'h05 :
		RG_rl_81_t1 = TR_93 ;
	7'h06 :
		RG_rl_81_t1 = TR_93 ;
	7'h07 :
		RG_rl_81_t1 = TR_93 ;
	7'h08 :
		RG_rl_81_t1 = TR_93 ;
	7'h09 :
		RG_rl_81_t1 = TR_93 ;
	7'h0a :
		RG_rl_81_t1 = TR_93 ;
	7'h0b :
		RG_rl_81_t1 = TR_93 ;
	7'h0c :
		RG_rl_81_t1 = TR_93 ;
	7'h0d :
		RG_rl_81_t1 = TR_93 ;
	7'h0e :
		RG_rl_81_t1 = TR_93 ;
	7'h0f :
		RG_rl_81_t1 = TR_93 ;
	7'h10 :
		RG_rl_81_t1 = TR_93 ;
	7'h11 :
		RG_rl_81_t1 = TR_93 ;
	7'h12 :
		RG_rl_81_t1 = TR_93 ;
	7'h13 :
		RG_rl_81_t1 = TR_93 ;
	7'h14 :
		RG_rl_81_t1 = TR_93 ;
	7'h15 :
		RG_rl_81_t1 = TR_93 ;
	7'h16 :
		RG_rl_81_t1 = TR_93 ;
	7'h17 :
		RG_rl_81_t1 = TR_93 ;
	7'h18 :
		RG_rl_81_t1 = TR_93 ;
	7'h19 :
		RG_rl_81_t1 = TR_93 ;
	7'h1a :
		RG_rl_81_t1 = TR_93 ;
	7'h1b :
		RG_rl_81_t1 = TR_93 ;
	7'h1c :
		RG_rl_81_t1 = TR_93 ;
	7'h1d :
		RG_rl_81_t1 = TR_93 ;
	7'h1e :
		RG_rl_81_t1 = TR_93 ;
	7'h1f :
		RG_rl_81_t1 = TR_93 ;
	7'h20 :
		RG_rl_81_t1 = TR_93 ;
	7'h21 :
		RG_rl_81_t1 = TR_93 ;
	7'h22 :
		RG_rl_81_t1 = TR_93 ;
	7'h23 :
		RG_rl_81_t1 = TR_93 ;
	7'h24 :
		RG_rl_81_t1 = TR_93 ;
	7'h25 :
		RG_rl_81_t1 = TR_93 ;
	7'h26 :
		RG_rl_81_t1 = TR_93 ;
	7'h27 :
		RG_rl_81_t1 = TR_93 ;
	7'h28 :
		RG_rl_81_t1 = TR_93 ;
	7'h29 :
		RG_rl_81_t1 = TR_93 ;
	7'h2a :
		RG_rl_81_t1 = TR_93 ;
	7'h2b :
		RG_rl_81_t1 = TR_93 ;
	7'h2c :
		RG_rl_81_t1 = TR_93 ;
	7'h2d :
		RG_rl_81_t1 = TR_93 ;
	7'h2e :
		RG_rl_81_t1 = TR_93 ;
	7'h2f :
		RG_rl_81_t1 = TR_93 ;
	7'h30 :
		RG_rl_81_t1 = TR_93 ;
	7'h31 :
		RG_rl_81_t1 = TR_93 ;
	7'h32 :
		RG_rl_81_t1 = TR_93 ;
	7'h33 :
		RG_rl_81_t1 = TR_93 ;
	7'h34 :
		RG_rl_81_t1 = TR_93 ;
	7'h35 :
		RG_rl_81_t1 = TR_93 ;
	7'h36 :
		RG_rl_81_t1 = TR_93 ;
	7'h37 :
		RG_rl_81_t1 = TR_93 ;
	7'h38 :
		RG_rl_81_t1 = TR_93 ;
	7'h39 :
		RG_rl_81_t1 = TR_93 ;
	7'h3a :
		RG_rl_81_t1 = TR_93 ;
	7'h3b :
		RG_rl_81_t1 = TR_93 ;
	7'h3c :
		RG_rl_81_t1 = TR_93 ;
	7'h3d :
		RG_rl_81_t1 = TR_93 ;
	7'h3e :
		RG_rl_81_t1 = TR_93 ;
	7'h3f :
		RG_rl_81_t1 = TR_93 ;
	7'h40 :
		RG_rl_81_t1 = TR_93 ;
	7'h41 :
		RG_rl_81_t1 = TR_93 ;
	7'h42 :
		RG_rl_81_t1 = TR_93 ;
	7'h43 :
		RG_rl_81_t1 = TR_93 ;
	7'h44 :
		RG_rl_81_t1 = TR_93 ;
	7'h45 :
		RG_rl_81_t1 = TR_93 ;
	7'h46 :
		RG_rl_81_t1 = TR_93 ;
	7'h47 :
		RG_rl_81_t1 = TR_93 ;
	7'h48 :
		RG_rl_81_t1 = TR_93 ;
	7'h49 :
		RG_rl_81_t1 = TR_93 ;
	7'h4a :
		RG_rl_81_t1 = TR_93 ;
	7'h4b :
		RG_rl_81_t1 = TR_93 ;
	7'h4c :
		RG_rl_81_t1 = TR_93 ;
	7'h4d :
		RG_rl_81_t1 = TR_93 ;
	7'h4e :
		RG_rl_81_t1 = TR_93 ;
	7'h4f :
		RG_rl_81_t1 = TR_93 ;
	7'h50 :
		RG_rl_81_t1 = TR_93 ;
	7'h51 :
		RG_rl_81_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h52 :
		RG_rl_81_t1 = TR_93 ;
	7'h53 :
		RG_rl_81_t1 = TR_93 ;
	7'h54 :
		RG_rl_81_t1 = TR_93 ;
	7'h55 :
		RG_rl_81_t1 = TR_93 ;
	7'h56 :
		RG_rl_81_t1 = TR_93 ;
	7'h57 :
		RG_rl_81_t1 = TR_93 ;
	7'h58 :
		RG_rl_81_t1 = TR_93 ;
	7'h59 :
		RG_rl_81_t1 = TR_93 ;
	7'h5a :
		RG_rl_81_t1 = TR_93 ;
	7'h5b :
		RG_rl_81_t1 = TR_93 ;
	7'h5c :
		RG_rl_81_t1 = TR_93 ;
	7'h5d :
		RG_rl_81_t1 = TR_93 ;
	7'h5e :
		RG_rl_81_t1 = TR_93 ;
	7'h5f :
		RG_rl_81_t1 = TR_93 ;
	7'h60 :
		RG_rl_81_t1 = TR_93 ;
	7'h61 :
		RG_rl_81_t1 = TR_93 ;
	7'h62 :
		RG_rl_81_t1 = TR_93 ;
	7'h63 :
		RG_rl_81_t1 = TR_93 ;
	7'h64 :
		RG_rl_81_t1 = TR_93 ;
	7'h65 :
		RG_rl_81_t1 = TR_93 ;
	7'h66 :
		RG_rl_81_t1 = TR_93 ;
	7'h67 :
		RG_rl_81_t1 = TR_93 ;
	7'h68 :
		RG_rl_81_t1 = TR_93 ;
	7'h69 :
		RG_rl_81_t1 = TR_93 ;
	7'h6a :
		RG_rl_81_t1 = TR_93 ;
	7'h6b :
		RG_rl_81_t1 = TR_93 ;
	7'h6c :
		RG_rl_81_t1 = TR_93 ;
	7'h6d :
		RG_rl_81_t1 = TR_93 ;
	7'h6e :
		RG_rl_81_t1 = TR_93 ;
	7'h6f :
		RG_rl_81_t1 = TR_93 ;
	7'h70 :
		RG_rl_81_t1 = TR_93 ;
	7'h71 :
		RG_rl_81_t1 = TR_93 ;
	7'h72 :
		RG_rl_81_t1 = TR_93 ;
	7'h73 :
		RG_rl_81_t1 = TR_93 ;
	7'h74 :
		RG_rl_81_t1 = TR_93 ;
	7'h75 :
		RG_rl_81_t1 = TR_93 ;
	7'h76 :
		RG_rl_81_t1 = TR_93 ;
	7'h77 :
		RG_rl_81_t1 = TR_93 ;
	7'h78 :
		RG_rl_81_t1 = TR_93 ;
	7'h79 :
		RG_rl_81_t1 = TR_93 ;
	7'h7a :
		RG_rl_81_t1 = TR_93 ;
	7'h7b :
		RG_rl_81_t1 = TR_93 ;
	7'h7c :
		RG_rl_81_t1 = TR_93 ;
	7'h7d :
		RG_rl_81_t1 = TR_93 ;
	7'h7e :
		RG_rl_81_t1 = TR_93 ;
	7'h7f :
		RG_rl_81_t1 = TR_93 ;
	default :
		RG_rl_81_t1 = 9'hx ;
	endcase
always @ ( RG_rl_81_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_22 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_81_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h51 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_81_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_22 )
		| ( { 9{ U_569 } } & RG_rl_81_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_81_en = ( U_570 | RG_rl_81_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_81_en )
		RG_rl_81 <= RG_rl_81_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_94 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_82_t1 = TR_94 ;
	7'h01 :
		RG_rl_82_t1 = TR_94 ;
	7'h02 :
		RG_rl_82_t1 = TR_94 ;
	7'h03 :
		RG_rl_82_t1 = TR_94 ;
	7'h04 :
		RG_rl_82_t1 = TR_94 ;
	7'h05 :
		RG_rl_82_t1 = TR_94 ;
	7'h06 :
		RG_rl_82_t1 = TR_94 ;
	7'h07 :
		RG_rl_82_t1 = TR_94 ;
	7'h08 :
		RG_rl_82_t1 = TR_94 ;
	7'h09 :
		RG_rl_82_t1 = TR_94 ;
	7'h0a :
		RG_rl_82_t1 = TR_94 ;
	7'h0b :
		RG_rl_82_t1 = TR_94 ;
	7'h0c :
		RG_rl_82_t1 = TR_94 ;
	7'h0d :
		RG_rl_82_t1 = TR_94 ;
	7'h0e :
		RG_rl_82_t1 = TR_94 ;
	7'h0f :
		RG_rl_82_t1 = TR_94 ;
	7'h10 :
		RG_rl_82_t1 = TR_94 ;
	7'h11 :
		RG_rl_82_t1 = TR_94 ;
	7'h12 :
		RG_rl_82_t1 = TR_94 ;
	7'h13 :
		RG_rl_82_t1 = TR_94 ;
	7'h14 :
		RG_rl_82_t1 = TR_94 ;
	7'h15 :
		RG_rl_82_t1 = TR_94 ;
	7'h16 :
		RG_rl_82_t1 = TR_94 ;
	7'h17 :
		RG_rl_82_t1 = TR_94 ;
	7'h18 :
		RG_rl_82_t1 = TR_94 ;
	7'h19 :
		RG_rl_82_t1 = TR_94 ;
	7'h1a :
		RG_rl_82_t1 = TR_94 ;
	7'h1b :
		RG_rl_82_t1 = TR_94 ;
	7'h1c :
		RG_rl_82_t1 = TR_94 ;
	7'h1d :
		RG_rl_82_t1 = TR_94 ;
	7'h1e :
		RG_rl_82_t1 = TR_94 ;
	7'h1f :
		RG_rl_82_t1 = TR_94 ;
	7'h20 :
		RG_rl_82_t1 = TR_94 ;
	7'h21 :
		RG_rl_82_t1 = TR_94 ;
	7'h22 :
		RG_rl_82_t1 = TR_94 ;
	7'h23 :
		RG_rl_82_t1 = TR_94 ;
	7'h24 :
		RG_rl_82_t1 = TR_94 ;
	7'h25 :
		RG_rl_82_t1 = TR_94 ;
	7'h26 :
		RG_rl_82_t1 = TR_94 ;
	7'h27 :
		RG_rl_82_t1 = TR_94 ;
	7'h28 :
		RG_rl_82_t1 = TR_94 ;
	7'h29 :
		RG_rl_82_t1 = TR_94 ;
	7'h2a :
		RG_rl_82_t1 = TR_94 ;
	7'h2b :
		RG_rl_82_t1 = TR_94 ;
	7'h2c :
		RG_rl_82_t1 = TR_94 ;
	7'h2d :
		RG_rl_82_t1 = TR_94 ;
	7'h2e :
		RG_rl_82_t1 = TR_94 ;
	7'h2f :
		RG_rl_82_t1 = TR_94 ;
	7'h30 :
		RG_rl_82_t1 = TR_94 ;
	7'h31 :
		RG_rl_82_t1 = TR_94 ;
	7'h32 :
		RG_rl_82_t1 = TR_94 ;
	7'h33 :
		RG_rl_82_t1 = TR_94 ;
	7'h34 :
		RG_rl_82_t1 = TR_94 ;
	7'h35 :
		RG_rl_82_t1 = TR_94 ;
	7'h36 :
		RG_rl_82_t1 = TR_94 ;
	7'h37 :
		RG_rl_82_t1 = TR_94 ;
	7'h38 :
		RG_rl_82_t1 = TR_94 ;
	7'h39 :
		RG_rl_82_t1 = TR_94 ;
	7'h3a :
		RG_rl_82_t1 = TR_94 ;
	7'h3b :
		RG_rl_82_t1 = TR_94 ;
	7'h3c :
		RG_rl_82_t1 = TR_94 ;
	7'h3d :
		RG_rl_82_t1 = TR_94 ;
	7'h3e :
		RG_rl_82_t1 = TR_94 ;
	7'h3f :
		RG_rl_82_t1 = TR_94 ;
	7'h40 :
		RG_rl_82_t1 = TR_94 ;
	7'h41 :
		RG_rl_82_t1 = TR_94 ;
	7'h42 :
		RG_rl_82_t1 = TR_94 ;
	7'h43 :
		RG_rl_82_t1 = TR_94 ;
	7'h44 :
		RG_rl_82_t1 = TR_94 ;
	7'h45 :
		RG_rl_82_t1 = TR_94 ;
	7'h46 :
		RG_rl_82_t1 = TR_94 ;
	7'h47 :
		RG_rl_82_t1 = TR_94 ;
	7'h48 :
		RG_rl_82_t1 = TR_94 ;
	7'h49 :
		RG_rl_82_t1 = TR_94 ;
	7'h4a :
		RG_rl_82_t1 = TR_94 ;
	7'h4b :
		RG_rl_82_t1 = TR_94 ;
	7'h4c :
		RG_rl_82_t1 = TR_94 ;
	7'h4d :
		RG_rl_82_t1 = TR_94 ;
	7'h4e :
		RG_rl_82_t1 = TR_94 ;
	7'h4f :
		RG_rl_82_t1 = TR_94 ;
	7'h50 :
		RG_rl_82_t1 = TR_94 ;
	7'h51 :
		RG_rl_82_t1 = TR_94 ;
	7'h52 :
		RG_rl_82_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h53 :
		RG_rl_82_t1 = TR_94 ;
	7'h54 :
		RG_rl_82_t1 = TR_94 ;
	7'h55 :
		RG_rl_82_t1 = TR_94 ;
	7'h56 :
		RG_rl_82_t1 = TR_94 ;
	7'h57 :
		RG_rl_82_t1 = TR_94 ;
	7'h58 :
		RG_rl_82_t1 = TR_94 ;
	7'h59 :
		RG_rl_82_t1 = TR_94 ;
	7'h5a :
		RG_rl_82_t1 = TR_94 ;
	7'h5b :
		RG_rl_82_t1 = TR_94 ;
	7'h5c :
		RG_rl_82_t1 = TR_94 ;
	7'h5d :
		RG_rl_82_t1 = TR_94 ;
	7'h5e :
		RG_rl_82_t1 = TR_94 ;
	7'h5f :
		RG_rl_82_t1 = TR_94 ;
	7'h60 :
		RG_rl_82_t1 = TR_94 ;
	7'h61 :
		RG_rl_82_t1 = TR_94 ;
	7'h62 :
		RG_rl_82_t1 = TR_94 ;
	7'h63 :
		RG_rl_82_t1 = TR_94 ;
	7'h64 :
		RG_rl_82_t1 = TR_94 ;
	7'h65 :
		RG_rl_82_t1 = TR_94 ;
	7'h66 :
		RG_rl_82_t1 = TR_94 ;
	7'h67 :
		RG_rl_82_t1 = TR_94 ;
	7'h68 :
		RG_rl_82_t1 = TR_94 ;
	7'h69 :
		RG_rl_82_t1 = TR_94 ;
	7'h6a :
		RG_rl_82_t1 = TR_94 ;
	7'h6b :
		RG_rl_82_t1 = TR_94 ;
	7'h6c :
		RG_rl_82_t1 = TR_94 ;
	7'h6d :
		RG_rl_82_t1 = TR_94 ;
	7'h6e :
		RG_rl_82_t1 = TR_94 ;
	7'h6f :
		RG_rl_82_t1 = TR_94 ;
	7'h70 :
		RG_rl_82_t1 = TR_94 ;
	7'h71 :
		RG_rl_82_t1 = TR_94 ;
	7'h72 :
		RG_rl_82_t1 = TR_94 ;
	7'h73 :
		RG_rl_82_t1 = TR_94 ;
	7'h74 :
		RG_rl_82_t1 = TR_94 ;
	7'h75 :
		RG_rl_82_t1 = TR_94 ;
	7'h76 :
		RG_rl_82_t1 = TR_94 ;
	7'h77 :
		RG_rl_82_t1 = TR_94 ;
	7'h78 :
		RG_rl_82_t1 = TR_94 ;
	7'h79 :
		RG_rl_82_t1 = TR_94 ;
	7'h7a :
		RG_rl_82_t1 = TR_94 ;
	7'h7b :
		RG_rl_82_t1 = TR_94 ;
	7'h7c :
		RG_rl_82_t1 = TR_94 ;
	7'h7d :
		RG_rl_82_t1 = TR_94 ;
	7'h7e :
		RG_rl_82_t1 = TR_94 ;
	7'h7f :
		RG_rl_82_t1 = TR_94 ;
	default :
		RG_rl_82_t1 = 9'hx ;
	endcase
always @ ( RG_rl_82_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_23 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_82_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h52 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_82_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_23 )
		| ( { 9{ U_569 } } & RG_rl_82_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_82_en = ( U_570 | RG_rl_82_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_82_en )
		RG_rl_82 <= RG_rl_82_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_95 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_83_t1 = TR_95 ;
	7'h01 :
		RG_rl_83_t1 = TR_95 ;
	7'h02 :
		RG_rl_83_t1 = TR_95 ;
	7'h03 :
		RG_rl_83_t1 = TR_95 ;
	7'h04 :
		RG_rl_83_t1 = TR_95 ;
	7'h05 :
		RG_rl_83_t1 = TR_95 ;
	7'h06 :
		RG_rl_83_t1 = TR_95 ;
	7'h07 :
		RG_rl_83_t1 = TR_95 ;
	7'h08 :
		RG_rl_83_t1 = TR_95 ;
	7'h09 :
		RG_rl_83_t1 = TR_95 ;
	7'h0a :
		RG_rl_83_t1 = TR_95 ;
	7'h0b :
		RG_rl_83_t1 = TR_95 ;
	7'h0c :
		RG_rl_83_t1 = TR_95 ;
	7'h0d :
		RG_rl_83_t1 = TR_95 ;
	7'h0e :
		RG_rl_83_t1 = TR_95 ;
	7'h0f :
		RG_rl_83_t1 = TR_95 ;
	7'h10 :
		RG_rl_83_t1 = TR_95 ;
	7'h11 :
		RG_rl_83_t1 = TR_95 ;
	7'h12 :
		RG_rl_83_t1 = TR_95 ;
	7'h13 :
		RG_rl_83_t1 = TR_95 ;
	7'h14 :
		RG_rl_83_t1 = TR_95 ;
	7'h15 :
		RG_rl_83_t1 = TR_95 ;
	7'h16 :
		RG_rl_83_t1 = TR_95 ;
	7'h17 :
		RG_rl_83_t1 = TR_95 ;
	7'h18 :
		RG_rl_83_t1 = TR_95 ;
	7'h19 :
		RG_rl_83_t1 = TR_95 ;
	7'h1a :
		RG_rl_83_t1 = TR_95 ;
	7'h1b :
		RG_rl_83_t1 = TR_95 ;
	7'h1c :
		RG_rl_83_t1 = TR_95 ;
	7'h1d :
		RG_rl_83_t1 = TR_95 ;
	7'h1e :
		RG_rl_83_t1 = TR_95 ;
	7'h1f :
		RG_rl_83_t1 = TR_95 ;
	7'h20 :
		RG_rl_83_t1 = TR_95 ;
	7'h21 :
		RG_rl_83_t1 = TR_95 ;
	7'h22 :
		RG_rl_83_t1 = TR_95 ;
	7'h23 :
		RG_rl_83_t1 = TR_95 ;
	7'h24 :
		RG_rl_83_t1 = TR_95 ;
	7'h25 :
		RG_rl_83_t1 = TR_95 ;
	7'h26 :
		RG_rl_83_t1 = TR_95 ;
	7'h27 :
		RG_rl_83_t1 = TR_95 ;
	7'h28 :
		RG_rl_83_t1 = TR_95 ;
	7'h29 :
		RG_rl_83_t1 = TR_95 ;
	7'h2a :
		RG_rl_83_t1 = TR_95 ;
	7'h2b :
		RG_rl_83_t1 = TR_95 ;
	7'h2c :
		RG_rl_83_t1 = TR_95 ;
	7'h2d :
		RG_rl_83_t1 = TR_95 ;
	7'h2e :
		RG_rl_83_t1 = TR_95 ;
	7'h2f :
		RG_rl_83_t1 = TR_95 ;
	7'h30 :
		RG_rl_83_t1 = TR_95 ;
	7'h31 :
		RG_rl_83_t1 = TR_95 ;
	7'h32 :
		RG_rl_83_t1 = TR_95 ;
	7'h33 :
		RG_rl_83_t1 = TR_95 ;
	7'h34 :
		RG_rl_83_t1 = TR_95 ;
	7'h35 :
		RG_rl_83_t1 = TR_95 ;
	7'h36 :
		RG_rl_83_t1 = TR_95 ;
	7'h37 :
		RG_rl_83_t1 = TR_95 ;
	7'h38 :
		RG_rl_83_t1 = TR_95 ;
	7'h39 :
		RG_rl_83_t1 = TR_95 ;
	7'h3a :
		RG_rl_83_t1 = TR_95 ;
	7'h3b :
		RG_rl_83_t1 = TR_95 ;
	7'h3c :
		RG_rl_83_t1 = TR_95 ;
	7'h3d :
		RG_rl_83_t1 = TR_95 ;
	7'h3e :
		RG_rl_83_t1 = TR_95 ;
	7'h3f :
		RG_rl_83_t1 = TR_95 ;
	7'h40 :
		RG_rl_83_t1 = TR_95 ;
	7'h41 :
		RG_rl_83_t1 = TR_95 ;
	7'h42 :
		RG_rl_83_t1 = TR_95 ;
	7'h43 :
		RG_rl_83_t1 = TR_95 ;
	7'h44 :
		RG_rl_83_t1 = TR_95 ;
	7'h45 :
		RG_rl_83_t1 = TR_95 ;
	7'h46 :
		RG_rl_83_t1 = TR_95 ;
	7'h47 :
		RG_rl_83_t1 = TR_95 ;
	7'h48 :
		RG_rl_83_t1 = TR_95 ;
	7'h49 :
		RG_rl_83_t1 = TR_95 ;
	7'h4a :
		RG_rl_83_t1 = TR_95 ;
	7'h4b :
		RG_rl_83_t1 = TR_95 ;
	7'h4c :
		RG_rl_83_t1 = TR_95 ;
	7'h4d :
		RG_rl_83_t1 = TR_95 ;
	7'h4e :
		RG_rl_83_t1 = TR_95 ;
	7'h4f :
		RG_rl_83_t1 = TR_95 ;
	7'h50 :
		RG_rl_83_t1 = TR_95 ;
	7'h51 :
		RG_rl_83_t1 = TR_95 ;
	7'h52 :
		RG_rl_83_t1 = TR_95 ;
	7'h53 :
		RG_rl_83_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h54 :
		RG_rl_83_t1 = TR_95 ;
	7'h55 :
		RG_rl_83_t1 = TR_95 ;
	7'h56 :
		RG_rl_83_t1 = TR_95 ;
	7'h57 :
		RG_rl_83_t1 = TR_95 ;
	7'h58 :
		RG_rl_83_t1 = TR_95 ;
	7'h59 :
		RG_rl_83_t1 = TR_95 ;
	7'h5a :
		RG_rl_83_t1 = TR_95 ;
	7'h5b :
		RG_rl_83_t1 = TR_95 ;
	7'h5c :
		RG_rl_83_t1 = TR_95 ;
	7'h5d :
		RG_rl_83_t1 = TR_95 ;
	7'h5e :
		RG_rl_83_t1 = TR_95 ;
	7'h5f :
		RG_rl_83_t1 = TR_95 ;
	7'h60 :
		RG_rl_83_t1 = TR_95 ;
	7'h61 :
		RG_rl_83_t1 = TR_95 ;
	7'h62 :
		RG_rl_83_t1 = TR_95 ;
	7'h63 :
		RG_rl_83_t1 = TR_95 ;
	7'h64 :
		RG_rl_83_t1 = TR_95 ;
	7'h65 :
		RG_rl_83_t1 = TR_95 ;
	7'h66 :
		RG_rl_83_t1 = TR_95 ;
	7'h67 :
		RG_rl_83_t1 = TR_95 ;
	7'h68 :
		RG_rl_83_t1 = TR_95 ;
	7'h69 :
		RG_rl_83_t1 = TR_95 ;
	7'h6a :
		RG_rl_83_t1 = TR_95 ;
	7'h6b :
		RG_rl_83_t1 = TR_95 ;
	7'h6c :
		RG_rl_83_t1 = TR_95 ;
	7'h6d :
		RG_rl_83_t1 = TR_95 ;
	7'h6e :
		RG_rl_83_t1 = TR_95 ;
	7'h6f :
		RG_rl_83_t1 = TR_95 ;
	7'h70 :
		RG_rl_83_t1 = TR_95 ;
	7'h71 :
		RG_rl_83_t1 = TR_95 ;
	7'h72 :
		RG_rl_83_t1 = TR_95 ;
	7'h73 :
		RG_rl_83_t1 = TR_95 ;
	7'h74 :
		RG_rl_83_t1 = TR_95 ;
	7'h75 :
		RG_rl_83_t1 = TR_95 ;
	7'h76 :
		RG_rl_83_t1 = TR_95 ;
	7'h77 :
		RG_rl_83_t1 = TR_95 ;
	7'h78 :
		RG_rl_83_t1 = TR_95 ;
	7'h79 :
		RG_rl_83_t1 = TR_95 ;
	7'h7a :
		RG_rl_83_t1 = TR_95 ;
	7'h7b :
		RG_rl_83_t1 = TR_95 ;
	7'h7c :
		RG_rl_83_t1 = TR_95 ;
	7'h7d :
		RG_rl_83_t1 = TR_95 ;
	7'h7e :
		RG_rl_83_t1 = TR_95 ;
	7'h7f :
		RG_rl_83_t1 = TR_95 ;
	default :
		RG_rl_83_t1 = 9'hx ;
	endcase
always @ ( RG_rl_83_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_24 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_83_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h53 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_83_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_24 )
		| ( { 9{ U_569 } } & RG_rl_83_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_83_en = ( U_570 | RG_rl_83_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_83_en )
		RG_rl_83 <= RG_rl_83_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_96 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_84_t1 = TR_96 ;
	7'h01 :
		RG_rl_84_t1 = TR_96 ;
	7'h02 :
		RG_rl_84_t1 = TR_96 ;
	7'h03 :
		RG_rl_84_t1 = TR_96 ;
	7'h04 :
		RG_rl_84_t1 = TR_96 ;
	7'h05 :
		RG_rl_84_t1 = TR_96 ;
	7'h06 :
		RG_rl_84_t1 = TR_96 ;
	7'h07 :
		RG_rl_84_t1 = TR_96 ;
	7'h08 :
		RG_rl_84_t1 = TR_96 ;
	7'h09 :
		RG_rl_84_t1 = TR_96 ;
	7'h0a :
		RG_rl_84_t1 = TR_96 ;
	7'h0b :
		RG_rl_84_t1 = TR_96 ;
	7'h0c :
		RG_rl_84_t1 = TR_96 ;
	7'h0d :
		RG_rl_84_t1 = TR_96 ;
	7'h0e :
		RG_rl_84_t1 = TR_96 ;
	7'h0f :
		RG_rl_84_t1 = TR_96 ;
	7'h10 :
		RG_rl_84_t1 = TR_96 ;
	7'h11 :
		RG_rl_84_t1 = TR_96 ;
	7'h12 :
		RG_rl_84_t1 = TR_96 ;
	7'h13 :
		RG_rl_84_t1 = TR_96 ;
	7'h14 :
		RG_rl_84_t1 = TR_96 ;
	7'h15 :
		RG_rl_84_t1 = TR_96 ;
	7'h16 :
		RG_rl_84_t1 = TR_96 ;
	7'h17 :
		RG_rl_84_t1 = TR_96 ;
	7'h18 :
		RG_rl_84_t1 = TR_96 ;
	7'h19 :
		RG_rl_84_t1 = TR_96 ;
	7'h1a :
		RG_rl_84_t1 = TR_96 ;
	7'h1b :
		RG_rl_84_t1 = TR_96 ;
	7'h1c :
		RG_rl_84_t1 = TR_96 ;
	7'h1d :
		RG_rl_84_t1 = TR_96 ;
	7'h1e :
		RG_rl_84_t1 = TR_96 ;
	7'h1f :
		RG_rl_84_t1 = TR_96 ;
	7'h20 :
		RG_rl_84_t1 = TR_96 ;
	7'h21 :
		RG_rl_84_t1 = TR_96 ;
	7'h22 :
		RG_rl_84_t1 = TR_96 ;
	7'h23 :
		RG_rl_84_t1 = TR_96 ;
	7'h24 :
		RG_rl_84_t1 = TR_96 ;
	7'h25 :
		RG_rl_84_t1 = TR_96 ;
	7'h26 :
		RG_rl_84_t1 = TR_96 ;
	7'h27 :
		RG_rl_84_t1 = TR_96 ;
	7'h28 :
		RG_rl_84_t1 = TR_96 ;
	7'h29 :
		RG_rl_84_t1 = TR_96 ;
	7'h2a :
		RG_rl_84_t1 = TR_96 ;
	7'h2b :
		RG_rl_84_t1 = TR_96 ;
	7'h2c :
		RG_rl_84_t1 = TR_96 ;
	7'h2d :
		RG_rl_84_t1 = TR_96 ;
	7'h2e :
		RG_rl_84_t1 = TR_96 ;
	7'h2f :
		RG_rl_84_t1 = TR_96 ;
	7'h30 :
		RG_rl_84_t1 = TR_96 ;
	7'h31 :
		RG_rl_84_t1 = TR_96 ;
	7'h32 :
		RG_rl_84_t1 = TR_96 ;
	7'h33 :
		RG_rl_84_t1 = TR_96 ;
	7'h34 :
		RG_rl_84_t1 = TR_96 ;
	7'h35 :
		RG_rl_84_t1 = TR_96 ;
	7'h36 :
		RG_rl_84_t1 = TR_96 ;
	7'h37 :
		RG_rl_84_t1 = TR_96 ;
	7'h38 :
		RG_rl_84_t1 = TR_96 ;
	7'h39 :
		RG_rl_84_t1 = TR_96 ;
	7'h3a :
		RG_rl_84_t1 = TR_96 ;
	7'h3b :
		RG_rl_84_t1 = TR_96 ;
	7'h3c :
		RG_rl_84_t1 = TR_96 ;
	7'h3d :
		RG_rl_84_t1 = TR_96 ;
	7'h3e :
		RG_rl_84_t1 = TR_96 ;
	7'h3f :
		RG_rl_84_t1 = TR_96 ;
	7'h40 :
		RG_rl_84_t1 = TR_96 ;
	7'h41 :
		RG_rl_84_t1 = TR_96 ;
	7'h42 :
		RG_rl_84_t1 = TR_96 ;
	7'h43 :
		RG_rl_84_t1 = TR_96 ;
	7'h44 :
		RG_rl_84_t1 = TR_96 ;
	7'h45 :
		RG_rl_84_t1 = TR_96 ;
	7'h46 :
		RG_rl_84_t1 = TR_96 ;
	7'h47 :
		RG_rl_84_t1 = TR_96 ;
	7'h48 :
		RG_rl_84_t1 = TR_96 ;
	7'h49 :
		RG_rl_84_t1 = TR_96 ;
	7'h4a :
		RG_rl_84_t1 = TR_96 ;
	7'h4b :
		RG_rl_84_t1 = TR_96 ;
	7'h4c :
		RG_rl_84_t1 = TR_96 ;
	7'h4d :
		RG_rl_84_t1 = TR_96 ;
	7'h4e :
		RG_rl_84_t1 = TR_96 ;
	7'h4f :
		RG_rl_84_t1 = TR_96 ;
	7'h50 :
		RG_rl_84_t1 = TR_96 ;
	7'h51 :
		RG_rl_84_t1 = TR_96 ;
	7'h52 :
		RG_rl_84_t1 = TR_96 ;
	7'h53 :
		RG_rl_84_t1 = TR_96 ;
	7'h54 :
		RG_rl_84_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h55 :
		RG_rl_84_t1 = TR_96 ;
	7'h56 :
		RG_rl_84_t1 = TR_96 ;
	7'h57 :
		RG_rl_84_t1 = TR_96 ;
	7'h58 :
		RG_rl_84_t1 = TR_96 ;
	7'h59 :
		RG_rl_84_t1 = TR_96 ;
	7'h5a :
		RG_rl_84_t1 = TR_96 ;
	7'h5b :
		RG_rl_84_t1 = TR_96 ;
	7'h5c :
		RG_rl_84_t1 = TR_96 ;
	7'h5d :
		RG_rl_84_t1 = TR_96 ;
	7'h5e :
		RG_rl_84_t1 = TR_96 ;
	7'h5f :
		RG_rl_84_t1 = TR_96 ;
	7'h60 :
		RG_rl_84_t1 = TR_96 ;
	7'h61 :
		RG_rl_84_t1 = TR_96 ;
	7'h62 :
		RG_rl_84_t1 = TR_96 ;
	7'h63 :
		RG_rl_84_t1 = TR_96 ;
	7'h64 :
		RG_rl_84_t1 = TR_96 ;
	7'h65 :
		RG_rl_84_t1 = TR_96 ;
	7'h66 :
		RG_rl_84_t1 = TR_96 ;
	7'h67 :
		RG_rl_84_t1 = TR_96 ;
	7'h68 :
		RG_rl_84_t1 = TR_96 ;
	7'h69 :
		RG_rl_84_t1 = TR_96 ;
	7'h6a :
		RG_rl_84_t1 = TR_96 ;
	7'h6b :
		RG_rl_84_t1 = TR_96 ;
	7'h6c :
		RG_rl_84_t1 = TR_96 ;
	7'h6d :
		RG_rl_84_t1 = TR_96 ;
	7'h6e :
		RG_rl_84_t1 = TR_96 ;
	7'h6f :
		RG_rl_84_t1 = TR_96 ;
	7'h70 :
		RG_rl_84_t1 = TR_96 ;
	7'h71 :
		RG_rl_84_t1 = TR_96 ;
	7'h72 :
		RG_rl_84_t1 = TR_96 ;
	7'h73 :
		RG_rl_84_t1 = TR_96 ;
	7'h74 :
		RG_rl_84_t1 = TR_96 ;
	7'h75 :
		RG_rl_84_t1 = TR_96 ;
	7'h76 :
		RG_rl_84_t1 = TR_96 ;
	7'h77 :
		RG_rl_84_t1 = TR_96 ;
	7'h78 :
		RG_rl_84_t1 = TR_96 ;
	7'h79 :
		RG_rl_84_t1 = TR_96 ;
	7'h7a :
		RG_rl_84_t1 = TR_96 ;
	7'h7b :
		RG_rl_84_t1 = TR_96 ;
	7'h7c :
		RG_rl_84_t1 = TR_96 ;
	7'h7d :
		RG_rl_84_t1 = TR_96 ;
	7'h7e :
		RG_rl_84_t1 = TR_96 ;
	7'h7f :
		RG_rl_84_t1 = TR_96 ;
	default :
		RG_rl_84_t1 = 9'hx ;
	endcase
always @ ( RG_rl_84_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_25 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_84_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h54 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_84_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_25 )
		| ( { 9{ U_569 } } & RG_rl_84_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_84_en = ( U_570 | RG_rl_84_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_84_en )
		RG_rl_84 <= RG_rl_84_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_97 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_85_t1 = TR_97 ;
	7'h01 :
		RG_rl_85_t1 = TR_97 ;
	7'h02 :
		RG_rl_85_t1 = TR_97 ;
	7'h03 :
		RG_rl_85_t1 = TR_97 ;
	7'h04 :
		RG_rl_85_t1 = TR_97 ;
	7'h05 :
		RG_rl_85_t1 = TR_97 ;
	7'h06 :
		RG_rl_85_t1 = TR_97 ;
	7'h07 :
		RG_rl_85_t1 = TR_97 ;
	7'h08 :
		RG_rl_85_t1 = TR_97 ;
	7'h09 :
		RG_rl_85_t1 = TR_97 ;
	7'h0a :
		RG_rl_85_t1 = TR_97 ;
	7'h0b :
		RG_rl_85_t1 = TR_97 ;
	7'h0c :
		RG_rl_85_t1 = TR_97 ;
	7'h0d :
		RG_rl_85_t1 = TR_97 ;
	7'h0e :
		RG_rl_85_t1 = TR_97 ;
	7'h0f :
		RG_rl_85_t1 = TR_97 ;
	7'h10 :
		RG_rl_85_t1 = TR_97 ;
	7'h11 :
		RG_rl_85_t1 = TR_97 ;
	7'h12 :
		RG_rl_85_t1 = TR_97 ;
	7'h13 :
		RG_rl_85_t1 = TR_97 ;
	7'h14 :
		RG_rl_85_t1 = TR_97 ;
	7'h15 :
		RG_rl_85_t1 = TR_97 ;
	7'h16 :
		RG_rl_85_t1 = TR_97 ;
	7'h17 :
		RG_rl_85_t1 = TR_97 ;
	7'h18 :
		RG_rl_85_t1 = TR_97 ;
	7'h19 :
		RG_rl_85_t1 = TR_97 ;
	7'h1a :
		RG_rl_85_t1 = TR_97 ;
	7'h1b :
		RG_rl_85_t1 = TR_97 ;
	7'h1c :
		RG_rl_85_t1 = TR_97 ;
	7'h1d :
		RG_rl_85_t1 = TR_97 ;
	7'h1e :
		RG_rl_85_t1 = TR_97 ;
	7'h1f :
		RG_rl_85_t1 = TR_97 ;
	7'h20 :
		RG_rl_85_t1 = TR_97 ;
	7'h21 :
		RG_rl_85_t1 = TR_97 ;
	7'h22 :
		RG_rl_85_t1 = TR_97 ;
	7'h23 :
		RG_rl_85_t1 = TR_97 ;
	7'h24 :
		RG_rl_85_t1 = TR_97 ;
	7'h25 :
		RG_rl_85_t1 = TR_97 ;
	7'h26 :
		RG_rl_85_t1 = TR_97 ;
	7'h27 :
		RG_rl_85_t1 = TR_97 ;
	7'h28 :
		RG_rl_85_t1 = TR_97 ;
	7'h29 :
		RG_rl_85_t1 = TR_97 ;
	7'h2a :
		RG_rl_85_t1 = TR_97 ;
	7'h2b :
		RG_rl_85_t1 = TR_97 ;
	7'h2c :
		RG_rl_85_t1 = TR_97 ;
	7'h2d :
		RG_rl_85_t1 = TR_97 ;
	7'h2e :
		RG_rl_85_t1 = TR_97 ;
	7'h2f :
		RG_rl_85_t1 = TR_97 ;
	7'h30 :
		RG_rl_85_t1 = TR_97 ;
	7'h31 :
		RG_rl_85_t1 = TR_97 ;
	7'h32 :
		RG_rl_85_t1 = TR_97 ;
	7'h33 :
		RG_rl_85_t1 = TR_97 ;
	7'h34 :
		RG_rl_85_t1 = TR_97 ;
	7'h35 :
		RG_rl_85_t1 = TR_97 ;
	7'h36 :
		RG_rl_85_t1 = TR_97 ;
	7'h37 :
		RG_rl_85_t1 = TR_97 ;
	7'h38 :
		RG_rl_85_t1 = TR_97 ;
	7'h39 :
		RG_rl_85_t1 = TR_97 ;
	7'h3a :
		RG_rl_85_t1 = TR_97 ;
	7'h3b :
		RG_rl_85_t1 = TR_97 ;
	7'h3c :
		RG_rl_85_t1 = TR_97 ;
	7'h3d :
		RG_rl_85_t1 = TR_97 ;
	7'h3e :
		RG_rl_85_t1 = TR_97 ;
	7'h3f :
		RG_rl_85_t1 = TR_97 ;
	7'h40 :
		RG_rl_85_t1 = TR_97 ;
	7'h41 :
		RG_rl_85_t1 = TR_97 ;
	7'h42 :
		RG_rl_85_t1 = TR_97 ;
	7'h43 :
		RG_rl_85_t1 = TR_97 ;
	7'h44 :
		RG_rl_85_t1 = TR_97 ;
	7'h45 :
		RG_rl_85_t1 = TR_97 ;
	7'h46 :
		RG_rl_85_t1 = TR_97 ;
	7'h47 :
		RG_rl_85_t1 = TR_97 ;
	7'h48 :
		RG_rl_85_t1 = TR_97 ;
	7'h49 :
		RG_rl_85_t1 = TR_97 ;
	7'h4a :
		RG_rl_85_t1 = TR_97 ;
	7'h4b :
		RG_rl_85_t1 = TR_97 ;
	7'h4c :
		RG_rl_85_t1 = TR_97 ;
	7'h4d :
		RG_rl_85_t1 = TR_97 ;
	7'h4e :
		RG_rl_85_t1 = TR_97 ;
	7'h4f :
		RG_rl_85_t1 = TR_97 ;
	7'h50 :
		RG_rl_85_t1 = TR_97 ;
	7'h51 :
		RG_rl_85_t1 = TR_97 ;
	7'h52 :
		RG_rl_85_t1 = TR_97 ;
	7'h53 :
		RG_rl_85_t1 = TR_97 ;
	7'h54 :
		RG_rl_85_t1 = TR_97 ;
	7'h55 :
		RG_rl_85_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h56 :
		RG_rl_85_t1 = TR_97 ;
	7'h57 :
		RG_rl_85_t1 = TR_97 ;
	7'h58 :
		RG_rl_85_t1 = TR_97 ;
	7'h59 :
		RG_rl_85_t1 = TR_97 ;
	7'h5a :
		RG_rl_85_t1 = TR_97 ;
	7'h5b :
		RG_rl_85_t1 = TR_97 ;
	7'h5c :
		RG_rl_85_t1 = TR_97 ;
	7'h5d :
		RG_rl_85_t1 = TR_97 ;
	7'h5e :
		RG_rl_85_t1 = TR_97 ;
	7'h5f :
		RG_rl_85_t1 = TR_97 ;
	7'h60 :
		RG_rl_85_t1 = TR_97 ;
	7'h61 :
		RG_rl_85_t1 = TR_97 ;
	7'h62 :
		RG_rl_85_t1 = TR_97 ;
	7'h63 :
		RG_rl_85_t1 = TR_97 ;
	7'h64 :
		RG_rl_85_t1 = TR_97 ;
	7'h65 :
		RG_rl_85_t1 = TR_97 ;
	7'h66 :
		RG_rl_85_t1 = TR_97 ;
	7'h67 :
		RG_rl_85_t1 = TR_97 ;
	7'h68 :
		RG_rl_85_t1 = TR_97 ;
	7'h69 :
		RG_rl_85_t1 = TR_97 ;
	7'h6a :
		RG_rl_85_t1 = TR_97 ;
	7'h6b :
		RG_rl_85_t1 = TR_97 ;
	7'h6c :
		RG_rl_85_t1 = TR_97 ;
	7'h6d :
		RG_rl_85_t1 = TR_97 ;
	7'h6e :
		RG_rl_85_t1 = TR_97 ;
	7'h6f :
		RG_rl_85_t1 = TR_97 ;
	7'h70 :
		RG_rl_85_t1 = TR_97 ;
	7'h71 :
		RG_rl_85_t1 = TR_97 ;
	7'h72 :
		RG_rl_85_t1 = TR_97 ;
	7'h73 :
		RG_rl_85_t1 = TR_97 ;
	7'h74 :
		RG_rl_85_t1 = TR_97 ;
	7'h75 :
		RG_rl_85_t1 = TR_97 ;
	7'h76 :
		RG_rl_85_t1 = TR_97 ;
	7'h77 :
		RG_rl_85_t1 = TR_97 ;
	7'h78 :
		RG_rl_85_t1 = TR_97 ;
	7'h79 :
		RG_rl_85_t1 = TR_97 ;
	7'h7a :
		RG_rl_85_t1 = TR_97 ;
	7'h7b :
		RG_rl_85_t1 = TR_97 ;
	7'h7c :
		RG_rl_85_t1 = TR_97 ;
	7'h7d :
		RG_rl_85_t1 = TR_97 ;
	7'h7e :
		RG_rl_85_t1 = TR_97 ;
	7'h7f :
		RG_rl_85_t1 = TR_97 ;
	default :
		RG_rl_85_t1 = 9'hx ;
	endcase
always @ ( RG_rl_85_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_26 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_85_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h55 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_85_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_26 )
		| ( { 9{ U_569 } } & RG_rl_85_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_85_en = ( U_570 | RG_rl_85_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_85_en )
		RG_rl_85 <= RG_rl_85_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_98 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_86_t1 = TR_98 ;
	7'h01 :
		RG_rl_86_t1 = TR_98 ;
	7'h02 :
		RG_rl_86_t1 = TR_98 ;
	7'h03 :
		RG_rl_86_t1 = TR_98 ;
	7'h04 :
		RG_rl_86_t1 = TR_98 ;
	7'h05 :
		RG_rl_86_t1 = TR_98 ;
	7'h06 :
		RG_rl_86_t1 = TR_98 ;
	7'h07 :
		RG_rl_86_t1 = TR_98 ;
	7'h08 :
		RG_rl_86_t1 = TR_98 ;
	7'h09 :
		RG_rl_86_t1 = TR_98 ;
	7'h0a :
		RG_rl_86_t1 = TR_98 ;
	7'h0b :
		RG_rl_86_t1 = TR_98 ;
	7'h0c :
		RG_rl_86_t1 = TR_98 ;
	7'h0d :
		RG_rl_86_t1 = TR_98 ;
	7'h0e :
		RG_rl_86_t1 = TR_98 ;
	7'h0f :
		RG_rl_86_t1 = TR_98 ;
	7'h10 :
		RG_rl_86_t1 = TR_98 ;
	7'h11 :
		RG_rl_86_t1 = TR_98 ;
	7'h12 :
		RG_rl_86_t1 = TR_98 ;
	7'h13 :
		RG_rl_86_t1 = TR_98 ;
	7'h14 :
		RG_rl_86_t1 = TR_98 ;
	7'h15 :
		RG_rl_86_t1 = TR_98 ;
	7'h16 :
		RG_rl_86_t1 = TR_98 ;
	7'h17 :
		RG_rl_86_t1 = TR_98 ;
	7'h18 :
		RG_rl_86_t1 = TR_98 ;
	7'h19 :
		RG_rl_86_t1 = TR_98 ;
	7'h1a :
		RG_rl_86_t1 = TR_98 ;
	7'h1b :
		RG_rl_86_t1 = TR_98 ;
	7'h1c :
		RG_rl_86_t1 = TR_98 ;
	7'h1d :
		RG_rl_86_t1 = TR_98 ;
	7'h1e :
		RG_rl_86_t1 = TR_98 ;
	7'h1f :
		RG_rl_86_t1 = TR_98 ;
	7'h20 :
		RG_rl_86_t1 = TR_98 ;
	7'h21 :
		RG_rl_86_t1 = TR_98 ;
	7'h22 :
		RG_rl_86_t1 = TR_98 ;
	7'h23 :
		RG_rl_86_t1 = TR_98 ;
	7'h24 :
		RG_rl_86_t1 = TR_98 ;
	7'h25 :
		RG_rl_86_t1 = TR_98 ;
	7'h26 :
		RG_rl_86_t1 = TR_98 ;
	7'h27 :
		RG_rl_86_t1 = TR_98 ;
	7'h28 :
		RG_rl_86_t1 = TR_98 ;
	7'h29 :
		RG_rl_86_t1 = TR_98 ;
	7'h2a :
		RG_rl_86_t1 = TR_98 ;
	7'h2b :
		RG_rl_86_t1 = TR_98 ;
	7'h2c :
		RG_rl_86_t1 = TR_98 ;
	7'h2d :
		RG_rl_86_t1 = TR_98 ;
	7'h2e :
		RG_rl_86_t1 = TR_98 ;
	7'h2f :
		RG_rl_86_t1 = TR_98 ;
	7'h30 :
		RG_rl_86_t1 = TR_98 ;
	7'h31 :
		RG_rl_86_t1 = TR_98 ;
	7'h32 :
		RG_rl_86_t1 = TR_98 ;
	7'h33 :
		RG_rl_86_t1 = TR_98 ;
	7'h34 :
		RG_rl_86_t1 = TR_98 ;
	7'h35 :
		RG_rl_86_t1 = TR_98 ;
	7'h36 :
		RG_rl_86_t1 = TR_98 ;
	7'h37 :
		RG_rl_86_t1 = TR_98 ;
	7'h38 :
		RG_rl_86_t1 = TR_98 ;
	7'h39 :
		RG_rl_86_t1 = TR_98 ;
	7'h3a :
		RG_rl_86_t1 = TR_98 ;
	7'h3b :
		RG_rl_86_t1 = TR_98 ;
	7'h3c :
		RG_rl_86_t1 = TR_98 ;
	7'h3d :
		RG_rl_86_t1 = TR_98 ;
	7'h3e :
		RG_rl_86_t1 = TR_98 ;
	7'h3f :
		RG_rl_86_t1 = TR_98 ;
	7'h40 :
		RG_rl_86_t1 = TR_98 ;
	7'h41 :
		RG_rl_86_t1 = TR_98 ;
	7'h42 :
		RG_rl_86_t1 = TR_98 ;
	7'h43 :
		RG_rl_86_t1 = TR_98 ;
	7'h44 :
		RG_rl_86_t1 = TR_98 ;
	7'h45 :
		RG_rl_86_t1 = TR_98 ;
	7'h46 :
		RG_rl_86_t1 = TR_98 ;
	7'h47 :
		RG_rl_86_t1 = TR_98 ;
	7'h48 :
		RG_rl_86_t1 = TR_98 ;
	7'h49 :
		RG_rl_86_t1 = TR_98 ;
	7'h4a :
		RG_rl_86_t1 = TR_98 ;
	7'h4b :
		RG_rl_86_t1 = TR_98 ;
	7'h4c :
		RG_rl_86_t1 = TR_98 ;
	7'h4d :
		RG_rl_86_t1 = TR_98 ;
	7'h4e :
		RG_rl_86_t1 = TR_98 ;
	7'h4f :
		RG_rl_86_t1 = TR_98 ;
	7'h50 :
		RG_rl_86_t1 = TR_98 ;
	7'h51 :
		RG_rl_86_t1 = TR_98 ;
	7'h52 :
		RG_rl_86_t1 = TR_98 ;
	7'h53 :
		RG_rl_86_t1 = TR_98 ;
	7'h54 :
		RG_rl_86_t1 = TR_98 ;
	7'h55 :
		RG_rl_86_t1 = TR_98 ;
	7'h56 :
		RG_rl_86_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h57 :
		RG_rl_86_t1 = TR_98 ;
	7'h58 :
		RG_rl_86_t1 = TR_98 ;
	7'h59 :
		RG_rl_86_t1 = TR_98 ;
	7'h5a :
		RG_rl_86_t1 = TR_98 ;
	7'h5b :
		RG_rl_86_t1 = TR_98 ;
	7'h5c :
		RG_rl_86_t1 = TR_98 ;
	7'h5d :
		RG_rl_86_t1 = TR_98 ;
	7'h5e :
		RG_rl_86_t1 = TR_98 ;
	7'h5f :
		RG_rl_86_t1 = TR_98 ;
	7'h60 :
		RG_rl_86_t1 = TR_98 ;
	7'h61 :
		RG_rl_86_t1 = TR_98 ;
	7'h62 :
		RG_rl_86_t1 = TR_98 ;
	7'h63 :
		RG_rl_86_t1 = TR_98 ;
	7'h64 :
		RG_rl_86_t1 = TR_98 ;
	7'h65 :
		RG_rl_86_t1 = TR_98 ;
	7'h66 :
		RG_rl_86_t1 = TR_98 ;
	7'h67 :
		RG_rl_86_t1 = TR_98 ;
	7'h68 :
		RG_rl_86_t1 = TR_98 ;
	7'h69 :
		RG_rl_86_t1 = TR_98 ;
	7'h6a :
		RG_rl_86_t1 = TR_98 ;
	7'h6b :
		RG_rl_86_t1 = TR_98 ;
	7'h6c :
		RG_rl_86_t1 = TR_98 ;
	7'h6d :
		RG_rl_86_t1 = TR_98 ;
	7'h6e :
		RG_rl_86_t1 = TR_98 ;
	7'h6f :
		RG_rl_86_t1 = TR_98 ;
	7'h70 :
		RG_rl_86_t1 = TR_98 ;
	7'h71 :
		RG_rl_86_t1 = TR_98 ;
	7'h72 :
		RG_rl_86_t1 = TR_98 ;
	7'h73 :
		RG_rl_86_t1 = TR_98 ;
	7'h74 :
		RG_rl_86_t1 = TR_98 ;
	7'h75 :
		RG_rl_86_t1 = TR_98 ;
	7'h76 :
		RG_rl_86_t1 = TR_98 ;
	7'h77 :
		RG_rl_86_t1 = TR_98 ;
	7'h78 :
		RG_rl_86_t1 = TR_98 ;
	7'h79 :
		RG_rl_86_t1 = TR_98 ;
	7'h7a :
		RG_rl_86_t1 = TR_98 ;
	7'h7b :
		RG_rl_86_t1 = TR_98 ;
	7'h7c :
		RG_rl_86_t1 = TR_98 ;
	7'h7d :
		RG_rl_86_t1 = TR_98 ;
	7'h7e :
		RG_rl_86_t1 = TR_98 ;
	7'h7f :
		RG_rl_86_t1 = TR_98 ;
	default :
		RG_rl_86_t1 = 9'hx ;
	endcase
always @ ( RG_rl_86_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_27 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_86_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h56 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_86_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_27 )
		| ( { 9{ U_569 } } & RG_rl_86_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_86_en = ( U_570 | RG_rl_86_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_86_en )
		RG_rl_86 <= RG_rl_86_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_99 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_87_t1 = TR_99 ;
	7'h01 :
		RG_rl_87_t1 = TR_99 ;
	7'h02 :
		RG_rl_87_t1 = TR_99 ;
	7'h03 :
		RG_rl_87_t1 = TR_99 ;
	7'h04 :
		RG_rl_87_t1 = TR_99 ;
	7'h05 :
		RG_rl_87_t1 = TR_99 ;
	7'h06 :
		RG_rl_87_t1 = TR_99 ;
	7'h07 :
		RG_rl_87_t1 = TR_99 ;
	7'h08 :
		RG_rl_87_t1 = TR_99 ;
	7'h09 :
		RG_rl_87_t1 = TR_99 ;
	7'h0a :
		RG_rl_87_t1 = TR_99 ;
	7'h0b :
		RG_rl_87_t1 = TR_99 ;
	7'h0c :
		RG_rl_87_t1 = TR_99 ;
	7'h0d :
		RG_rl_87_t1 = TR_99 ;
	7'h0e :
		RG_rl_87_t1 = TR_99 ;
	7'h0f :
		RG_rl_87_t1 = TR_99 ;
	7'h10 :
		RG_rl_87_t1 = TR_99 ;
	7'h11 :
		RG_rl_87_t1 = TR_99 ;
	7'h12 :
		RG_rl_87_t1 = TR_99 ;
	7'h13 :
		RG_rl_87_t1 = TR_99 ;
	7'h14 :
		RG_rl_87_t1 = TR_99 ;
	7'h15 :
		RG_rl_87_t1 = TR_99 ;
	7'h16 :
		RG_rl_87_t1 = TR_99 ;
	7'h17 :
		RG_rl_87_t1 = TR_99 ;
	7'h18 :
		RG_rl_87_t1 = TR_99 ;
	7'h19 :
		RG_rl_87_t1 = TR_99 ;
	7'h1a :
		RG_rl_87_t1 = TR_99 ;
	7'h1b :
		RG_rl_87_t1 = TR_99 ;
	7'h1c :
		RG_rl_87_t1 = TR_99 ;
	7'h1d :
		RG_rl_87_t1 = TR_99 ;
	7'h1e :
		RG_rl_87_t1 = TR_99 ;
	7'h1f :
		RG_rl_87_t1 = TR_99 ;
	7'h20 :
		RG_rl_87_t1 = TR_99 ;
	7'h21 :
		RG_rl_87_t1 = TR_99 ;
	7'h22 :
		RG_rl_87_t1 = TR_99 ;
	7'h23 :
		RG_rl_87_t1 = TR_99 ;
	7'h24 :
		RG_rl_87_t1 = TR_99 ;
	7'h25 :
		RG_rl_87_t1 = TR_99 ;
	7'h26 :
		RG_rl_87_t1 = TR_99 ;
	7'h27 :
		RG_rl_87_t1 = TR_99 ;
	7'h28 :
		RG_rl_87_t1 = TR_99 ;
	7'h29 :
		RG_rl_87_t1 = TR_99 ;
	7'h2a :
		RG_rl_87_t1 = TR_99 ;
	7'h2b :
		RG_rl_87_t1 = TR_99 ;
	7'h2c :
		RG_rl_87_t1 = TR_99 ;
	7'h2d :
		RG_rl_87_t1 = TR_99 ;
	7'h2e :
		RG_rl_87_t1 = TR_99 ;
	7'h2f :
		RG_rl_87_t1 = TR_99 ;
	7'h30 :
		RG_rl_87_t1 = TR_99 ;
	7'h31 :
		RG_rl_87_t1 = TR_99 ;
	7'h32 :
		RG_rl_87_t1 = TR_99 ;
	7'h33 :
		RG_rl_87_t1 = TR_99 ;
	7'h34 :
		RG_rl_87_t1 = TR_99 ;
	7'h35 :
		RG_rl_87_t1 = TR_99 ;
	7'h36 :
		RG_rl_87_t1 = TR_99 ;
	7'h37 :
		RG_rl_87_t1 = TR_99 ;
	7'h38 :
		RG_rl_87_t1 = TR_99 ;
	7'h39 :
		RG_rl_87_t1 = TR_99 ;
	7'h3a :
		RG_rl_87_t1 = TR_99 ;
	7'h3b :
		RG_rl_87_t1 = TR_99 ;
	7'h3c :
		RG_rl_87_t1 = TR_99 ;
	7'h3d :
		RG_rl_87_t1 = TR_99 ;
	7'h3e :
		RG_rl_87_t1 = TR_99 ;
	7'h3f :
		RG_rl_87_t1 = TR_99 ;
	7'h40 :
		RG_rl_87_t1 = TR_99 ;
	7'h41 :
		RG_rl_87_t1 = TR_99 ;
	7'h42 :
		RG_rl_87_t1 = TR_99 ;
	7'h43 :
		RG_rl_87_t1 = TR_99 ;
	7'h44 :
		RG_rl_87_t1 = TR_99 ;
	7'h45 :
		RG_rl_87_t1 = TR_99 ;
	7'h46 :
		RG_rl_87_t1 = TR_99 ;
	7'h47 :
		RG_rl_87_t1 = TR_99 ;
	7'h48 :
		RG_rl_87_t1 = TR_99 ;
	7'h49 :
		RG_rl_87_t1 = TR_99 ;
	7'h4a :
		RG_rl_87_t1 = TR_99 ;
	7'h4b :
		RG_rl_87_t1 = TR_99 ;
	7'h4c :
		RG_rl_87_t1 = TR_99 ;
	7'h4d :
		RG_rl_87_t1 = TR_99 ;
	7'h4e :
		RG_rl_87_t1 = TR_99 ;
	7'h4f :
		RG_rl_87_t1 = TR_99 ;
	7'h50 :
		RG_rl_87_t1 = TR_99 ;
	7'h51 :
		RG_rl_87_t1 = TR_99 ;
	7'h52 :
		RG_rl_87_t1 = TR_99 ;
	7'h53 :
		RG_rl_87_t1 = TR_99 ;
	7'h54 :
		RG_rl_87_t1 = TR_99 ;
	7'h55 :
		RG_rl_87_t1 = TR_99 ;
	7'h56 :
		RG_rl_87_t1 = TR_99 ;
	7'h57 :
		RG_rl_87_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h58 :
		RG_rl_87_t1 = TR_99 ;
	7'h59 :
		RG_rl_87_t1 = TR_99 ;
	7'h5a :
		RG_rl_87_t1 = TR_99 ;
	7'h5b :
		RG_rl_87_t1 = TR_99 ;
	7'h5c :
		RG_rl_87_t1 = TR_99 ;
	7'h5d :
		RG_rl_87_t1 = TR_99 ;
	7'h5e :
		RG_rl_87_t1 = TR_99 ;
	7'h5f :
		RG_rl_87_t1 = TR_99 ;
	7'h60 :
		RG_rl_87_t1 = TR_99 ;
	7'h61 :
		RG_rl_87_t1 = TR_99 ;
	7'h62 :
		RG_rl_87_t1 = TR_99 ;
	7'h63 :
		RG_rl_87_t1 = TR_99 ;
	7'h64 :
		RG_rl_87_t1 = TR_99 ;
	7'h65 :
		RG_rl_87_t1 = TR_99 ;
	7'h66 :
		RG_rl_87_t1 = TR_99 ;
	7'h67 :
		RG_rl_87_t1 = TR_99 ;
	7'h68 :
		RG_rl_87_t1 = TR_99 ;
	7'h69 :
		RG_rl_87_t1 = TR_99 ;
	7'h6a :
		RG_rl_87_t1 = TR_99 ;
	7'h6b :
		RG_rl_87_t1 = TR_99 ;
	7'h6c :
		RG_rl_87_t1 = TR_99 ;
	7'h6d :
		RG_rl_87_t1 = TR_99 ;
	7'h6e :
		RG_rl_87_t1 = TR_99 ;
	7'h6f :
		RG_rl_87_t1 = TR_99 ;
	7'h70 :
		RG_rl_87_t1 = TR_99 ;
	7'h71 :
		RG_rl_87_t1 = TR_99 ;
	7'h72 :
		RG_rl_87_t1 = TR_99 ;
	7'h73 :
		RG_rl_87_t1 = TR_99 ;
	7'h74 :
		RG_rl_87_t1 = TR_99 ;
	7'h75 :
		RG_rl_87_t1 = TR_99 ;
	7'h76 :
		RG_rl_87_t1 = TR_99 ;
	7'h77 :
		RG_rl_87_t1 = TR_99 ;
	7'h78 :
		RG_rl_87_t1 = TR_99 ;
	7'h79 :
		RG_rl_87_t1 = TR_99 ;
	7'h7a :
		RG_rl_87_t1 = TR_99 ;
	7'h7b :
		RG_rl_87_t1 = TR_99 ;
	7'h7c :
		RG_rl_87_t1 = TR_99 ;
	7'h7d :
		RG_rl_87_t1 = TR_99 ;
	7'h7e :
		RG_rl_87_t1 = TR_99 ;
	7'h7f :
		RG_rl_87_t1 = TR_99 ;
	default :
		RG_rl_87_t1 = 9'hx ;
	endcase
always @ ( RG_rl_87_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_28 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_87_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h57 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_87_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_28 )
		| ( { 9{ U_569 } } & RG_rl_87_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_87_en = ( U_570 | RG_rl_87_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_87_en )
		RG_rl_87 <= RG_rl_87_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_100 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_88_t1 = TR_100 ;
	7'h01 :
		RG_rl_88_t1 = TR_100 ;
	7'h02 :
		RG_rl_88_t1 = TR_100 ;
	7'h03 :
		RG_rl_88_t1 = TR_100 ;
	7'h04 :
		RG_rl_88_t1 = TR_100 ;
	7'h05 :
		RG_rl_88_t1 = TR_100 ;
	7'h06 :
		RG_rl_88_t1 = TR_100 ;
	7'h07 :
		RG_rl_88_t1 = TR_100 ;
	7'h08 :
		RG_rl_88_t1 = TR_100 ;
	7'h09 :
		RG_rl_88_t1 = TR_100 ;
	7'h0a :
		RG_rl_88_t1 = TR_100 ;
	7'h0b :
		RG_rl_88_t1 = TR_100 ;
	7'h0c :
		RG_rl_88_t1 = TR_100 ;
	7'h0d :
		RG_rl_88_t1 = TR_100 ;
	7'h0e :
		RG_rl_88_t1 = TR_100 ;
	7'h0f :
		RG_rl_88_t1 = TR_100 ;
	7'h10 :
		RG_rl_88_t1 = TR_100 ;
	7'h11 :
		RG_rl_88_t1 = TR_100 ;
	7'h12 :
		RG_rl_88_t1 = TR_100 ;
	7'h13 :
		RG_rl_88_t1 = TR_100 ;
	7'h14 :
		RG_rl_88_t1 = TR_100 ;
	7'h15 :
		RG_rl_88_t1 = TR_100 ;
	7'h16 :
		RG_rl_88_t1 = TR_100 ;
	7'h17 :
		RG_rl_88_t1 = TR_100 ;
	7'h18 :
		RG_rl_88_t1 = TR_100 ;
	7'h19 :
		RG_rl_88_t1 = TR_100 ;
	7'h1a :
		RG_rl_88_t1 = TR_100 ;
	7'h1b :
		RG_rl_88_t1 = TR_100 ;
	7'h1c :
		RG_rl_88_t1 = TR_100 ;
	7'h1d :
		RG_rl_88_t1 = TR_100 ;
	7'h1e :
		RG_rl_88_t1 = TR_100 ;
	7'h1f :
		RG_rl_88_t1 = TR_100 ;
	7'h20 :
		RG_rl_88_t1 = TR_100 ;
	7'h21 :
		RG_rl_88_t1 = TR_100 ;
	7'h22 :
		RG_rl_88_t1 = TR_100 ;
	7'h23 :
		RG_rl_88_t1 = TR_100 ;
	7'h24 :
		RG_rl_88_t1 = TR_100 ;
	7'h25 :
		RG_rl_88_t1 = TR_100 ;
	7'h26 :
		RG_rl_88_t1 = TR_100 ;
	7'h27 :
		RG_rl_88_t1 = TR_100 ;
	7'h28 :
		RG_rl_88_t1 = TR_100 ;
	7'h29 :
		RG_rl_88_t1 = TR_100 ;
	7'h2a :
		RG_rl_88_t1 = TR_100 ;
	7'h2b :
		RG_rl_88_t1 = TR_100 ;
	7'h2c :
		RG_rl_88_t1 = TR_100 ;
	7'h2d :
		RG_rl_88_t1 = TR_100 ;
	7'h2e :
		RG_rl_88_t1 = TR_100 ;
	7'h2f :
		RG_rl_88_t1 = TR_100 ;
	7'h30 :
		RG_rl_88_t1 = TR_100 ;
	7'h31 :
		RG_rl_88_t1 = TR_100 ;
	7'h32 :
		RG_rl_88_t1 = TR_100 ;
	7'h33 :
		RG_rl_88_t1 = TR_100 ;
	7'h34 :
		RG_rl_88_t1 = TR_100 ;
	7'h35 :
		RG_rl_88_t1 = TR_100 ;
	7'h36 :
		RG_rl_88_t1 = TR_100 ;
	7'h37 :
		RG_rl_88_t1 = TR_100 ;
	7'h38 :
		RG_rl_88_t1 = TR_100 ;
	7'h39 :
		RG_rl_88_t1 = TR_100 ;
	7'h3a :
		RG_rl_88_t1 = TR_100 ;
	7'h3b :
		RG_rl_88_t1 = TR_100 ;
	7'h3c :
		RG_rl_88_t1 = TR_100 ;
	7'h3d :
		RG_rl_88_t1 = TR_100 ;
	7'h3e :
		RG_rl_88_t1 = TR_100 ;
	7'h3f :
		RG_rl_88_t1 = TR_100 ;
	7'h40 :
		RG_rl_88_t1 = TR_100 ;
	7'h41 :
		RG_rl_88_t1 = TR_100 ;
	7'h42 :
		RG_rl_88_t1 = TR_100 ;
	7'h43 :
		RG_rl_88_t1 = TR_100 ;
	7'h44 :
		RG_rl_88_t1 = TR_100 ;
	7'h45 :
		RG_rl_88_t1 = TR_100 ;
	7'h46 :
		RG_rl_88_t1 = TR_100 ;
	7'h47 :
		RG_rl_88_t1 = TR_100 ;
	7'h48 :
		RG_rl_88_t1 = TR_100 ;
	7'h49 :
		RG_rl_88_t1 = TR_100 ;
	7'h4a :
		RG_rl_88_t1 = TR_100 ;
	7'h4b :
		RG_rl_88_t1 = TR_100 ;
	7'h4c :
		RG_rl_88_t1 = TR_100 ;
	7'h4d :
		RG_rl_88_t1 = TR_100 ;
	7'h4e :
		RG_rl_88_t1 = TR_100 ;
	7'h4f :
		RG_rl_88_t1 = TR_100 ;
	7'h50 :
		RG_rl_88_t1 = TR_100 ;
	7'h51 :
		RG_rl_88_t1 = TR_100 ;
	7'h52 :
		RG_rl_88_t1 = TR_100 ;
	7'h53 :
		RG_rl_88_t1 = TR_100 ;
	7'h54 :
		RG_rl_88_t1 = TR_100 ;
	7'h55 :
		RG_rl_88_t1 = TR_100 ;
	7'h56 :
		RG_rl_88_t1 = TR_100 ;
	7'h57 :
		RG_rl_88_t1 = TR_100 ;
	7'h58 :
		RG_rl_88_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h59 :
		RG_rl_88_t1 = TR_100 ;
	7'h5a :
		RG_rl_88_t1 = TR_100 ;
	7'h5b :
		RG_rl_88_t1 = TR_100 ;
	7'h5c :
		RG_rl_88_t1 = TR_100 ;
	7'h5d :
		RG_rl_88_t1 = TR_100 ;
	7'h5e :
		RG_rl_88_t1 = TR_100 ;
	7'h5f :
		RG_rl_88_t1 = TR_100 ;
	7'h60 :
		RG_rl_88_t1 = TR_100 ;
	7'h61 :
		RG_rl_88_t1 = TR_100 ;
	7'h62 :
		RG_rl_88_t1 = TR_100 ;
	7'h63 :
		RG_rl_88_t1 = TR_100 ;
	7'h64 :
		RG_rl_88_t1 = TR_100 ;
	7'h65 :
		RG_rl_88_t1 = TR_100 ;
	7'h66 :
		RG_rl_88_t1 = TR_100 ;
	7'h67 :
		RG_rl_88_t1 = TR_100 ;
	7'h68 :
		RG_rl_88_t1 = TR_100 ;
	7'h69 :
		RG_rl_88_t1 = TR_100 ;
	7'h6a :
		RG_rl_88_t1 = TR_100 ;
	7'h6b :
		RG_rl_88_t1 = TR_100 ;
	7'h6c :
		RG_rl_88_t1 = TR_100 ;
	7'h6d :
		RG_rl_88_t1 = TR_100 ;
	7'h6e :
		RG_rl_88_t1 = TR_100 ;
	7'h6f :
		RG_rl_88_t1 = TR_100 ;
	7'h70 :
		RG_rl_88_t1 = TR_100 ;
	7'h71 :
		RG_rl_88_t1 = TR_100 ;
	7'h72 :
		RG_rl_88_t1 = TR_100 ;
	7'h73 :
		RG_rl_88_t1 = TR_100 ;
	7'h74 :
		RG_rl_88_t1 = TR_100 ;
	7'h75 :
		RG_rl_88_t1 = TR_100 ;
	7'h76 :
		RG_rl_88_t1 = TR_100 ;
	7'h77 :
		RG_rl_88_t1 = TR_100 ;
	7'h78 :
		RG_rl_88_t1 = TR_100 ;
	7'h79 :
		RG_rl_88_t1 = TR_100 ;
	7'h7a :
		RG_rl_88_t1 = TR_100 ;
	7'h7b :
		RG_rl_88_t1 = TR_100 ;
	7'h7c :
		RG_rl_88_t1 = TR_100 ;
	7'h7d :
		RG_rl_88_t1 = TR_100 ;
	7'h7e :
		RG_rl_88_t1 = TR_100 ;
	7'h7f :
		RG_rl_88_t1 = TR_100 ;
	default :
		RG_rl_88_t1 = 9'hx ;
	endcase
always @ ( RG_rl_88_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_29 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_88_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h58 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_88_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_29 )
		| ( { 9{ U_569 } } & RG_rl_88_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_88_en = ( U_570 | RG_rl_88_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_88_en )
		RG_rl_88 <= RG_rl_88_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_101 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_89_t1 = TR_101 ;
	7'h01 :
		RG_rl_89_t1 = TR_101 ;
	7'h02 :
		RG_rl_89_t1 = TR_101 ;
	7'h03 :
		RG_rl_89_t1 = TR_101 ;
	7'h04 :
		RG_rl_89_t1 = TR_101 ;
	7'h05 :
		RG_rl_89_t1 = TR_101 ;
	7'h06 :
		RG_rl_89_t1 = TR_101 ;
	7'h07 :
		RG_rl_89_t1 = TR_101 ;
	7'h08 :
		RG_rl_89_t1 = TR_101 ;
	7'h09 :
		RG_rl_89_t1 = TR_101 ;
	7'h0a :
		RG_rl_89_t1 = TR_101 ;
	7'h0b :
		RG_rl_89_t1 = TR_101 ;
	7'h0c :
		RG_rl_89_t1 = TR_101 ;
	7'h0d :
		RG_rl_89_t1 = TR_101 ;
	7'h0e :
		RG_rl_89_t1 = TR_101 ;
	7'h0f :
		RG_rl_89_t1 = TR_101 ;
	7'h10 :
		RG_rl_89_t1 = TR_101 ;
	7'h11 :
		RG_rl_89_t1 = TR_101 ;
	7'h12 :
		RG_rl_89_t1 = TR_101 ;
	7'h13 :
		RG_rl_89_t1 = TR_101 ;
	7'h14 :
		RG_rl_89_t1 = TR_101 ;
	7'h15 :
		RG_rl_89_t1 = TR_101 ;
	7'h16 :
		RG_rl_89_t1 = TR_101 ;
	7'h17 :
		RG_rl_89_t1 = TR_101 ;
	7'h18 :
		RG_rl_89_t1 = TR_101 ;
	7'h19 :
		RG_rl_89_t1 = TR_101 ;
	7'h1a :
		RG_rl_89_t1 = TR_101 ;
	7'h1b :
		RG_rl_89_t1 = TR_101 ;
	7'h1c :
		RG_rl_89_t1 = TR_101 ;
	7'h1d :
		RG_rl_89_t1 = TR_101 ;
	7'h1e :
		RG_rl_89_t1 = TR_101 ;
	7'h1f :
		RG_rl_89_t1 = TR_101 ;
	7'h20 :
		RG_rl_89_t1 = TR_101 ;
	7'h21 :
		RG_rl_89_t1 = TR_101 ;
	7'h22 :
		RG_rl_89_t1 = TR_101 ;
	7'h23 :
		RG_rl_89_t1 = TR_101 ;
	7'h24 :
		RG_rl_89_t1 = TR_101 ;
	7'h25 :
		RG_rl_89_t1 = TR_101 ;
	7'h26 :
		RG_rl_89_t1 = TR_101 ;
	7'h27 :
		RG_rl_89_t1 = TR_101 ;
	7'h28 :
		RG_rl_89_t1 = TR_101 ;
	7'h29 :
		RG_rl_89_t1 = TR_101 ;
	7'h2a :
		RG_rl_89_t1 = TR_101 ;
	7'h2b :
		RG_rl_89_t1 = TR_101 ;
	7'h2c :
		RG_rl_89_t1 = TR_101 ;
	7'h2d :
		RG_rl_89_t1 = TR_101 ;
	7'h2e :
		RG_rl_89_t1 = TR_101 ;
	7'h2f :
		RG_rl_89_t1 = TR_101 ;
	7'h30 :
		RG_rl_89_t1 = TR_101 ;
	7'h31 :
		RG_rl_89_t1 = TR_101 ;
	7'h32 :
		RG_rl_89_t1 = TR_101 ;
	7'h33 :
		RG_rl_89_t1 = TR_101 ;
	7'h34 :
		RG_rl_89_t1 = TR_101 ;
	7'h35 :
		RG_rl_89_t1 = TR_101 ;
	7'h36 :
		RG_rl_89_t1 = TR_101 ;
	7'h37 :
		RG_rl_89_t1 = TR_101 ;
	7'h38 :
		RG_rl_89_t1 = TR_101 ;
	7'h39 :
		RG_rl_89_t1 = TR_101 ;
	7'h3a :
		RG_rl_89_t1 = TR_101 ;
	7'h3b :
		RG_rl_89_t1 = TR_101 ;
	7'h3c :
		RG_rl_89_t1 = TR_101 ;
	7'h3d :
		RG_rl_89_t1 = TR_101 ;
	7'h3e :
		RG_rl_89_t1 = TR_101 ;
	7'h3f :
		RG_rl_89_t1 = TR_101 ;
	7'h40 :
		RG_rl_89_t1 = TR_101 ;
	7'h41 :
		RG_rl_89_t1 = TR_101 ;
	7'h42 :
		RG_rl_89_t1 = TR_101 ;
	7'h43 :
		RG_rl_89_t1 = TR_101 ;
	7'h44 :
		RG_rl_89_t1 = TR_101 ;
	7'h45 :
		RG_rl_89_t1 = TR_101 ;
	7'h46 :
		RG_rl_89_t1 = TR_101 ;
	7'h47 :
		RG_rl_89_t1 = TR_101 ;
	7'h48 :
		RG_rl_89_t1 = TR_101 ;
	7'h49 :
		RG_rl_89_t1 = TR_101 ;
	7'h4a :
		RG_rl_89_t1 = TR_101 ;
	7'h4b :
		RG_rl_89_t1 = TR_101 ;
	7'h4c :
		RG_rl_89_t1 = TR_101 ;
	7'h4d :
		RG_rl_89_t1 = TR_101 ;
	7'h4e :
		RG_rl_89_t1 = TR_101 ;
	7'h4f :
		RG_rl_89_t1 = TR_101 ;
	7'h50 :
		RG_rl_89_t1 = TR_101 ;
	7'h51 :
		RG_rl_89_t1 = TR_101 ;
	7'h52 :
		RG_rl_89_t1 = TR_101 ;
	7'h53 :
		RG_rl_89_t1 = TR_101 ;
	7'h54 :
		RG_rl_89_t1 = TR_101 ;
	7'h55 :
		RG_rl_89_t1 = TR_101 ;
	7'h56 :
		RG_rl_89_t1 = TR_101 ;
	7'h57 :
		RG_rl_89_t1 = TR_101 ;
	7'h58 :
		RG_rl_89_t1 = TR_101 ;
	7'h59 :
		RG_rl_89_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5a :
		RG_rl_89_t1 = TR_101 ;
	7'h5b :
		RG_rl_89_t1 = TR_101 ;
	7'h5c :
		RG_rl_89_t1 = TR_101 ;
	7'h5d :
		RG_rl_89_t1 = TR_101 ;
	7'h5e :
		RG_rl_89_t1 = TR_101 ;
	7'h5f :
		RG_rl_89_t1 = TR_101 ;
	7'h60 :
		RG_rl_89_t1 = TR_101 ;
	7'h61 :
		RG_rl_89_t1 = TR_101 ;
	7'h62 :
		RG_rl_89_t1 = TR_101 ;
	7'h63 :
		RG_rl_89_t1 = TR_101 ;
	7'h64 :
		RG_rl_89_t1 = TR_101 ;
	7'h65 :
		RG_rl_89_t1 = TR_101 ;
	7'h66 :
		RG_rl_89_t1 = TR_101 ;
	7'h67 :
		RG_rl_89_t1 = TR_101 ;
	7'h68 :
		RG_rl_89_t1 = TR_101 ;
	7'h69 :
		RG_rl_89_t1 = TR_101 ;
	7'h6a :
		RG_rl_89_t1 = TR_101 ;
	7'h6b :
		RG_rl_89_t1 = TR_101 ;
	7'h6c :
		RG_rl_89_t1 = TR_101 ;
	7'h6d :
		RG_rl_89_t1 = TR_101 ;
	7'h6e :
		RG_rl_89_t1 = TR_101 ;
	7'h6f :
		RG_rl_89_t1 = TR_101 ;
	7'h70 :
		RG_rl_89_t1 = TR_101 ;
	7'h71 :
		RG_rl_89_t1 = TR_101 ;
	7'h72 :
		RG_rl_89_t1 = TR_101 ;
	7'h73 :
		RG_rl_89_t1 = TR_101 ;
	7'h74 :
		RG_rl_89_t1 = TR_101 ;
	7'h75 :
		RG_rl_89_t1 = TR_101 ;
	7'h76 :
		RG_rl_89_t1 = TR_101 ;
	7'h77 :
		RG_rl_89_t1 = TR_101 ;
	7'h78 :
		RG_rl_89_t1 = TR_101 ;
	7'h79 :
		RG_rl_89_t1 = TR_101 ;
	7'h7a :
		RG_rl_89_t1 = TR_101 ;
	7'h7b :
		RG_rl_89_t1 = TR_101 ;
	7'h7c :
		RG_rl_89_t1 = TR_101 ;
	7'h7d :
		RG_rl_89_t1 = TR_101 ;
	7'h7e :
		RG_rl_89_t1 = TR_101 ;
	7'h7f :
		RG_rl_89_t1 = TR_101 ;
	default :
		RG_rl_89_t1 = 9'hx ;
	endcase
always @ ( RG_rl_89_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_30 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_89_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h59 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_89_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_30 )
		| ( { 9{ U_569 } } & RG_rl_89_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_89_en = ( U_570 | RG_rl_89_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_89_en )
		RG_rl_89 <= RG_rl_89_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_102 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_90_t1 = TR_102 ;
	7'h01 :
		RG_rl_90_t1 = TR_102 ;
	7'h02 :
		RG_rl_90_t1 = TR_102 ;
	7'h03 :
		RG_rl_90_t1 = TR_102 ;
	7'h04 :
		RG_rl_90_t1 = TR_102 ;
	7'h05 :
		RG_rl_90_t1 = TR_102 ;
	7'h06 :
		RG_rl_90_t1 = TR_102 ;
	7'h07 :
		RG_rl_90_t1 = TR_102 ;
	7'h08 :
		RG_rl_90_t1 = TR_102 ;
	7'h09 :
		RG_rl_90_t1 = TR_102 ;
	7'h0a :
		RG_rl_90_t1 = TR_102 ;
	7'h0b :
		RG_rl_90_t1 = TR_102 ;
	7'h0c :
		RG_rl_90_t1 = TR_102 ;
	7'h0d :
		RG_rl_90_t1 = TR_102 ;
	7'h0e :
		RG_rl_90_t1 = TR_102 ;
	7'h0f :
		RG_rl_90_t1 = TR_102 ;
	7'h10 :
		RG_rl_90_t1 = TR_102 ;
	7'h11 :
		RG_rl_90_t1 = TR_102 ;
	7'h12 :
		RG_rl_90_t1 = TR_102 ;
	7'h13 :
		RG_rl_90_t1 = TR_102 ;
	7'h14 :
		RG_rl_90_t1 = TR_102 ;
	7'h15 :
		RG_rl_90_t1 = TR_102 ;
	7'h16 :
		RG_rl_90_t1 = TR_102 ;
	7'h17 :
		RG_rl_90_t1 = TR_102 ;
	7'h18 :
		RG_rl_90_t1 = TR_102 ;
	7'h19 :
		RG_rl_90_t1 = TR_102 ;
	7'h1a :
		RG_rl_90_t1 = TR_102 ;
	7'h1b :
		RG_rl_90_t1 = TR_102 ;
	7'h1c :
		RG_rl_90_t1 = TR_102 ;
	7'h1d :
		RG_rl_90_t1 = TR_102 ;
	7'h1e :
		RG_rl_90_t1 = TR_102 ;
	7'h1f :
		RG_rl_90_t1 = TR_102 ;
	7'h20 :
		RG_rl_90_t1 = TR_102 ;
	7'h21 :
		RG_rl_90_t1 = TR_102 ;
	7'h22 :
		RG_rl_90_t1 = TR_102 ;
	7'h23 :
		RG_rl_90_t1 = TR_102 ;
	7'h24 :
		RG_rl_90_t1 = TR_102 ;
	7'h25 :
		RG_rl_90_t1 = TR_102 ;
	7'h26 :
		RG_rl_90_t1 = TR_102 ;
	7'h27 :
		RG_rl_90_t1 = TR_102 ;
	7'h28 :
		RG_rl_90_t1 = TR_102 ;
	7'h29 :
		RG_rl_90_t1 = TR_102 ;
	7'h2a :
		RG_rl_90_t1 = TR_102 ;
	7'h2b :
		RG_rl_90_t1 = TR_102 ;
	7'h2c :
		RG_rl_90_t1 = TR_102 ;
	7'h2d :
		RG_rl_90_t1 = TR_102 ;
	7'h2e :
		RG_rl_90_t1 = TR_102 ;
	7'h2f :
		RG_rl_90_t1 = TR_102 ;
	7'h30 :
		RG_rl_90_t1 = TR_102 ;
	7'h31 :
		RG_rl_90_t1 = TR_102 ;
	7'h32 :
		RG_rl_90_t1 = TR_102 ;
	7'h33 :
		RG_rl_90_t1 = TR_102 ;
	7'h34 :
		RG_rl_90_t1 = TR_102 ;
	7'h35 :
		RG_rl_90_t1 = TR_102 ;
	7'h36 :
		RG_rl_90_t1 = TR_102 ;
	7'h37 :
		RG_rl_90_t1 = TR_102 ;
	7'h38 :
		RG_rl_90_t1 = TR_102 ;
	7'h39 :
		RG_rl_90_t1 = TR_102 ;
	7'h3a :
		RG_rl_90_t1 = TR_102 ;
	7'h3b :
		RG_rl_90_t1 = TR_102 ;
	7'h3c :
		RG_rl_90_t1 = TR_102 ;
	7'h3d :
		RG_rl_90_t1 = TR_102 ;
	7'h3e :
		RG_rl_90_t1 = TR_102 ;
	7'h3f :
		RG_rl_90_t1 = TR_102 ;
	7'h40 :
		RG_rl_90_t1 = TR_102 ;
	7'h41 :
		RG_rl_90_t1 = TR_102 ;
	7'h42 :
		RG_rl_90_t1 = TR_102 ;
	7'h43 :
		RG_rl_90_t1 = TR_102 ;
	7'h44 :
		RG_rl_90_t1 = TR_102 ;
	7'h45 :
		RG_rl_90_t1 = TR_102 ;
	7'h46 :
		RG_rl_90_t1 = TR_102 ;
	7'h47 :
		RG_rl_90_t1 = TR_102 ;
	7'h48 :
		RG_rl_90_t1 = TR_102 ;
	7'h49 :
		RG_rl_90_t1 = TR_102 ;
	7'h4a :
		RG_rl_90_t1 = TR_102 ;
	7'h4b :
		RG_rl_90_t1 = TR_102 ;
	7'h4c :
		RG_rl_90_t1 = TR_102 ;
	7'h4d :
		RG_rl_90_t1 = TR_102 ;
	7'h4e :
		RG_rl_90_t1 = TR_102 ;
	7'h4f :
		RG_rl_90_t1 = TR_102 ;
	7'h50 :
		RG_rl_90_t1 = TR_102 ;
	7'h51 :
		RG_rl_90_t1 = TR_102 ;
	7'h52 :
		RG_rl_90_t1 = TR_102 ;
	7'h53 :
		RG_rl_90_t1 = TR_102 ;
	7'h54 :
		RG_rl_90_t1 = TR_102 ;
	7'h55 :
		RG_rl_90_t1 = TR_102 ;
	7'h56 :
		RG_rl_90_t1 = TR_102 ;
	7'h57 :
		RG_rl_90_t1 = TR_102 ;
	7'h58 :
		RG_rl_90_t1 = TR_102 ;
	7'h59 :
		RG_rl_90_t1 = TR_102 ;
	7'h5a :
		RG_rl_90_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5b :
		RG_rl_90_t1 = TR_102 ;
	7'h5c :
		RG_rl_90_t1 = TR_102 ;
	7'h5d :
		RG_rl_90_t1 = TR_102 ;
	7'h5e :
		RG_rl_90_t1 = TR_102 ;
	7'h5f :
		RG_rl_90_t1 = TR_102 ;
	7'h60 :
		RG_rl_90_t1 = TR_102 ;
	7'h61 :
		RG_rl_90_t1 = TR_102 ;
	7'h62 :
		RG_rl_90_t1 = TR_102 ;
	7'h63 :
		RG_rl_90_t1 = TR_102 ;
	7'h64 :
		RG_rl_90_t1 = TR_102 ;
	7'h65 :
		RG_rl_90_t1 = TR_102 ;
	7'h66 :
		RG_rl_90_t1 = TR_102 ;
	7'h67 :
		RG_rl_90_t1 = TR_102 ;
	7'h68 :
		RG_rl_90_t1 = TR_102 ;
	7'h69 :
		RG_rl_90_t1 = TR_102 ;
	7'h6a :
		RG_rl_90_t1 = TR_102 ;
	7'h6b :
		RG_rl_90_t1 = TR_102 ;
	7'h6c :
		RG_rl_90_t1 = TR_102 ;
	7'h6d :
		RG_rl_90_t1 = TR_102 ;
	7'h6e :
		RG_rl_90_t1 = TR_102 ;
	7'h6f :
		RG_rl_90_t1 = TR_102 ;
	7'h70 :
		RG_rl_90_t1 = TR_102 ;
	7'h71 :
		RG_rl_90_t1 = TR_102 ;
	7'h72 :
		RG_rl_90_t1 = TR_102 ;
	7'h73 :
		RG_rl_90_t1 = TR_102 ;
	7'h74 :
		RG_rl_90_t1 = TR_102 ;
	7'h75 :
		RG_rl_90_t1 = TR_102 ;
	7'h76 :
		RG_rl_90_t1 = TR_102 ;
	7'h77 :
		RG_rl_90_t1 = TR_102 ;
	7'h78 :
		RG_rl_90_t1 = TR_102 ;
	7'h79 :
		RG_rl_90_t1 = TR_102 ;
	7'h7a :
		RG_rl_90_t1 = TR_102 ;
	7'h7b :
		RG_rl_90_t1 = TR_102 ;
	7'h7c :
		RG_rl_90_t1 = TR_102 ;
	7'h7d :
		RG_rl_90_t1 = TR_102 ;
	7'h7e :
		RG_rl_90_t1 = TR_102 ;
	7'h7f :
		RG_rl_90_t1 = TR_102 ;
	default :
		RG_rl_90_t1 = 9'hx ;
	endcase
always @ ( RG_rl_90_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_31 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_90_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h5a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_90_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_31 )
		| ( { 9{ U_569 } } & RG_rl_90_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_90_en = ( U_570 | RG_rl_90_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_90_en )
		RG_rl_90 <= RG_rl_90_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_103 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_91_t1 = TR_103 ;
	7'h01 :
		RG_rl_91_t1 = TR_103 ;
	7'h02 :
		RG_rl_91_t1 = TR_103 ;
	7'h03 :
		RG_rl_91_t1 = TR_103 ;
	7'h04 :
		RG_rl_91_t1 = TR_103 ;
	7'h05 :
		RG_rl_91_t1 = TR_103 ;
	7'h06 :
		RG_rl_91_t1 = TR_103 ;
	7'h07 :
		RG_rl_91_t1 = TR_103 ;
	7'h08 :
		RG_rl_91_t1 = TR_103 ;
	7'h09 :
		RG_rl_91_t1 = TR_103 ;
	7'h0a :
		RG_rl_91_t1 = TR_103 ;
	7'h0b :
		RG_rl_91_t1 = TR_103 ;
	7'h0c :
		RG_rl_91_t1 = TR_103 ;
	7'h0d :
		RG_rl_91_t1 = TR_103 ;
	7'h0e :
		RG_rl_91_t1 = TR_103 ;
	7'h0f :
		RG_rl_91_t1 = TR_103 ;
	7'h10 :
		RG_rl_91_t1 = TR_103 ;
	7'h11 :
		RG_rl_91_t1 = TR_103 ;
	7'h12 :
		RG_rl_91_t1 = TR_103 ;
	7'h13 :
		RG_rl_91_t1 = TR_103 ;
	7'h14 :
		RG_rl_91_t1 = TR_103 ;
	7'h15 :
		RG_rl_91_t1 = TR_103 ;
	7'h16 :
		RG_rl_91_t1 = TR_103 ;
	7'h17 :
		RG_rl_91_t1 = TR_103 ;
	7'h18 :
		RG_rl_91_t1 = TR_103 ;
	7'h19 :
		RG_rl_91_t1 = TR_103 ;
	7'h1a :
		RG_rl_91_t1 = TR_103 ;
	7'h1b :
		RG_rl_91_t1 = TR_103 ;
	7'h1c :
		RG_rl_91_t1 = TR_103 ;
	7'h1d :
		RG_rl_91_t1 = TR_103 ;
	7'h1e :
		RG_rl_91_t1 = TR_103 ;
	7'h1f :
		RG_rl_91_t1 = TR_103 ;
	7'h20 :
		RG_rl_91_t1 = TR_103 ;
	7'h21 :
		RG_rl_91_t1 = TR_103 ;
	7'h22 :
		RG_rl_91_t1 = TR_103 ;
	7'h23 :
		RG_rl_91_t1 = TR_103 ;
	7'h24 :
		RG_rl_91_t1 = TR_103 ;
	7'h25 :
		RG_rl_91_t1 = TR_103 ;
	7'h26 :
		RG_rl_91_t1 = TR_103 ;
	7'h27 :
		RG_rl_91_t1 = TR_103 ;
	7'h28 :
		RG_rl_91_t1 = TR_103 ;
	7'h29 :
		RG_rl_91_t1 = TR_103 ;
	7'h2a :
		RG_rl_91_t1 = TR_103 ;
	7'h2b :
		RG_rl_91_t1 = TR_103 ;
	7'h2c :
		RG_rl_91_t1 = TR_103 ;
	7'h2d :
		RG_rl_91_t1 = TR_103 ;
	7'h2e :
		RG_rl_91_t1 = TR_103 ;
	7'h2f :
		RG_rl_91_t1 = TR_103 ;
	7'h30 :
		RG_rl_91_t1 = TR_103 ;
	7'h31 :
		RG_rl_91_t1 = TR_103 ;
	7'h32 :
		RG_rl_91_t1 = TR_103 ;
	7'h33 :
		RG_rl_91_t1 = TR_103 ;
	7'h34 :
		RG_rl_91_t1 = TR_103 ;
	7'h35 :
		RG_rl_91_t1 = TR_103 ;
	7'h36 :
		RG_rl_91_t1 = TR_103 ;
	7'h37 :
		RG_rl_91_t1 = TR_103 ;
	7'h38 :
		RG_rl_91_t1 = TR_103 ;
	7'h39 :
		RG_rl_91_t1 = TR_103 ;
	7'h3a :
		RG_rl_91_t1 = TR_103 ;
	7'h3b :
		RG_rl_91_t1 = TR_103 ;
	7'h3c :
		RG_rl_91_t1 = TR_103 ;
	7'h3d :
		RG_rl_91_t1 = TR_103 ;
	7'h3e :
		RG_rl_91_t1 = TR_103 ;
	7'h3f :
		RG_rl_91_t1 = TR_103 ;
	7'h40 :
		RG_rl_91_t1 = TR_103 ;
	7'h41 :
		RG_rl_91_t1 = TR_103 ;
	7'h42 :
		RG_rl_91_t1 = TR_103 ;
	7'h43 :
		RG_rl_91_t1 = TR_103 ;
	7'h44 :
		RG_rl_91_t1 = TR_103 ;
	7'h45 :
		RG_rl_91_t1 = TR_103 ;
	7'h46 :
		RG_rl_91_t1 = TR_103 ;
	7'h47 :
		RG_rl_91_t1 = TR_103 ;
	7'h48 :
		RG_rl_91_t1 = TR_103 ;
	7'h49 :
		RG_rl_91_t1 = TR_103 ;
	7'h4a :
		RG_rl_91_t1 = TR_103 ;
	7'h4b :
		RG_rl_91_t1 = TR_103 ;
	7'h4c :
		RG_rl_91_t1 = TR_103 ;
	7'h4d :
		RG_rl_91_t1 = TR_103 ;
	7'h4e :
		RG_rl_91_t1 = TR_103 ;
	7'h4f :
		RG_rl_91_t1 = TR_103 ;
	7'h50 :
		RG_rl_91_t1 = TR_103 ;
	7'h51 :
		RG_rl_91_t1 = TR_103 ;
	7'h52 :
		RG_rl_91_t1 = TR_103 ;
	7'h53 :
		RG_rl_91_t1 = TR_103 ;
	7'h54 :
		RG_rl_91_t1 = TR_103 ;
	7'h55 :
		RG_rl_91_t1 = TR_103 ;
	7'h56 :
		RG_rl_91_t1 = TR_103 ;
	7'h57 :
		RG_rl_91_t1 = TR_103 ;
	7'h58 :
		RG_rl_91_t1 = TR_103 ;
	7'h59 :
		RG_rl_91_t1 = TR_103 ;
	7'h5a :
		RG_rl_91_t1 = TR_103 ;
	7'h5b :
		RG_rl_91_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5c :
		RG_rl_91_t1 = TR_103 ;
	7'h5d :
		RG_rl_91_t1 = TR_103 ;
	7'h5e :
		RG_rl_91_t1 = TR_103 ;
	7'h5f :
		RG_rl_91_t1 = TR_103 ;
	7'h60 :
		RG_rl_91_t1 = TR_103 ;
	7'h61 :
		RG_rl_91_t1 = TR_103 ;
	7'h62 :
		RG_rl_91_t1 = TR_103 ;
	7'h63 :
		RG_rl_91_t1 = TR_103 ;
	7'h64 :
		RG_rl_91_t1 = TR_103 ;
	7'h65 :
		RG_rl_91_t1 = TR_103 ;
	7'h66 :
		RG_rl_91_t1 = TR_103 ;
	7'h67 :
		RG_rl_91_t1 = TR_103 ;
	7'h68 :
		RG_rl_91_t1 = TR_103 ;
	7'h69 :
		RG_rl_91_t1 = TR_103 ;
	7'h6a :
		RG_rl_91_t1 = TR_103 ;
	7'h6b :
		RG_rl_91_t1 = TR_103 ;
	7'h6c :
		RG_rl_91_t1 = TR_103 ;
	7'h6d :
		RG_rl_91_t1 = TR_103 ;
	7'h6e :
		RG_rl_91_t1 = TR_103 ;
	7'h6f :
		RG_rl_91_t1 = TR_103 ;
	7'h70 :
		RG_rl_91_t1 = TR_103 ;
	7'h71 :
		RG_rl_91_t1 = TR_103 ;
	7'h72 :
		RG_rl_91_t1 = TR_103 ;
	7'h73 :
		RG_rl_91_t1 = TR_103 ;
	7'h74 :
		RG_rl_91_t1 = TR_103 ;
	7'h75 :
		RG_rl_91_t1 = TR_103 ;
	7'h76 :
		RG_rl_91_t1 = TR_103 ;
	7'h77 :
		RG_rl_91_t1 = TR_103 ;
	7'h78 :
		RG_rl_91_t1 = TR_103 ;
	7'h79 :
		RG_rl_91_t1 = TR_103 ;
	7'h7a :
		RG_rl_91_t1 = TR_103 ;
	7'h7b :
		RG_rl_91_t1 = TR_103 ;
	7'h7c :
		RG_rl_91_t1 = TR_103 ;
	7'h7d :
		RG_rl_91_t1 = TR_103 ;
	7'h7e :
		RG_rl_91_t1 = TR_103 ;
	7'h7f :
		RG_rl_91_t1 = TR_103 ;
	default :
		RG_rl_91_t1 = 9'hx ;
	endcase
always @ ( RG_rl_91_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_32 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_91_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h5b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_91_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_32 )
		| ( { 9{ U_569 } } & RG_rl_91_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_91_en = ( U_570 | RG_rl_91_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_91_en )
		RG_rl_91 <= RG_rl_91_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_104 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_92_t1 = TR_104 ;
	7'h01 :
		RG_rl_92_t1 = TR_104 ;
	7'h02 :
		RG_rl_92_t1 = TR_104 ;
	7'h03 :
		RG_rl_92_t1 = TR_104 ;
	7'h04 :
		RG_rl_92_t1 = TR_104 ;
	7'h05 :
		RG_rl_92_t1 = TR_104 ;
	7'h06 :
		RG_rl_92_t1 = TR_104 ;
	7'h07 :
		RG_rl_92_t1 = TR_104 ;
	7'h08 :
		RG_rl_92_t1 = TR_104 ;
	7'h09 :
		RG_rl_92_t1 = TR_104 ;
	7'h0a :
		RG_rl_92_t1 = TR_104 ;
	7'h0b :
		RG_rl_92_t1 = TR_104 ;
	7'h0c :
		RG_rl_92_t1 = TR_104 ;
	7'h0d :
		RG_rl_92_t1 = TR_104 ;
	7'h0e :
		RG_rl_92_t1 = TR_104 ;
	7'h0f :
		RG_rl_92_t1 = TR_104 ;
	7'h10 :
		RG_rl_92_t1 = TR_104 ;
	7'h11 :
		RG_rl_92_t1 = TR_104 ;
	7'h12 :
		RG_rl_92_t1 = TR_104 ;
	7'h13 :
		RG_rl_92_t1 = TR_104 ;
	7'h14 :
		RG_rl_92_t1 = TR_104 ;
	7'h15 :
		RG_rl_92_t1 = TR_104 ;
	7'h16 :
		RG_rl_92_t1 = TR_104 ;
	7'h17 :
		RG_rl_92_t1 = TR_104 ;
	7'h18 :
		RG_rl_92_t1 = TR_104 ;
	7'h19 :
		RG_rl_92_t1 = TR_104 ;
	7'h1a :
		RG_rl_92_t1 = TR_104 ;
	7'h1b :
		RG_rl_92_t1 = TR_104 ;
	7'h1c :
		RG_rl_92_t1 = TR_104 ;
	7'h1d :
		RG_rl_92_t1 = TR_104 ;
	7'h1e :
		RG_rl_92_t1 = TR_104 ;
	7'h1f :
		RG_rl_92_t1 = TR_104 ;
	7'h20 :
		RG_rl_92_t1 = TR_104 ;
	7'h21 :
		RG_rl_92_t1 = TR_104 ;
	7'h22 :
		RG_rl_92_t1 = TR_104 ;
	7'h23 :
		RG_rl_92_t1 = TR_104 ;
	7'h24 :
		RG_rl_92_t1 = TR_104 ;
	7'h25 :
		RG_rl_92_t1 = TR_104 ;
	7'h26 :
		RG_rl_92_t1 = TR_104 ;
	7'h27 :
		RG_rl_92_t1 = TR_104 ;
	7'h28 :
		RG_rl_92_t1 = TR_104 ;
	7'h29 :
		RG_rl_92_t1 = TR_104 ;
	7'h2a :
		RG_rl_92_t1 = TR_104 ;
	7'h2b :
		RG_rl_92_t1 = TR_104 ;
	7'h2c :
		RG_rl_92_t1 = TR_104 ;
	7'h2d :
		RG_rl_92_t1 = TR_104 ;
	7'h2e :
		RG_rl_92_t1 = TR_104 ;
	7'h2f :
		RG_rl_92_t1 = TR_104 ;
	7'h30 :
		RG_rl_92_t1 = TR_104 ;
	7'h31 :
		RG_rl_92_t1 = TR_104 ;
	7'h32 :
		RG_rl_92_t1 = TR_104 ;
	7'h33 :
		RG_rl_92_t1 = TR_104 ;
	7'h34 :
		RG_rl_92_t1 = TR_104 ;
	7'h35 :
		RG_rl_92_t1 = TR_104 ;
	7'h36 :
		RG_rl_92_t1 = TR_104 ;
	7'h37 :
		RG_rl_92_t1 = TR_104 ;
	7'h38 :
		RG_rl_92_t1 = TR_104 ;
	7'h39 :
		RG_rl_92_t1 = TR_104 ;
	7'h3a :
		RG_rl_92_t1 = TR_104 ;
	7'h3b :
		RG_rl_92_t1 = TR_104 ;
	7'h3c :
		RG_rl_92_t1 = TR_104 ;
	7'h3d :
		RG_rl_92_t1 = TR_104 ;
	7'h3e :
		RG_rl_92_t1 = TR_104 ;
	7'h3f :
		RG_rl_92_t1 = TR_104 ;
	7'h40 :
		RG_rl_92_t1 = TR_104 ;
	7'h41 :
		RG_rl_92_t1 = TR_104 ;
	7'h42 :
		RG_rl_92_t1 = TR_104 ;
	7'h43 :
		RG_rl_92_t1 = TR_104 ;
	7'h44 :
		RG_rl_92_t1 = TR_104 ;
	7'h45 :
		RG_rl_92_t1 = TR_104 ;
	7'h46 :
		RG_rl_92_t1 = TR_104 ;
	7'h47 :
		RG_rl_92_t1 = TR_104 ;
	7'h48 :
		RG_rl_92_t1 = TR_104 ;
	7'h49 :
		RG_rl_92_t1 = TR_104 ;
	7'h4a :
		RG_rl_92_t1 = TR_104 ;
	7'h4b :
		RG_rl_92_t1 = TR_104 ;
	7'h4c :
		RG_rl_92_t1 = TR_104 ;
	7'h4d :
		RG_rl_92_t1 = TR_104 ;
	7'h4e :
		RG_rl_92_t1 = TR_104 ;
	7'h4f :
		RG_rl_92_t1 = TR_104 ;
	7'h50 :
		RG_rl_92_t1 = TR_104 ;
	7'h51 :
		RG_rl_92_t1 = TR_104 ;
	7'h52 :
		RG_rl_92_t1 = TR_104 ;
	7'h53 :
		RG_rl_92_t1 = TR_104 ;
	7'h54 :
		RG_rl_92_t1 = TR_104 ;
	7'h55 :
		RG_rl_92_t1 = TR_104 ;
	7'h56 :
		RG_rl_92_t1 = TR_104 ;
	7'h57 :
		RG_rl_92_t1 = TR_104 ;
	7'h58 :
		RG_rl_92_t1 = TR_104 ;
	7'h59 :
		RG_rl_92_t1 = TR_104 ;
	7'h5a :
		RG_rl_92_t1 = TR_104 ;
	7'h5b :
		RG_rl_92_t1 = TR_104 ;
	7'h5c :
		RG_rl_92_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5d :
		RG_rl_92_t1 = TR_104 ;
	7'h5e :
		RG_rl_92_t1 = TR_104 ;
	7'h5f :
		RG_rl_92_t1 = TR_104 ;
	7'h60 :
		RG_rl_92_t1 = TR_104 ;
	7'h61 :
		RG_rl_92_t1 = TR_104 ;
	7'h62 :
		RG_rl_92_t1 = TR_104 ;
	7'h63 :
		RG_rl_92_t1 = TR_104 ;
	7'h64 :
		RG_rl_92_t1 = TR_104 ;
	7'h65 :
		RG_rl_92_t1 = TR_104 ;
	7'h66 :
		RG_rl_92_t1 = TR_104 ;
	7'h67 :
		RG_rl_92_t1 = TR_104 ;
	7'h68 :
		RG_rl_92_t1 = TR_104 ;
	7'h69 :
		RG_rl_92_t1 = TR_104 ;
	7'h6a :
		RG_rl_92_t1 = TR_104 ;
	7'h6b :
		RG_rl_92_t1 = TR_104 ;
	7'h6c :
		RG_rl_92_t1 = TR_104 ;
	7'h6d :
		RG_rl_92_t1 = TR_104 ;
	7'h6e :
		RG_rl_92_t1 = TR_104 ;
	7'h6f :
		RG_rl_92_t1 = TR_104 ;
	7'h70 :
		RG_rl_92_t1 = TR_104 ;
	7'h71 :
		RG_rl_92_t1 = TR_104 ;
	7'h72 :
		RG_rl_92_t1 = TR_104 ;
	7'h73 :
		RG_rl_92_t1 = TR_104 ;
	7'h74 :
		RG_rl_92_t1 = TR_104 ;
	7'h75 :
		RG_rl_92_t1 = TR_104 ;
	7'h76 :
		RG_rl_92_t1 = TR_104 ;
	7'h77 :
		RG_rl_92_t1 = TR_104 ;
	7'h78 :
		RG_rl_92_t1 = TR_104 ;
	7'h79 :
		RG_rl_92_t1 = TR_104 ;
	7'h7a :
		RG_rl_92_t1 = TR_104 ;
	7'h7b :
		RG_rl_92_t1 = TR_104 ;
	7'h7c :
		RG_rl_92_t1 = TR_104 ;
	7'h7d :
		RG_rl_92_t1 = TR_104 ;
	7'h7e :
		RG_rl_92_t1 = TR_104 ;
	7'h7f :
		RG_rl_92_t1 = TR_104 ;
	default :
		RG_rl_92_t1 = 9'hx ;
	endcase
always @ ( RG_rl_92_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_33 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_92_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h5c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_92_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_33 )
		| ( { 9{ U_569 } } & RG_rl_92_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_92_en = ( U_570 | RG_rl_92_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_92_en )
		RG_rl_92 <= RG_rl_92_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_105 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_93_t1 = TR_105 ;
	7'h01 :
		RG_rl_93_t1 = TR_105 ;
	7'h02 :
		RG_rl_93_t1 = TR_105 ;
	7'h03 :
		RG_rl_93_t1 = TR_105 ;
	7'h04 :
		RG_rl_93_t1 = TR_105 ;
	7'h05 :
		RG_rl_93_t1 = TR_105 ;
	7'h06 :
		RG_rl_93_t1 = TR_105 ;
	7'h07 :
		RG_rl_93_t1 = TR_105 ;
	7'h08 :
		RG_rl_93_t1 = TR_105 ;
	7'h09 :
		RG_rl_93_t1 = TR_105 ;
	7'h0a :
		RG_rl_93_t1 = TR_105 ;
	7'h0b :
		RG_rl_93_t1 = TR_105 ;
	7'h0c :
		RG_rl_93_t1 = TR_105 ;
	7'h0d :
		RG_rl_93_t1 = TR_105 ;
	7'h0e :
		RG_rl_93_t1 = TR_105 ;
	7'h0f :
		RG_rl_93_t1 = TR_105 ;
	7'h10 :
		RG_rl_93_t1 = TR_105 ;
	7'h11 :
		RG_rl_93_t1 = TR_105 ;
	7'h12 :
		RG_rl_93_t1 = TR_105 ;
	7'h13 :
		RG_rl_93_t1 = TR_105 ;
	7'h14 :
		RG_rl_93_t1 = TR_105 ;
	7'h15 :
		RG_rl_93_t1 = TR_105 ;
	7'h16 :
		RG_rl_93_t1 = TR_105 ;
	7'h17 :
		RG_rl_93_t1 = TR_105 ;
	7'h18 :
		RG_rl_93_t1 = TR_105 ;
	7'h19 :
		RG_rl_93_t1 = TR_105 ;
	7'h1a :
		RG_rl_93_t1 = TR_105 ;
	7'h1b :
		RG_rl_93_t1 = TR_105 ;
	7'h1c :
		RG_rl_93_t1 = TR_105 ;
	7'h1d :
		RG_rl_93_t1 = TR_105 ;
	7'h1e :
		RG_rl_93_t1 = TR_105 ;
	7'h1f :
		RG_rl_93_t1 = TR_105 ;
	7'h20 :
		RG_rl_93_t1 = TR_105 ;
	7'h21 :
		RG_rl_93_t1 = TR_105 ;
	7'h22 :
		RG_rl_93_t1 = TR_105 ;
	7'h23 :
		RG_rl_93_t1 = TR_105 ;
	7'h24 :
		RG_rl_93_t1 = TR_105 ;
	7'h25 :
		RG_rl_93_t1 = TR_105 ;
	7'h26 :
		RG_rl_93_t1 = TR_105 ;
	7'h27 :
		RG_rl_93_t1 = TR_105 ;
	7'h28 :
		RG_rl_93_t1 = TR_105 ;
	7'h29 :
		RG_rl_93_t1 = TR_105 ;
	7'h2a :
		RG_rl_93_t1 = TR_105 ;
	7'h2b :
		RG_rl_93_t1 = TR_105 ;
	7'h2c :
		RG_rl_93_t1 = TR_105 ;
	7'h2d :
		RG_rl_93_t1 = TR_105 ;
	7'h2e :
		RG_rl_93_t1 = TR_105 ;
	7'h2f :
		RG_rl_93_t1 = TR_105 ;
	7'h30 :
		RG_rl_93_t1 = TR_105 ;
	7'h31 :
		RG_rl_93_t1 = TR_105 ;
	7'h32 :
		RG_rl_93_t1 = TR_105 ;
	7'h33 :
		RG_rl_93_t1 = TR_105 ;
	7'h34 :
		RG_rl_93_t1 = TR_105 ;
	7'h35 :
		RG_rl_93_t1 = TR_105 ;
	7'h36 :
		RG_rl_93_t1 = TR_105 ;
	7'h37 :
		RG_rl_93_t1 = TR_105 ;
	7'h38 :
		RG_rl_93_t1 = TR_105 ;
	7'h39 :
		RG_rl_93_t1 = TR_105 ;
	7'h3a :
		RG_rl_93_t1 = TR_105 ;
	7'h3b :
		RG_rl_93_t1 = TR_105 ;
	7'h3c :
		RG_rl_93_t1 = TR_105 ;
	7'h3d :
		RG_rl_93_t1 = TR_105 ;
	7'h3e :
		RG_rl_93_t1 = TR_105 ;
	7'h3f :
		RG_rl_93_t1 = TR_105 ;
	7'h40 :
		RG_rl_93_t1 = TR_105 ;
	7'h41 :
		RG_rl_93_t1 = TR_105 ;
	7'h42 :
		RG_rl_93_t1 = TR_105 ;
	7'h43 :
		RG_rl_93_t1 = TR_105 ;
	7'h44 :
		RG_rl_93_t1 = TR_105 ;
	7'h45 :
		RG_rl_93_t1 = TR_105 ;
	7'h46 :
		RG_rl_93_t1 = TR_105 ;
	7'h47 :
		RG_rl_93_t1 = TR_105 ;
	7'h48 :
		RG_rl_93_t1 = TR_105 ;
	7'h49 :
		RG_rl_93_t1 = TR_105 ;
	7'h4a :
		RG_rl_93_t1 = TR_105 ;
	7'h4b :
		RG_rl_93_t1 = TR_105 ;
	7'h4c :
		RG_rl_93_t1 = TR_105 ;
	7'h4d :
		RG_rl_93_t1 = TR_105 ;
	7'h4e :
		RG_rl_93_t1 = TR_105 ;
	7'h4f :
		RG_rl_93_t1 = TR_105 ;
	7'h50 :
		RG_rl_93_t1 = TR_105 ;
	7'h51 :
		RG_rl_93_t1 = TR_105 ;
	7'h52 :
		RG_rl_93_t1 = TR_105 ;
	7'h53 :
		RG_rl_93_t1 = TR_105 ;
	7'h54 :
		RG_rl_93_t1 = TR_105 ;
	7'h55 :
		RG_rl_93_t1 = TR_105 ;
	7'h56 :
		RG_rl_93_t1 = TR_105 ;
	7'h57 :
		RG_rl_93_t1 = TR_105 ;
	7'h58 :
		RG_rl_93_t1 = TR_105 ;
	7'h59 :
		RG_rl_93_t1 = TR_105 ;
	7'h5a :
		RG_rl_93_t1 = TR_105 ;
	7'h5b :
		RG_rl_93_t1 = TR_105 ;
	7'h5c :
		RG_rl_93_t1 = TR_105 ;
	7'h5d :
		RG_rl_93_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5e :
		RG_rl_93_t1 = TR_105 ;
	7'h5f :
		RG_rl_93_t1 = TR_105 ;
	7'h60 :
		RG_rl_93_t1 = TR_105 ;
	7'h61 :
		RG_rl_93_t1 = TR_105 ;
	7'h62 :
		RG_rl_93_t1 = TR_105 ;
	7'h63 :
		RG_rl_93_t1 = TR_105 ;
	7'h64 :
		RG_rl_93_t1 = TR_105 ;
	7'h65 :
		RG_rl_93_t1 = TR_105 ;
	7'h66 :
		RG_rl_93_t1 = TR_105 ;
	7'h67 :
		RG_rl_93_t1 = TR_105 ;
	7'h68 :
		RG_rl_93_t1 = TR_105 ;
	7'h69 :
		RG_rl_93_t1 = TR_105 ;
	7'h6a :
		RG_rl_93_t1 = TR_105 ;
	7'h6b :
		RG_rl_93_t1 = TR_105 ;
	7'h6c :
		RG_rl_93_t1 = TR_105 ;
	7'h6d :
		RG_rl_93_t1 = TR_105 ;
	7'h6e :
		RG_rl_93_t1 = TR_105 ;
	7'h6f :
		RG_rl_93_t1 = TR_105 ;
	7'h70 :
		RG_rl_93_t1 = TR_105 ;
	7'h71 :
		RG_rl_93_t1 = TR_105 ;
	7'h72 :
		RG_rl_93_t1 = TR_105 ;
	7'h73 :
		RG_rl_93_t1 = TR_105 ;
	7'h74 :
		RG_rl_93_t1 = TR_105 ;
	7'h75 :
		RG_rl_93_t1 = TR_105 ;
	7'h76 :
		RG_rl_93_t1 = TR_105 ;
	7'h77 :
		RG_rl_93_t1 = TR_105 ;
	7'h78 :
		RG_rl_93_t1 = TR_105 ;
	7'h79 :
		RG_rl_93_t1 = TR_105 ;
	7'h7a :
		RG_rl_93_t1 = TR_105 ;
	7'h7b :
		RG_rl_93_t1 = TR_105 ;
	7'h7c :
		RG_rl_93_t1 = TR_105 ;
	7'h7d :
		RG_rl_93_t1 = TR_105 ;
	7'h7e :
		RG_rl_93_t1 = TR_105 ;
	7'h7f :
		RG_rl_93_t1 = TR_105 ;
	default :
		RG_rl_93_t1 = 9'hx ;
	endcase
always @ ( RG_rl_93_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_34 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_93_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h5d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_93_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_34 )
		| ( { 9{ U_569 } } & RG_rl_93_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_93_en = ( U_570 | RG_rl_93_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_93_en )
		RG_rl_93 <= RG_rl_93_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_106 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_94_t1 = TR_106 ;
	7'h01 :
		RG_rl_94_t1 = TR_106 ;
	7'h02 :
		RG_rl_94_t1 = TR_106 ;
	7'h03 :
		RG_rl_94_t1 = TR_106 ;
	7'h04 :
		RG_rl_94_t1 = TR_106 ;
	7'h05 :
		RG_rl_94_t1 = TR_106 ;
	7'h06 :
		RG_rl_94_t1 = TR_106 ;
	7'h07 :
		RG_rl_94_t1 = TR_106 ;
	7'h08 :
		RG_rl_94_t1 = TR_106 ;
	7'h09 :
		RG_rl_94_t1 = TR_106 ;
	7'h0a :
		RG_rl_94_t1 = TR_106 ;
	7'h0b :
		RG_rl_94_t1 = TR_106 ;
	7'h0c :
		RG_rl_94_t1 = TR_106 ;
	7'h0d :
		RG_rl_94_t1 = TR_106 ;
	7'h0e :
		RG_rl_94_t1 = TR_106 ;
	7'h0f :
		RG_rl_94_t1 = TR_106 ;
	7'h10 :
		RG_rl_94_t1 = TR_106 ;
	7'h11 :
		RG_rl_94_t1 = TR_106 ;
	7'h12 :
		RG_rl_94_t1 = TR_106 ;
	7'h13 :
		RG_rl_94_t1 = TR_106 ;
	7'h14 :
		RG_rl_94_t1 = TR_106 ;
	7'h15 :
		RG_rl_94_t1 = TR_106 ;
	7'h16 :
		RG_rl_94_t1 = TR_106 ;
	7'h17 :
		RG_rl_94_t1 = TR_106 ;
	7'h18 :
		RG_rl_94_t1 = TR_106 ;
	7'h19 :
		RG_rl_94_t1 = TR_106 ;
	7'h1a :
		RG_rl_94_t1 = TR_106 ;
	7'h1b :
		RG_rl_94_t1 = TR_106 ;
	7'h1c :
		RG_rl_94_t1 = TR_106 ;
	7'h1d :
		RG_rl_94_t1 = TR_106 ;
	7'h1e :
		RG_rl_94_t1 = TR_106 ;
	7'h1f :
		RG_rl_94_t1 = TR_106 ;
	7'h20 :
		RG_rl_94_t1 = TR_106 ;
	7'h21 :
		RG_rl_94_t1 = TR_106 ;
	7'h22 :
		RG_rl_94_t1 = TR_106 ;
	7'h23 :
		RG_rl_94_t1 = TR_106 ;
	7'h24 :
		RG_rl_94_t1 = TR_106 ;
	7'h25 :
		RG_rl_94_t1 = TR_106 ;
	7'h26 :
		RG_rl_94_t1 = TR_106 ;
	7'h27 :
		RG_rl_94_t1 = TR_106 ;
	7'h28 :
		RG_rl_94_t1 = TR_106 ;
	7'h29 :
		RG_rl_94_t1 = TR_106 ;
	7'h2a :
		RG_rl_94_t1 = TR_106 ;
	7'h2b :
		RG_rl_94_t1 = TR_106 ;
	7'h2c :
		RG_rl_94_t1 = TR_106 ;
	7'h2d :
		RG_rl_94_t1 = TR_106 ;
	7'h2e :
		RG_rl_94_t1 = TR_106 ;
	7'h2f :
		RG_rl_94_t1 = TR_106 ;
	7'h30 :
		RG_rl_94_t1 = TR_106 ;
	7'h31 :
		RG_rl_94_t1 = TR_106 ;
	7'h32 :
		RG_rl_94_t1 = TR_106 ;
	7'h33 :
		RG_rl_94_t1 = TR_106 ;
	7'h34 :
		RG_rl_94_t1 = TR_106 ;
	7'h35 :
		RG_rl_94_t1 = TR_106 ;
	7'h36 :
		RG_rl_94_t1 = TR_106 ;
	7'h37 :
		RG_rl_94_t1 = TR_106 ;
	7'h38 :
		RG_rl_94_t1 = TR_106 ;
	7'h39 :
		RG_rl_94_t1 = TR_106 ;
	7'h3a :
		RG_rl_94_t1 = TR_106 ;
	7'h3b :
		RG_rl_94_t1 = TR_106 ;
	7'h3c :
		RG_rl_94_t1 = TR_106 ;
	7'h3d :
		RG_rl_94_t1 = TR_106 ;
	7'h3e :
		RG_rl_94_t1 = TR_106 ;
	7'h3f :
		RG_rl_94_t1 = TR_106 ;
	7'h40 :
		RG_rl_94_t1 = TR_106 ;
	7'h41 :
		RG_rl_94_t1 = TR_106 ;
	7'h42 :
		RG_rl_94_t1 = TR_106 ;
	7'h43 :
		RG_rl_94_t1 = TR_106 ;
	7'h44 :
		RG_rl_94_t1 = TR_106 ;
	7'h45 :
		RG_rl_94_t1 = TR_106 ;
	7'h46 :
		RG_rl_94_t1 = TR_106 ;
	7'h47 :
		RG_rl_94_t1 = TR_106 ;
	7'h48 :
		RG_rl_94_t1 = TR_106 ;
	7'h49 :
		RG_rl_94_t1 = TR_106 ;
	7'h4a :
		RG_rl_94_t1 = TR_106 ;
	7'h4b :
		RG_rl_94_t1 = TR_106 ;
	7'h4c :
		RG_rl_94_t1 = TR_106 ;
	7'h4d :
		RG_rl_94_t1 = TR_106 ;
	7'h4e :
		RG_rl_94_t1 = TR_106 ;
	7'h4f :
		RG_rl_94_t1 = TR_106 ;
	7'h50 :
		RG_rl_94_t1 = TR_106 ;
	7'h51 :
		RG_rl_94_t1 = TR_106 ;
	7'h52 :
		RG_rl_94_t1 = TR_106 ;
	7'h53 :
		RG_rl_94_t1 = TR_106 ;
	7'h54 :
		RG_rl_94_t1 = TR_106 ;
	7'h55 :
		RG_rl_94_t1 = TR_106 ;
	7'h56 :
		RG_rl_94_t1 = TR_106 ;
	7'h57 :
		RG_rl_94_t1 = TR_106 ;
	7'h58 :
		RG_rl_94_t1 = TR_106 ;
	7'h59 :
		RG_rl_94_t1 = TR_106 ;
	7'h5a :
		RG_rl_94_t1 = TR_106 ;
	7'h5b :
		RG_rl_94_t1 = TR_106 ;
	7'h5c :
		RG_rl_94_t1 = TR_106 ;
	7'h5d :
		RG_rl_94_t1 = TR_106 ;
	7'h5e :
		RG_rl_94_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h5f :
		RG_rl_94_t1 = TR_106 ;
	7'h60 :
		RG_rl_94_t1 = TR_106 ;
	7'h61 :
		RG_rl_94_t1 = TR_106 ;
	7'h62 :
		RG_rl_94_t1 = TR_106 ;
	7'h63 :
		RG_rl_94_t1 = TR_106 ;
	7'h64 :
		RG_rl_94_t1 = TR_106 ;
	7'h65 :
		RG_rl_94_t1 = TR_106 ;
	7'h66 :
		RG_rl_94_t1 = TR_106 ;
	7'h67 :
		RG_rl_94_t1 = TR_106 ;
	7'h68 :
		RG_rl_94_t1 = TR_106 ;
	7'h69 :
		RG_rl_94_t1 = TR_106 ;
	7'h6a :
		RG_rl_94_t1 = TR_106 ;
	7'h6b :
		RG_rl_94_t1 = TR_106 ;
	7'h6c :
		RG_rl_94_t1 = TR_106 ;
	7'h6d :
		RG_rl_94_t1 = TR_106 ;
	7'h6e :
		RG_rl_94_t1 = TR_106 ;
	7'h6f :
		RG_rl_94_t1 = TR_106 ;
	7'h70 :
		RG_rl_94_t1 = TR_106 ;
	7'h71 :
		RG_rl_94_t1 = TR_106 ;
	7'h72 :
		RG_rl_94_t1 = TR_106 ;
	7'h73 :
		RG_rl_94_t1 = TR_106 ;
	7'h74 :
		RG_rl_94_t1 = TR_106 ;
	7'h75 :
		RG_rl_94_t1 = TR_106 ;
	7'h76 :
		RG_rl_94_t1 = TR_106 ;
	7'h77 :
		RG_rl_94_t1 = TR_106 ;
	7'h78 :
		RG_rl_94_t1 = TR_106 ;
	7'h79 :
		RG_rl_94_t1 = TR_106 ;
	7'h7a :
		RG_rl_94_t1 = TR_106 ;
	7'h7b :
		RG_rl_94_t1 = TR_106 ;
	7'h7c :
		RG_rl_94_t1 = TR_106 ;
	7'h7d :
		RG_rl_94_t1 = TR_106 ;
	7'h7e :
		RG_rl_94_t1 = TR_106 ;
	7'h7f :
		RG_rl_94_t1 = TR_106 ;
	default :
		RG_rl_94_t1 = 9'hx ;
	endcase
always @ ( RG_rl_94_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_35 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_94_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h5e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_94_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_35 )
		| ( { 9{ U_569 } } & RG_rl_94_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_94_en = ( U_570 | RG_rl_94_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_94_en )
		RG_rl_94 <= RG_rl_94_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_107 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_95_t1 = TR_107 ;
	7'h01 :
		RG_rl_95_t1 = TR_107 ;
	7'h02 :
		RG_rl_95_t1 = TR_107 ;
	7'h03 :
		RG_rl_95_t1 = TR_107 ;
	7'h04 :
		RG_rl_95_t1 = TR_107 ;
	7'h05 :
		RG_rl_95_t1 = TR_107 ;
	7'h06 :
		RG_rl_95_t1 = TR_107 ;
	7'h07 :
		RG_rl_95_t1 = TR_107 ;
	7'h08 :
		RG_rl_95_t1 = TR_107 ;
	7'h09 :
		RG_rl_95_t1 = TR_107 ;
	7'h0a :
		RG_rl_95_t1 = TR_107 ;
	7'h0b :
		RG_rl_95_t1 = TR_107 ;
	7'h0c :
		RG_rl_95_t1 = TR_107 ;
	7'h0d :
		RG_rl_95_t1 = TR_107 ;
	7'h0e :
		RG_rl_95_t1 = TR_107 ;
	7'h0f :
		RG_rl_95_t1 = TR_107 ;
	7'h10 :
		RG_rl_95_t1 = TR_107 ;
	7'h11 :
		RG_rl_95_t1 = TR_107 ;
	7'h12 :
		RG_rl_95_t1 = TR_107 ;
	7'h13 :
		RG_rl_95_t1 = TR_107 ;
	7'h14 :
		RG_rl_95_t1 = TR_107 ;
	7'h15 :
		RG_rl_95_t1 = TR_107 ;
	7'h16 :
		RG_rl_95_t1 = TR_107 ;
	7'h17 :
		RG_rl_95_t1 = TR_107 ;
	7'h18 :
		RG_rl_95_t1 = TR_107 ;
	7'h19 :
		RG_rl_95_t1 = TR_107 ;
	7'h1a :
		RG_rl_95_t1 = TR_107 ;
	7'h1b :
		RG_rl_95_t1 = TR_107 ;
	7'h1c :
		RG_rl_95_t1 = TR_107 ;
	7'h1d :
		RG_rl_95_t1 = TR_107 ;
	7'h1e :
		RG_rl_95_t1 = TR_107 ;
	7'h1f :
		RG_rl_95_t1 = TR_107 ;
	7'h20 :
		RG_rl_95_t1 = TR_107 ;
	7'h21 :
		RG_rl_95_t1 = TR_107 ;
	7'h22 :
		RG_rl_95_t1 = TR_107 ;
	7'h23 :
		RG_rl_95_t1 = TR_107 ;
	7'h24 :
		RG_rl_95_t1 = TR_107 ;
	7'h25 :
		RG_rl_95_t1 = TR_107 ;
	7'h26 :
		RG_rl_95_t1 = TR_107 ;
	7'h27 :
		RG_rl_95_t1 = TR_107 ;
	7'h28 :
		RG_rl_95_t1 = TR_107 ;
	7'h29 :
		RG_rl_95_t1 = TR_107 ;
	7'h2a :
		RG_rl_95_t1 = TR_107 ;
	7'h2b :
		RG_rl_95_t1 = TR_107 ;
	7'h2c :
		RG_rl_95_t1 = TR_107 ;
	7'h2d :
		RG_rl_95_t1 = TR_107 ;
	7'h2e :
		RG_rl_95_t1 = TR_107 ;
	7'h2f :
		RG_rl_95_t1 = TR_107 ;
	7'h30 :
		RG_rl_95_t1 = TR_107 ;
	7'h31 :
		RG_rl_95_t1 = TR_107 ;
	7'h32 :
		RG_rl_95_t1 = TR_107 ;
	7'h33 :
		RG_rl_95_t1 = TR_107 ;
	7'h34 :
		RG_rl_95_t1 = TR_107 ;
	7'h35 :
		RG_rl_95_t1 = TR_107 ;
	7'h36 :
		RG_rl_95_t1 = TR_107 ;
	7'h37 :
		RG_rl_95_t1 = TR_107 ;
	7'h38 :
		RG_rl_95_t1 = TR_107 ;
	7'h39 :
		RG_rl_95_t1 = TR_107 ;
	7'h3a :
		RG_rl_95_t1 = TR_107 ;
	7'h3b :
		RG_rl_95_t1 = TR_107 ;
	7'h3c :
		RG_rl_95_t1 = TR_107 ;
	7'h3d :
		RG_rl_95_t1 = TR_107 ;
	7'h3e :
		RG_rl_95_t1 = TR_107 ;
	7'h3f :
		RG_rl_95_t1 = TR_107 ;
	7'h40 :
		RG_rl_95_t1 = TR_107 ;
	7'h41 :
		RG_rl_95_t1 = TR_107 ;
	7'h42 :
		RG_rl_95_t1 = TR_107 ;
	7'h43 :
		RG_rl_95_t1 = TR_107 ;
	7'h44 :
		RG_rl_95_t1 = TR_107 ;
	7'h45 :
		RG_rl_95_t1 = TR_107 ;
	7'h46 :
		RG_rl_95_t1 = TR_107 ;
	7'h47 :
		RG_rl_95_t1 = TR_107 ;
	7'h48 :
		RG_rl_95_t1 = TR_107 ;
	7'h49 :
		RG_rl_95_t1 = TR_107 ;
	7'h4a :
		RG_rl_95_t1 = TR_107 ;
	7'h4b :
		RG_rl_95_t1 = TR_107 ;
	7'h4c :
		RG_rl_95_t1 = TR_107 ;
	7'h4d :
		RG_rl_95_t1 = TR_107 ;
	7'h4e :
		RG_rl_95_t1 = TR_107 ;
	7'h4f :
		RG_rl_95_t1 = TR_107 ;
	7'h50 :
		RG_rl_95_t1 = TR_107 ;
	7'h51 :
		RG_rl_95_t1 = TR_107 ;
	7'h52 :
		RG_rl_95_t1 = TR_107 ;
	7'h53 :
		RG_rl_95_t1 = TR_107 ;
	7'h54 :
		RG_rl_95_t1 = TR_107 ;
	7'h55 :
		RG_rl_95_t1 = TR_107 ;
	7'h56 :
		RG_rl_95_t1 = TR_107 ;
	7'h57 :
		RG_rl_95_t1 = TR_107 ;
	7'h58 :
		RG_rl_95_t1 = TR_107 ;
	7'h59 :
		RG_rl_95_t1 = TR_107 ;
	7'h5a :
		RG_rl_95_t1 = TR_107 ;
	7'h5b :
		RG_rl_95_t1 = TR_107 ;
	7'h5c :
		RG_rl_95_t1 = TR_107 ;
	7'h5d :
		RG_rl_95_t1 = TR_107 ;
	7'h5e :
		RG_rl_95_t1 = TR_107 ;
	7'h5f :
		RG_rl_95_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h60 :
		RG_rl_95_t1 = TR_107 ;
	7'h61 :
		RG_rl_95_t1 = TR_107 ;
	7'h62 :
		RG_rl_95_t1 = TR_107 ;
	7'h63 :
		RG_rl_95_t1 = TR_107 ;
	7'h64 :
		RG_rl_95_t1 = TR_107 ;
	7'h65 :
		RG_rl_95_t1 = TR_107 ;
	7'h66 :
		RG_rl_95_t1 = TR_107 ;
	7'h67 :
		RG_rl_95_t1 = TR_107 ;
	7'h68 :
		RG_rl_95_t1 = TR_107 ;
	7'h69 :
		RG_rl_95_t1 = TR_107 ;
	7'h6a :
		RG_rl_95_t1 = TR_107 ;
	7'h6b :
		RG_rl_95_t1 = TR_107 ;
	7'h6c :
		RG_rl_95_t1 = TR_107 ;
	7'h6d :
		RG_rl_95_t1 = TR_107 ;
	7'h6e :
		RG_rl_95_t1 = TR_107 ;
	7'h6f :
		RG_rl_95_t1 = TR_107 ;
	7'h70 :
		RG_rl_95_t1 = TR_107 ;
	7'h71 :
		RG_rl_95_t1 = TR_107 ;
	7'h72 :
		RG_rl_95_t1 = TR_107 ;
	7'h73 :
		RG_rl_95_t1 = TR_107 ;
	7'h74 :
		RG_rl_95_t1 = TR_107 ;
	7'h75 :
		RG_rl_95_t1 = TR_107 ;
	7'h76 :
		RG_rl_95_t1 = TR_107 ;
	7'h77 :
		RG_rl_95_t1 = TR_107 ;
	7'h78 :
		RG_rl_95_t1 = TR_107 ;
	7'h79 :
		RG_rl_95_t1 = TR_107 ;
	7'h7a :
		RG_rl_95_t1 = TR_107 ;
	7'h7b :
		RG_rl_95_t1 = TR_107 ;
	7'h7c :
		RG_rl_95_t1 = TR_107 ;
	7'h7d :
		RG_rl_95_t1 = TR_107 ;
	7'h7e :
		RG_rl_95_t1 = TR_107 ;
	7'h7f :
		RG_rl_95_t1 = TR_107 ;
	default :
		RG_rl_95_t1 = 9'hx ;
	endcase
always @ ( RG_rl_95_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_36 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_95_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h5f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_95_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_36 )
		| ( { 9{ U_569 } } & RG_rl_95_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_95_en = ( U_570 | RG_rl_95_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_95_en )
		RG_rl_95 <= RG_rl_95_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_108 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_96_t1 = TR_108 ;
	7'h01 :
		RG_rl_96_t1 = TR_108 ;
	7'h02 :
		RG_rl_96_t1 = TR_108 ;
	7'h03 :
		RG_rl_96_t1 = TR_108 ;
	7'h04 :
		RG_rl_96_t1 = TR_108 ;
	7'h05 :
		RG_rl_96_t1 = TR_108 ;
	7'h06 :
		RG_rl_96_t1 = TR_108 ;
	7'h07 :
		RG_rl_96_t1 = TR_108 ;
	7'h08 :
		RG_rl_96_t1 = TR_108 ;
	7'h09 :
		RG_rl_96_t1 = TR_108 ;
	7'h0a :
		RG_rl_96_t1 = TR_108 ;
	7'h0b :
		RG_rl_96_t1 = TR_108 ;
	7'h0c :
		RG_rl_96_t1 = TR_108 ;
	7'h0d :
		RG_rl_96_t1 = TR_108 ;
	7'h0e :
		RG_rl_96_t1 = TR_108 ;
	7'h0f :
		RG_rl_96_t1 = TR_108 ;
	7'h10 :
		RG_rl_96_t1 = TR_108 ;
	7'h11 :
		RG_rl_96_t1 = TR_108 ;
	7'h12 :
		RG_rl_96_t1 = TR_108 ;
	7'h13 :
		RG_rl_96_t1 = TR_108 ;
	7'h14 :
		RG_rl_96_t1 = TR_108 ;
	7'h15 :
		RG_rl_96_t1 = TR_108 ;
	7'h16 :
		RG_rl_96_t1 = TR_108 ;
	7'h17 :
		RG_rl_96_t1 = TR_108 ;
	7'h18 :
		RG_rl_96_t1 = TR_108 ;
	7'h19 :
		RG_rl_96_t1 = TR_108 ;
	7'h1a :
		RG_rl_96_t1 = TR_108 ;
	7'h1b :
		RG_rl_96_t1 = TR_108 ;
	7'h1c :
		RG_rl_96_t1 = TR_108 ;
	7'h1d :
		RG_rl_96_t1 = TR_108 ;
	7'h1e :
		RG_rl_96_t1 = TR_108 ;
	7'h1f :
		RG_rl_96_t1 = TR_108 ;
	7'h20 :
		RG_rl_96_t1 = TR_108 ;
	7'h21 :
		RG_rl_96_t1 = TR_108 ;
	7'h22 :
		RG_rl_96_t1 = TR_108 ;
	7'h23 :
		RG_rl_96_t1 = TR_108 ;
	7'h24 :
		RG_rl_96_t1 = TR_108 ;
	7'h25 :
		RG_rl_96_t1 = TR_108 ;
	7'h26 :
		RG_rl_96_t1 = TR_108 ;
	7'h27 :
		RG_rl_96_t1 = TR_108 ;
	7'h28 :
		RG_rl_96_t1 = TR_108 ;
	7'h29 :
		RG_rl_96_t1 = TR_108 ;
	7'h2a :
		RG_rl_96_t1 = TR_108 ;
	7'h2b :
		RG_rl_96_t1 = TR_108 ;
	7'h2c :
		RG_rl_96_t1 = TR_108 ;
	7'h2d :
		RG_rl_96_t1 = TR_108 ;
	7'h2e :
		RG_rl_96_t1 = TR_108 ;
	7'h2f :
		RG_rl_96_t1 = TR_108 ;
	7'h30 :
		RG_rl_96_t1 = TR_108 ;
	7'h31 :
		RG_rl_96_t1 = TR_108 ;
	7'h32 :
		RG_rl_96_t1 = TR_108 ;
	7'h33 :
		RG_rl_96_t1 = TR_108 ;
	7'h34 :
		RG_rl_96_t1 = TR_108 ;
	7'h35 :
		RG_rl_96_t1 = TR_108 ;
	7'h36 :
		RG_rl_96_t1 = TR_108 ;
	7'h37 :
		RG_rl_96_t1 = TR_108 ;
	7'h38 :
		RG_rl_96_t1 = TR_108 ;
	7'h39 :
		RG_rl_96_t1 = TR_108 ;
	7'h3a :
		RG_rl_96_t1 = TR_108 ;
	7'h3b :
		RG_rl_96_t1 = TR_108 ;
	7'h3c :
		RG_rl_96_t1 = TR_108 ;
	7'h3d :
		RG_rl_96_t1 = TR_108 ;
	7'h3e :
		RG_rl_96_t1 = TR_108 ;
	7'h3f :
		RG_rl_96_t1 = TR_108 ;
	7'h40 :
		RG_rl_96_t1 = TR_108 ;
	7'h41 :
		RG_rl_96_t1 = TR_108 ;
	7'h42 :
		RG_rl_96_t1 = TR_108 ;
	7'h43 :
		RG_rl_96_t1 = TR_108 ;
	7'h44 :
		RG_rl_96_t1 = TR_108 ;
	7'h45 :
		RG_rl_96_t1 = TR_108 ;
	7'h46 :
		RG_rl_96_t1 = TR_108 ;
	7'h47 :
		RG_rl_96_t1 = TR_108 ;
	7'h48 :
		RG_rl_96_t1 = TR_108 ;
	7'h49 :
		RG_rl_96_t1 = TR_108 ;
	7'h4a :
		RG_rl_96_t1 = TR_108 ;
	7'h4b :
		RG_rl_96_t1 = TR_108 ;
	7'h4c :
		RG_rl_96_t1 = TR_108 ;
	7'h4d :
		RG_rl_96_t1 = TR_108 ;
	7'h4e :
		RG_rl_96_t1 = TR_108 ;
	7'h4f :
		RG_rl_96_t1 = TR_108 ;
	7'h50 :
		RG_rl_96_t1 = TR_108 ;
	7'h51 :
		RG_rl_96_t1 = TR_108 ;
	7'h52 :
		RG_rl_96_t1 = TR_108 ;
	7'h53 :
		RG_rl_96_t1 = TR_108 ;
	7'h54 :
		RG_rl_96_t1 = TR_108 ;
	7'h55 :
		RG_rl_96_t1 = TR_108 ;
	7'h56 :
		RG_rl_96_t1 = TR_108 ;
	7'h57 :
		RG_rl_96_t1 = TR_108 ;
	7'h58 :
		RG_rl_96_t1 = TR_108 ;
	7'h59 :
		RG_rl_96_t1 = TR_108 ;
	7'h5a :
		RG_rl_96_t1 = TR_108 ;
	7'h5b :
		RG_rl_96_t1 = TR_108 ;
	7'h5c :
		RG_rl_96_t1 = TR_108 ;
	7'h5d :
		RG_rl_96_t1 = TR_108 ;
	7'h5e :
		RG_rl_96_t1 = TR_108 ;
	7'h5f :
		RG_rl_96_t1 = TR_108 ;
	7'h60 :
		RG_rl_96_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h61 :
		RG_rl_96_t1 = TR_108 ;
	7'h62 :
		RG_rl_96_t1 = TR_108 ;
	7'h63 :
		RG_rl_96_t1 = TR_108 ;
	7'h64 :
		RG_rl_96_t1 = TR_108 ;
	7'h65 :
		RG_rl_96_t1 = TR_108 ;
	7'h66 :
		RG_rl_96_t1 = TR_108 ;
	7'h67 :
		RG_rl_96_t1 = TR_108 ;
	7'h68 :
		RG_rl_96_t1 = TR_108 ;
	7'h69 :
		RG_rl_96_t1 = TR_108 ;
	7'h6a :
		RG_rl_96_t1 = TR_108 ;
	7'h6b :
		RG_rl_96_t1 = TR_108 ;
	7'h6c :
		RG_rl_96_t1 = TR_108 ;
	7'h6d :
		RG_rl_96_t1 = TR_108 ;
	7'h6e :
		RG_rl_96_t1 = TR_108 ;
	7'h6f :
		RG_rl_96_t1 = TR_108 ;
	7'h70 :
		RG_rl_96_t1 = TR_108 ;
	7'h71 :
		RG_rl_96_t1 = TR_108 ;
	7'h72 :
		RG_rl_96_t1 = TR_108 ;
	7'h73 :
		RG_rl_96_t1 = TR_108 ;
	7'h74 :
		RG_rl_96_t1 = TR_108 ;
	7'h75 :
		RG_rl_96_t1 = TR_108 ;
	7'h76 :
		RG_rl_96_t1 = TR_108 ;
	7'h77 :
		RG_rl_96_t1 = TR_108 ;
	7'h78 :
		RG_rl_96_t1 = TR_108 ;
	7'h79 :
		RG_rl_96_t1 = TR_108 ;
	7'h7a :
		RG_rl_96_t1 = TR_108 ;
	7'h7b :
		RG_rl_96_t1 = TR_108 ;
	7'h7c :
		RG_rl_96_t1 = TR_108 ;
	7'h7d :
		RG_rl_96_t1 = TR_108 ;
	7'h7e :
		RG_rl_96_t1 = TR_108 ;
	7'h7f :
		RG_rl_96_t1 = TR_108 ;
	default :
		RG_rl_96_t1 = 9'hx ;
	endcase
always @ ( RG_rl_96_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_37 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_96_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h60 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_96_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_37 )
		| ( { 9{ U_569 } } & RG_rl_96_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_96_en = ( U_570 | RG_rl_96_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_96_en )
		RG_rl_96 <= RG_rl_96_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_109 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_97_t1 = TR_109 ;
	7'h01 :
		RG_rl_97_t1 = TR_109 ;
	7'h02 :
		RG_rl_97_t1 = TR_109 ;
	7'h03 :
		RG_rl_97_t1 = TR_109 ;
	7'h04 :
		RG_rl_97_t1 = TR_109 ;
	7'h05 :
		RG_rl_97_t1 = TR_109 ;
	7'h06 :
		RG_rl_97_t1 = TR_109 ;
	7'h07 :
		RG_rl_97_t1 = TR_109 ;
	7'h08 :
		RG_rl_97_t1 = TR_109 ;
	7'h09 :
		RG_rl_97_t1 = TR_109 ;
	7'h0a :
		RG_rl_97_t1 = TR_109 ;
	7'h0b :
		RG_rl_97_t1 = TR_109 ;
	7'h0c :
		RG_rl_97_t1 = TR_109 ;
	7'h0d :
		RG_rl_97_t1 = TR_109 ;
	7'h0e :
		RG_rl_97_t1 = TR_109 ;
	7'h0f :
		RG_rl_97_t1 = TR_109 ;
	7'h10 :
		RG_rl_97_t1 = TR_109 ;
	7'h11 :
		RG_rl_97_t1 = TR_109 ;
	7'h12 :
		RG_rl_97_t1 = TR_109 ;
	7'h13 :
		RG_rl_97_t1 = TR_109 ;
	7'h14 :
		RG_rl_97_t1 = TR_109 ;
	7'h15 :
		RG_rl_97_t1 = TR_109 ;
	7'h16 :
		RG_rl_97_t1 = TR_109 ;
	7'h17 :
		RG_rl_97_t1 = TR_109 ;
	7'h18 :
		RG_rl_97_t1 = TR_109 ;
	7'h19 :
		RG_rl_97_t1 = TR_109 ;
	7'h1a :
		RG_rl_97_t1 = TR_109 ;
	7'h1b :
		RG_rl_97_t1 = TR_109 ;
	7'h1c :
		RG_rl_97_t1 = TR_109 ;
	7'h1d :
		RG_rl_97_t1 = TR_109 ;
	7'h1e :
		RG_rl_97_t1 = TR_109 ;
	7'h1f :
		RG_rl_97_t1 = TR_109 ;
	7'h20 :
		RG_rl_97_t1 = TR_109 ;
	7'h21 :
		RG_rl_97_t1 = TR_109 ;
	7'h22 :
		RG_rl_97_t1 = TR_109 ;
	7'h23 :
		RG_rl_97_t1 = TR_109 ;
	7'h24 :
		RG_rl_97_t1 = TR_109 ;
	7'h25 :
		RG_rl_97_t1 = TR_109 ;
	7'h26 :
		RG_rl_97_t1 = TR_109 ;
	7'h27 :
		RG_rl_97_t1 = TR_109 ;
	7'h28 :
		RG_rl_97_t1 = TR_109 ;
	7'h29 :
		RG_rl_97_t1 = TR_109 ;
	7'h2a :
		RG_rl_97_t1 = TR_109 ;
	7'h2b :
		RG_rl_97_t1 = TR_109 ;
	7'h2c :
		RG_rl_97_t1 = TR_109 ;
	7'h2d :
		RG_rl_97_t1 = TR_109 ;
	7'h2e :
		RG_rl_97_t1 = TR_109 ;
	7'h2f :
		RG_rl_97_t1 = TR_109 ;
	7'h30 :
		RG_rl_97_t1 = TR_109 ;
	7'h31 :
		RG_rl_97_t1 = TR_109 ;
	7'h32 :
		RG_rl_97_t1 = TR_109 ;
	7'h33 :
		RG_rl_97_t1 = TR_109 ;
	7'h34 :
		RG_rl_97_t1 = TR_109 ;
	7'h35 :
		RG_rl_97_t1 = TR_109 ;
	7'h36 :
		RG_rl_97_t1 = TR_109 ;
	7'h37 :
		RG_rl_97_t1 = TR_109 ;
	7'h38 :
		RG_rl_97_t1 = TR_109 ;
	7'h39 :
		RG_rl_97_t1 = TR_109 ;
	7'h3a :
		RG_rl_97_t1 = TR_109 ;
	7'h3b :
		RG_rl_97_t1 = TR_109 ;
	7'h3c :
		RG_rl_97_t1 = TR_109 ;
	7'h3d :
		RG_rl_97_t1 = TR_109 ;
	7'h3e :
		RG_rl_97_t1 = TR_109 ;
	7'h3f :
		RG_rl_97_t1 = TR_109 ;
	7'h40 :
		RG_rl_97_t1 = TR_109 ;
	7'h41 :
		RG_rl_97_t1 = TR_109 ;
	7'h42 :
		RG_rl_97_t1 = TR_109 ;
	7'h43 :
		RG_rl_97_t1 = TR_109 ;
	7'h44 :
		RG_rl_97_t1 = TR_109 ;
	7'h45 :
		RG_rl_97_t1 = TR_109 ;
	7'h46 :
		RG_rl_97_t1 = TR_109 ;
	7'h47 :
		RG_rl_97_t1 = TR_109 ;
	7'h48 :
		RG_rl_97_t1 = TR_109 ;
	7'h49 :
		RG_rl_97_t1 = TR_109 ;
	7'h4a :
		RG_rl_97_t1 = TR_109 ;
	7'h4b :
		RG_rl_97_t1 = TR_109 ;
	7'h4c :
		RG_rl_97_t1 = TR_109 ;
	7'h4d :
		RG_rl_97_t1 = TR_109 ;
	7'h4e :
		RG_rl_97_t1 = TR_109 ;
	7'h4f :
		RG_rl_97_t1 = TR_109 ;
	7'h50 :
		RG_rl_97_t1 = TR_109 ;
	7'h51 :
		RG_rl_97_t1 = TR_109 ;
	7'h52 :
		RG_rl_97_t1 = TR_109 ;
	7'h53 :
		RG_rl_97_t1 = TR_109 ;
	7'h54 :
		RG_rl_97_t1 = TR_109 ;
	7'h55 :
		RG_rl_97_t1 = TR_109 ;
	7'h56 :
		RG_rl_97_t1 = TR_109 ;
	7'h57 :
		RG_rl_97_t1 = TR_109 ;
	7'h58 :
		RG_rl_97_t1 = TR_109 ;
	7'h59 :
		RG_rl_97_t1 = TR_109 ;
	7'h5a :
		RG_rl_97_t1 = TR_109 ;
	7'h5b :
		RG_rl_97_t1 = TR_109 ;
	7'h5c :
		RG_rl_97_t1 = TR_109 ;
	7'h5d :
		RG_rl_97_t1 = TR_109 ;
	7'h5e :
		RG_rl_97_t1 = TR_109 ;
	7'h5f :
		RG_rl_97_t1 = TR_109 ;
	7'h60 :
		RG_rl_97_t1 = TR_109 ;
	7'h61 :
		RG_rl_97_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h62 :
		RG_rl_97_t1 = TR_109 ;
	7'h63 :
		RG_rl_97_t1 = TR_109 ;
	7'h64 :
		RG_rl_97_t1 = TR_109 ;
	7'h65 :
		RG_rl_97_t1 = TR_109 ;
	7'h66 :
		RG_rl_97_t1 = TR_109 ;
	7'h67 :
		RG_rl_97_t1 = TR_109 ;
	7'h68 :
		RG_rl_97_t1 = TR_109 ;
	7'h69 :
		RG_rl_97_t1 = TR_109 ;
	7'h6a :
		RG_rl_97_t1 = TR_109 ;
	7'h6b :
		RG_rl_97_t1 = TR_109 ;
	7'h6c :
		RG_rl_97_t1 = TR_109 ;
	7'h6d :
		RG_rl_97_t1 = TR_109 ;
	7'h6e :
		RG_rl_97_t1 = TR_109 ;
	7'h6f :
		RG_rl_97_t1 = TR_109 ;
	7'h70 :
		RG_rl_97_t1 = TR_109 ;
	7'h71 :
		RG_rl_97_t1 = TR_109 ;
	7'h72 :
		RG_rl_97_t1 = TR_109 ;
	7'h73 :
		RG_rl_97_t1 = TR_109 ;
	7'h74 :
		RG_rl_97_t1 = TR_109 ;
	7'h75 :
		RG_rl_97_t1 = TR_109 ;
	7'h76 :
		RG_rl_97_t1 = TR_109 ;
	7'h77 :
		RG_rl_97_t1 = TR_109 ;
	7'h78 :
		RG_rl_97_t1 = TR_109 ;
	7'h79 :
		RG_rl_97_t1 = TR_109 ;
	7'h7a :
		RG_rl_97_t1 = TR_109 ;
	7'h7b :
		RG_rl_97_t1 = TR_109 ;
	7'h7c :
		RG_rl_97_t1 = TR_109 ;
	7'h7d :
		RG_rl_97_t1 = TR_109 ;
	7'h7e :
		RG_rl_97_t1 = TR_109 ;
	7'h7f :
		RG_rl_97_t1 = TR_109 ;
	default :
		RG_rl_97_t1 = 9'hx ;
	endcase
always @ ( RG_rl_97_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_38 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_97_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h61 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_97_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_38 )
		| ( { 9{ U_569 } } & RG_rl_97_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_97_en = ( U_570 | RG_rl_97_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_97_en )
		RG_rl_97 <= RG_rl_97_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_110 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_98_t1 = TR_110 ;
	7'h01 :
		RG_rl_98_t1 = TR_110 ;
	7'h02 :
		RG_rl_98_t1 = TR_110 ;
	7'h03 :
		RG_rl_98_t1 = TR_110 ;
	7'h04 :
		RG_rl_98_t1 = TR_110 ;
	7'h05 :
		RG_rl_98_t1 = TR_110 ;
	7'h06 :
		RG_rl_98_t1 = TR_110 ;
	7'h07 :
		RG_rl_98_t1 = TR_110 ;
	7'h08 :
		RG_rl_98_t1 = TR_110 ;
	7'h09 :
		RG_rl_98_t1 = TR_110 ;
	7'h0a :
		RG_rl_98_t1 = TR_110 ;
	7'h0b :
		RG_rl_98_t1 = TR_110 ;
	7'h0c :
		RG_rl_98_t1 = TR_110 ;
	7'h0d :
		RG_rl_98_t1 = TR_110 ;
	7'h0e :
		RG_rl_98_t1 = TR_110 ;
	7'h0f :
		RG_rl_98_t1 = TR_110 ;
	7'h10 :
		RG_rl_98_t1 = TR_110 ;
	7'h11 :
		RG_rl_98_t1 = TR_110 ;
	7'h12 :
		RG_rl_98_t1 = TR_110 ;
	7'h13 :
		RG_rl_98_t1 = TR_110 ;
	7'h14 :
		RG_rl_98_t1 = TR_110 ;
	7'h15 :
		RG_rl_98_t1 = TR_110 ;
	7'h16 :
		RG_rl_98_t1 = TR_110 ;
	7'h17 :
		RG_rl_98_t1 = TR_110 ;
	7'h18 :
		RG_rl_98_t1 = TR_110 ;
	7'h19 :
		RG_rl_98_t1 = TR_110 ;
	7'h1a :
		RG_rl_98_t1 = TR_110 ;
	7'h1b :
		RG_rl_98_t1 = TR_110 ;
	7'h1c :
		RG_rl_98_t1 = TR_110 ;
	7'h1d :
		RG_rl_98_t1 = TR_110 ;
	7'h1e :
		RG_rl_98_t1 = TR_110 ;
	7'h1f :
		RG_rl_98_t1 = TR_110 ;
	7'h20 :
		RG_rl_98_t1 = TR_110 ;
	7'h21 :
		RG_rl_98_t1 = TR_110 ;
	7'h22 :
		RG_rl_98_t1 = TR_110 ;
	7'h23 :
		RG_rl_98_t1 = TR_110 ;
	7'h24 :
		RG_rl_98_t1 = TR_110 ;
	7'h25 :
		RG_rl_98_t1 = TR_110 ;
	7'h26 :
		RG_rl_98_t1 = TR_110 ;
	7'h27 :
		RG_rl_98_t1 = TR_110 ;
	7'h28 :
		RG_rl_98_t1 = TR_110 ;
	7'h29 :
		RG_rl_98_t1 = TR_110 ;
	7'h2a :
		RG_rl_98_t1 = TR_110 ;
	7'h2b :
		RG_rl_98_t1 = TR_110 ;
	7'h2c :
		RG_rl_98_t1 = TR_110 ;
	7'h2d :
		RG_rl_98_t1 = TR_110 ;
	7'h2e :
		RG_rl_98_t1 = TR_110 ;
	7'h2f :
		RG_rl_98_t1 = TR_110 ;
	7'h30 :
		RG_rl_98_t1 = TR_110 ;
	7'h31 :
		RG_rl_98_t1 = TR_110 ;
	7'h32 :
		RG_rl_98_t1 = TR_110 ;
	7'h33 :
		RG_rl_98_t1 = TR_110 ;
	7'h34 :
		RG_rl_98_t1 = TR_110 ;
	7'h35 :
		RG_rl_98_t1 = TR_110 ;
	7'h36 :
		RG_rl_98_t1 = TR_110 ;
	7'h37 :
		RG_rl_98_t1 = TR_110 ;
	7'h38 :
		RG_rl_98_t1 = TR_110 ;
	7'h39 :
		RG_rl_98_t1 = TR_110 ;
	7'h3a :
		RG_rl_98_t1 = TR_110 ;
	7'h3b :
		RG_rl_98_t1 = TR_110 ;
	7'h3c :
		RG_rl_98_t1 = TR_110 ;
	7'h3d :
		RG_rl_98_t1 = TR_110 ;
	7'h3e :
		RG_rl_98_t1 = TR_110 ;
	7'h3f :
		RG_rl_98_t1 = TR_110 ;
	7'h40 :
		RG_rl_98_t1 = TR_110 ;
	7'h41 :
		RG_rl_98_t1 = TR_110 ;
	7'h42 :
		RG_rl_98_t1 = TR_110 ;
	7'h43 :
		RG_rl_98_t1 = TR_110 ;
	7'h44 :
		RG_rl_98_t1 = TR_110 ;
	7'h45 :
		RG_rl_98_t1 = TR_110 ;
	7'h46 :
		RG_rl_98_t1 = TR_110 ;
	7'h47 :
		RG_rl_98_t1 = TR_110 ;
	7'h48 :
		RG_rl_98_t1 = TR_110 ;
	7'h49 :
		RG_rl_98_t1 = TR_110 ;
	7'h4a :
		RG_rl_98_t1 = TR_110 ;
	7'h4b :
		RG_rl_98_t1 = TR_110 ;
	7'h4c :
		RG_rl_98_t1 = TR_110 ;
	7'h4d :
		RG_rl_98_t1 = TR_110 ;
	7'h4e :
		RG_rl_98_t1 = TR_110 ;
	7'h4f :
		RG_rl_98_t1 = TR_110 ;
	7'h50 :
		RG_rl_98_t1 = TR_110 ;
	7'h51 :
		RG_rl_98_t1 = TR_110 ;
	7'h52 :
		RG_rl_98_t1 = TR_110 ;
	7'h53 :
		RG_rl_98_t1 = TR_110 ;
	7'h54 :
		RG_rl_98_t1 = TR_110 ;
	7'h55 :
		RG_rl_98_t1 = TR_110 ;
	7'h56 :
		RG_rl_98_t1 = TR_110 ;
	7'h57 :
		RG_rl_98_t1 = TR_110 ;
	7'h58 :
		RG_rl_98_t1 = TR_110 ;
	7'h59 :
		RG_rl_98_t1 = TR_110 ;
	7'h5a :
		RG_rl_98_t1 = TR_110 ;
	7'h5b :
		RG_rl_98_t1 = TR_110 ;
	7'h5c :
		RG_rl_98_t1 = TR_110 ;
	7'h5d :
		RG_rl_98_t1 = TR_110 ;
	7'h5e :
		RG_rl_98_t1 = TR_110 ;
	7'h5f :
		RG_rl_98_t1 = TR_110 ;
	7'h60 :
		RG_rl_98_t1 = TR_110 ;
	7'h61 :
		RG_rl_98_t1 = TR_110 ;
	7'h62 :
		RG_rl_98_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h63 :
		RG_rl_98_t1 = TR_110 ;
	7'h64 :
		RG_rl_98_t1 = TR_110 ;
	7'h65 :
		RG_rl_98_t1 = TR_110 ;
	7'h66 :
		RG_rl_98_t1 = TR_110 ;
	7'h67 :
		RG_rl_98_t1 = TR_110 ;
	7'h68 :
		RG_rl_98_t1 = TR_110 ;
	7'h69 :
		RG_rl_98_t1 = TR_110 ;
	7'h6a :
		RG_rl_98_t1 = TR_110 ;
	7'h6b :
		RG_rl_98_t1 = TR_110 ;
	7'h6c :
		RG_rl_98_t1 = TR_110 ;
	7'h6d :
		RG_rl_98_t1 = TR_110 ;
	7'h6e :
		RG_rl_98_t1 = TR_110 ;
	7'h6f :
		RG_rl_98_t1 = TR_110 ;
	7'h70 :
		RG_rl_98_t1 = TR_110 ;
	7'h71 :
		RG_rl_98_t1 = TR_110 ;
	7'h72 :
		RG_rl_98_t1 = TR_110 ;
	7'h73 :
		RG_rl_98_t1 = TR_110 ;
	7'h74 :
		RG_rl_98_t1 = TR_110 ;
	7'h75 :
		RG_rl_98_t1 = TR_110 ;
	7'h76 :
		RG_rl_98_t1 = TR_110 ;
	7'h77 :
		RG_rl_98_t1 = TR_110 ;
	7'h78 :
		RG_rl_98_t1 = TR_110 ;
	7'h79 :
		RG_rl_98_t1 = TR_110 ;
	7'h7a :
		RG_rl_98_t1 = TR_110 ;
	7'h7b :
		RG_rl_98_t1 = TR_110 ;
	7'h7c :
		RG_rl_98_t1 = TR_110 ;
	7'h7d :
		RG_rl_98_t1 = TR_110 ;
	7'h7e :
		RG_rl_98_t1 = TR_110 ;
	7'h7f :
		RG_rl_98_t1 = TR_110 ;
	default :
		RG_rl_98_t1 = 9'hx ;
	endcase
always @ ( RG_rl_98_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_39 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_98_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h62 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_98_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_39 )
		| ( { 9{ U_569 } } & RG_rl_98_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_98_en = ( U_570 | RG_rl_98_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_98_en )
		RG_rl_98 <= RG_rl_98_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_111 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_99_t1 = TR_111 ;
	7'h01 :
		RG_rl_99_t1 = TR_111 ;
	7'h02 :
		RG_rl_99_t1 = TR_111 ;
	7'h03 :
		RG_rl_99_t1 = TR_111 ;
	7'h04 :
		RG_rl_99_t1 = TR_111 ;
	7'h05 :
		RG_rl_99_t1 = TR_111 ;
	7'h06 :
		RG_rl_99_t1 = TR_111 ;
	7'h07 :
		RG_rl_99_t1 = TR_111 ;
	7'h08 :
		RG_rl_99_t1 = TR_111 ;
	7'h09 :
		RG_rl_99_t1 = TR_111 ;
	7'h0a :
		RG_rl_99_t1 = TR_111 ;
	7'h0b :
		RG_rl_99_t1 = TR_111 ;
	7'h0c :
		RG_rl_99_t1 = TR_111 ;
	7'h0d :
		RG_rl_99_t1 = TR_111 ;
	7'h0e :
		RG_rl_99_t1 = TR_111 ;
	7'h0f :
		RG_rl_99_t1 = TR_111 ;
	7'h10 :
		RG_rl_99_t1 = TR_111 ;
	7'h11 :
		RG_rl_99_t1 = TR_111 ;
	7'h12 :
		RG_rl_99_t1 = TR_111 ;
	7'h13 :
		RG_rl_99_t1 = TR_111 ;
	7'h14 :
		RG_rl_99_t1 = TR_111 ;
	7'h15 :
		RG_rl_99_t1 = TR_111 ;
	7'h16 :
		RG_rl_99_t1 = TR_111 ;
	7'h17 :
		RG_rl_99_t1 = TR_111 ;
	7'h18 :
		RG_rl_99_t1 = TR_111 ;
	7'h19 :
		RG_rl_99_t1 = TR_111 ;
	7'h1a :
		RG_rl_99_t1 = TR_111 ;
	7'h1b :
		RG_rl_99_t1 = TR_111 ;
	7'h1c :
		RG_rl_99_t1 = TR_111 ;
	7'h1d :
		RG_rl_99_t1 = TR_111 ;
	7'h1e :
		RG_rl_99_t1 = TR_111 ;
	7'h1f :
		RG_rl_99_t1 = TR_111 ;
	7'h20 :
		RG_rl_99_t1 = TR_111 ;
	7'h21 :
		RG_rl_99_t1 = TR_111 ;
	7'h22 :
		RG_rl_99_t1 = TR_111 ;
	7'h23 :
		RG_rl_99_t1 = TR_111 ;
	7'h24 :
		RG_rl_99_t1 = TR_111 ;
	7'h25 :
		RG_rl_99_t1 = TR_111 ;
	7'h26 :
		RG_rl_99_t1 = TR_111 ;
	7'h27 :
		RG_rl_99_t1 = TR_111 ;
	7'h28 :
		RG_rl_99_t1 = TR_111 ;
	7'h29 :
		RG_rl_99_t1 = TR_111 ;
	7'h2a :
		RG_rl_99_t1 = TR_111 ;
	7'h2b :
		RG_rl_99_t1 = TR_111 ;
	7'h2c :
		RG_rl_99_t1 = TR_111 ;
	7'h2d :
		RG_rl_99_t1 = TR_111 ;
	7'h2e :
		RG_rl_99_t1 = TR_111 ;
	7'h2f :
		RG_rl_99_t1 = TR_111 ;
	7'h30 :
		RG_rl_99_t1 = TR_111 ;
	7'h31 :
		RG_rl_99_t1 = TR_111 ;
	7'h32 :
		RG_rl_99_t1 = TR_111 ;
	7'h33 :
		RG_rl_99_t1 = TR_111 ;
	7'h34 :
		RG_rl_99_t1 = TR_111 ;
	7'h35 :
		RG_rl_99_t1 = TR_111 ;
	7'h36 :
		RG_rl_99_t1 = TR_111 ;
	7'h37 :
		RG_rl_99_t1 = TR_111 ;
	7'h38 :
		RG_rl_99_t1 = TR_111 ;
	7'h39 :
		RG_rl_99_t1 = TR_111 ;
	7'h3a :
		RG_rl_99_t1 = TR_111 ;
	7'h3b :
		RG_rl_99_t1 = TR_111 ;
	7'h3c :
		RG_rl_99_t1 = TR_111 ;
	7'h3d :
		RG_rl_99_t1 = TR_111 ;
	7'h3e :
		RG_rl_99_t1 = TR_111 ;
	7'h3f :
		RG_rl_99_t1 = TR_111 ;
	7'h40 :
		RG_rl_99_t1 = TR_111 ;
	7'h41 :
		RG_rl_99_t1 = TR_111 ;
	7'h42 :
		RG_rl_99_t1 = TR_111 ;
	7'h43 :
		RG_rl_99_t1 = TR_111 ;
	7'h44 :
		RG_rl_99_t1 = TR_111 ;
	7'h45 :
		RG_rl_99_t1 = TR_111 ;
	7'h46 :
		RG_rl_99_t1 = TR_111 ;
	7'h47 :
		RG_rl_99_t1 = TR_111 ;
	7'h48 :
		RG_rl_99_t1 = TR_111 ;
	7'h49 :
		RG_rl_99_t1 = TR_111 ;
	7'h4a :
		RG_rl_99_t1 = TR_111 ;
	7'h4b :
		RG_rl_99_t1 = TR_111 ;
	7'h4c :
		RG_rl_99_t1 = TR_111 ;
	7'h4d :
		RG_rl_99_t1 = TR_111 ;
	7'h4e :
		RG_rl_99_t1 = TR_111 ;
	7'h4f :
		RG_rl_99_t1 = TR_111 ;
	7'h50 :
		RG_rl_99_t1 = TR_111 ;
	7'h51 :
		RG_rl_99_t1 = TR_111 ;
	7'h52 :
		RG_rl_99_t1 = TR_111 ;
	7'h53 :
		RG_rl_99_t1 = TR_111 ;
	7'h54 :
		RG_rl_99_t1 = TR_111 ;
	7'h55 :
		RG_rl_99_t1 = TR_111 ;
	7'h56 :
		RG_rl_99_t1 = TR_111 ;
	7'h57 :
		RG_rl_99_t1 = TR_111 ;
	7'h58 :
		RG_rl_99_t1 = TR_111 ;
	7'h59 :
		RG_rl_99_t1 = TR_111 ;
	7'h5a :
		RG_rl_99_t1 = TR_111 ;
	7'h5b :
		RG_rl_99_t1 = TR_111 ;
	7'h5c :
		RG_rl_99_t1 = TR_111 ;
	7'h5d :
		RG_rl_99_t1 = TR_111 ;
	7'h5e :
		RG_rl_99_t1 = TR_111 ;
	7'h5f :
		RG_rl_99_t1 = TR_111 ;
	7'h60 :
		RG_rl_99_t1 = TR_111 ;
	7'h61 :
		RG_rl_99_t1 = TR_111 ;
	7'h62 :
		RG_rl_99_t1 = TR_111 ;
	7'h63 :
		RG_rl_99_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h64 :
		RG_rl_99_t1 = TR_111 ;
	7'h65 :
		RG_rl_99_t1 = TR_111 ;
	7'h66 :
		RG_rl_99_t1 = TR_111 ;
	7'h67 :
		RG_rl_99_t1 = TR_111 ;
	7'h68 :
		RG_rl_99_t1 = TR_111 ;
	7'h69 :
		RG_rl_99_t1 = TR_111 ;
	7'h6a :
		RG_rl_99_t1 = TR_111 ;
	7'h6b :
		RG_rl_99_t1 = TR_111 ;
	7'h6c :
		RG_rl_99_t1 = TR_111 ;
	7'h6d :
		RG_rl_99_t1 = TR_111 ;
	7'h6e :
		RG_rl_99_t1 = TR_111 ;
	7'h6f :
		RG_rl_99_t1 = TR_111 ;
	7'h70 :
		RG_rl_99_t1 = TR_111 ;
	7'h71 :
		RG_rl_99_t1 = TR_111 ;
	7'h72 :
		RG_rl_99_t1 = TR_111 ;
	7'h73 :
		RG_rl_99_t1 = TR_111 ;
	7'h74 :
		RG_rl_99_t1 = TR_111 ;
	7'h75 :
		RG_rl_99_t1 = TR_111 ;
	7'h76 :
		RG_rl_99_t1 = TR_111 ;
	7'h77 :
		RG_rl_99_t1 = TR_111 ;
	7'h78 :
		RG_rl_99_t1 = TR_111 ;
	7'h79 :
		RG_rl_99_t1 = TR_111 ;
	7'h7a :
		RG_rl_99_t1 = TR_111 ;
	7'h7b :
		RG_rl_99_t1 = TR_111 ;
	7'h7c :
		RG_rl_99_t1 = TR_111 ;
	7'h7d :
		RG_rl_99_t1 = TR_111 ;
	7'h7e :
		RG_rl_99_t1 = TR_111 ;
	7'h7f :
		RG_rl_99_t1 = TR_111 ;
	default :
		RG_rl_99_t1 = 9'hx ;
	endcase
always @ ( RG_rl_99_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_40 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_99_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h63 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_99_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_40 )
		| ( { 9{ U_569 } } & RG_rl_99_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_99_en = ( U_570 | RG_rl_99_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_99_en )
		RG_rl_99 <= RG_rl_99_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_112 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_100_t1 = TR_112 ;
	7'h01 :
		RG_rl_100_t1 = TR_112 ;
	7'h02 :
		RG_rl_100_t1 = TR_112 ;
	7'h03 :
		RG_rl_100_t1 = TR_112 ;
	7'h04 :
		RG_rl_100_t1 = TR_112 ;
	7'h05 :
		RG_rl_100_t1 = TR_112 ;
	7'h06 :
		RG_rl_100_t1 = TR_112 ;
	7'h07 :
		RG_rl_100_t1 = TR_112 ;
	7'h08 :
		RG_rl_100_t1 = TR_112 ;
	7'h09 :
		RG_rl_100_t1 = TR_112 ;
	7'h0a :
		RG_rl_100_t1 = TR_112 ;
	7'h0b :
		RG_rl_100_t1 = TR_112 ;
	7'h0c :
		RG_rl_100_t1 = TR_112 ;
	7'h0d :
		RG_rl_100_t1 = TR_112 ;
	7'h0e :
		RG_rl_100_t1 = TR_112 ;
	7'h0f :
		RG_rl_100_t1 = TR_112 ;
	7'h10 :
		RG_rl_100_t1 = TR_112 ;
	7'h11 :
		RG_rl_100_t1 = TR_112 ;
	7'h12 :
		RG_rl_100_t1 = TR_112 ;
	7'h13 :
		RG_rl_100_t1 = TR_112 ;
	7'h14 :
		RG_rl_100_t1 = TR_112 ;
	7'h15 :
		RG_rl_100_t1 = TR_112 ;
	7'h16 :
		RG_rl_100_t1 = TR_112 ;
	7'h17 :
		RG_rl_100_t1 = TR_112 ;
	7'h18 :
		RG_rl_100_t1 = TR_112 ;
	7'h19 :
		RG_rl_100_t1 = TR_112 ;
	7'h1a :
		RG_rl_100_t1 = TR_112 ;
	7'h1b :
		RG_rl_100_t1 = TR_112 ;
	7'h1c :
		RG_rl_100_t1 = TR_112 ;
	7'h1d :
		RG_rl_100_t1 = TR_112 ;
	7'h1e :
		RG_rl_100_t1 = TR_112 ;
	7'h1f :
		RG_rl_100_t1 = TR_112 ;
	7'h20 :
		RG_rl_100_t1 = TR_112 ;
	7'h21 :
		RG_rl_100_t1 = TR_112 ;
	7'h22 :
		RG_rl_100_t1 = TR_112 ;
	7'h23 :
		RG_rl_100_t1 = TR_112 ;
	7'h24 :
		RG_rl_100_t1 = TR_112 ;
	7'h25 :
		RG_rl_100_t1 = TR_112 ;
	7'h26 :
		RG_rl_100_t1 = TR_112 ;
	7'h27 :
		RG_rl_100_t1 = TR_112 ;
	7'h28 :
		RG_rl_100_t1 = TR_112 ;
	7'h29 :
		RG_rl_100_t1 = TR_112 ;
	7'h2a :
		RG_rl_100_t1 = TR_112 ;
	7'h2b :
		RG_rl_100_t1 = TR_112 ;
	7'h2c :
		RG_rl_100_t1 = TR_112 ;
	7'h2d :
		RG_rl_100_t1 = TR_112 ;
	7'h2e :
		RG_rl_100_t1 = TR_112 ;
	7'h2f :
		RG_rl_100_t1 = TR_112 ;
	7'h30 :
		RG_rl_100_t1 = TR_112 ;
	7'h31 :
		RG_rl_100_t1 = TR_112 ;
	7'h32 :
		RG_rl_100_t1 = TR_112 ;
	7'h33 :
		RG_rl_100_t1 = TR_112 ;
	7'h34 :
		RG_rl_100_t1 = TR_112 ;
	7'h35 :
		RG_rl_100_t1 = TR_112 ;
	7'h36 :
		RG_rl_100_t1 = TR_112 ;
	7'h37 :
		RG_rl_100_t1 = TR_112 ;
	7'h38 :
		RG_rl_100_t1 = TR_112 ;
	7'h39 :
		RG_rl_100_t1 = TR_112 ;
	7'h3a :
		RG_rl_100_t1 = TR_112 ;
	7'h3b :
		RG_rl_100_t1 = TR_112 ;
	7'h3c :
		RG_rl_100_t1 = TR_112 ;
	7'h3d :
		RG_rl_100_t1 = TR_112 ;
	7'h3e :
		RG_rl_100_t1 = TR_112 ;
	7'h3f :
		RG_rl_100_t1 = TR_112 ;
	7'h40 :
		RG_rl_100_t1 = TR_112 ;
	7'h41 :
		RG_rl_100_t1 = TR_112 ;
	7'h42 :
		RG_rl_100_t1 = TR_112 ;
	7'h43 :
		RG_rl_100_t1 = TR_112 ;
	7'h44 :
		RG_rl_100_t1 = TR_112 ;
	7'h45 :
		RG_rl_100_t1 = TR_112 ;
	7'h46 :
		RG_rl_100_t1 = TR_112 ;
	7'h47 :
		RG_rl_100_t1 = TR_112 ;
	7'h48 :
		RG_rl_100_t1 = TR_112 ;
	7'h49 :
		RG_rl_100_t1 = TR_112 ;
	7'h4a :
		RG_rl_100_t1 = TR_112 ;
	7'h4b :
		RG_rl_100_t1 = TR_112 ;
	7'h4c :
		RG_rl_100_t1 = TR_112 ;
	7'h4d :
		RG_rl_100_t1 = TR_112 ;
	7'h4e :
		RG_rl_100_t1 = TR_112 ;
	7'h4f :
		RG_rl_100_t1 = TR_112 ;
	7'h50 :
		RG_rl_100_t1 = TR_112 ;
	7'h51 :
		RG_rl_100_t1 = TR_112 ;
	7'h52 :
		RG_rl_100_t1 = TR_112 ;
	7'h53 :
		RG_rl_100_t1 = TR_112 ;
	7'h54 :
		RG_rl_100_t1 = TR_112 ;
	7'h55 :
		RG_rl_100_t1 = TR_112 ;
	7'h56 :
		RG_rl_100_t1 = TR_112 ;
	7'h57 :
		RG_rl_100_t1 = TR_112 ;
	7'h58 :
		RG_rl_100_t1 = TR_112 ;
	7'h59 :
		RG_rl_100_t1 = TR_112 ;
	7'h5a :
		RG_rl_100_t1 = TR_112 ;
	7'h5b :
		RG_rl_100_t1 = TR_112 ;
	7'h5c :
		RG_rl_100_t1 = TR_112 ;
	7'h5d :
		RG_rl_100_t1 = TR_112 ;
	7'h5e :
		RG_rl_100_t1 = TR_112 ;
	7'h5f :
		RG_rl_100_t1 = TR_112 ;
	7'h60 :
		RG_rl_100_t1 = TR_112 ;
	7'h61 :
		RG_rl_100_t1 = TR_112 ;
	7'h62 :
		RG_rl_100_t1 = TR_112 ;
	7'h63 :
		RG_rl_100_t1 = TR_112 ;
	7'h64 :
		RG_rl_100_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h65 :
		RG_rl_100_t1 = TR_112 ;
	7'h66 :
		RG_rl_100_t1 = TR_112 ;
	7'h67 :
		RG_rl_100_t1 = TR_112 ;
	7'h68 :
		RG_rl_100_t1 = TR_112 ;
	7'h69 :
		RG_rl_100_t1 = TR_112 ;
	7'h6a :
		RG_rl_100_t1 = TR_112 ;
	7'h6b :
		RG_rl_100_t1 = TR_112 ;
	7'h6c :
		RG_rl_100_t1 = TR_112 ;
	7'h6d :
		RG_rl_100_t1 = TR_112 ;
	7'h6e :
		RG_rl_100_t1 = TR_112 ;
	7'h6f :
		RG_rl_100_t1 = TR_112 ;
	7'h70 :
		RG_rl_100_t1 = TR_112 ;
	7'h71 :
		RG_rl_100_t1 = TR_112 ;
	7'h72 :
		RG_rl_100_t1 = TR_112 ;
	7'h73 :
		RG_rl_100_t1 = TR_112 ;
	7'h74 :
		RG_rl_100_t1 = TR_112 ;
	7'h75 :
		RG_rl_100_t1 = TR_112 ;
	7'h76 :
		RG_rl_100_t1 = TR_112 ;
	7'h77 :
		RG_rl_100_t1 = TR_112 ;
	7'h78 :
		RG_rl_100_t1 = TR_112 ;
	7'h79 :
		RG_rl_100_t1 = TR_112 ;
	7'h7a :
		RG_rl_100_t1 = TR_112 ;
	7'h7b :
		RG_rl_100_t1 = TR_112 ;
	7'h7c :
		RG_rl_100_t1 = TR_112 ;
	7'h7d :
		RG_rl_100_t1 = TR_112 ;
	7'h7e :
		RG_rl_100_t1 = TR_112 ;
	7'h7f :
		RG_rl_100_t1 = TR_112 ;
	default :
		RG_rl_100_t1 = 9'hx ;
	endcase
always @ ( RG_rl_100_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_41 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_100_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h64 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_100_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_41 )
		| ( { 9{ U_569 } } & RG_rl_100_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_100_en = ( U_570 | RG_rl_100_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_100_en )
		RG_rl_100 <= RG_rl_100_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_113 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_101_t1 = TR_113 ;
	7'h01 :
		RG_rl_101_t1 = TR_113 ;
	7'h02 :
		RG_rl_101_t1 = TR_113 ;
	7'h03 :
		RG_rl_101_t1 = TR_113 ;
	7'h04 :
		RG_rl_101_t1 = TR_113 ;
	7'h05 :
		RG_rl_101_t1 = TR_113 ;
	7'h06 :
		RG_rl_101_t1 = TR_113 ;
	7'h07 :
		RG_rl_101_t1 = TR_113 ;
	7'h08 :
		RG_rl_101_t1 = TR_113 ;
	7'h09 :
		RG_rl_101_t1 = TR_113 ;
	7'h0a :
		RG_rl_101_t1 = TR_113 ;
	7'h0b :
		RG_rl_101_t1 = TR_113 ;
	7'h0c :
		RG_rl_101_t1 = TR_113 ;
	7'h0d :
		RG_rl_101_t1 = TR_113 ;
	7'h0e :
		RG_rl_101_t1 = TR_113 ;
	7'h0f :
		RG_rl_101_t1 = TR_113 ;
	7'h10 :
		RG_rl_101_t1 = TR_113 ;
	7'h11 :
		RG_rl_101_t1 = TR_113 ;
	7'h12 :
		RG_rl_101_t1 = TR_113 ;
	7'h13 :
		RG_rl_101_t1 = TR_113 ;
	7'h14 :
		RG_rl_101_t1 = TR_113 ;
	7'h15 :
		RG_rl_101_t1 = TR_113 ;
	7'h16 :
		RG_rl_101_t1 = TR_113 ;
	7'h17 :
		RG_rl_101_t1 = TR_113 ;
	7'h18 :
		RG_rl_101_t1 = TR_113 ;
	7'h19 :
		RG_rl_101_t1 = TR_113 ;
	7'h1a :
		RG_rl_101_t1 = TR_113 ;
	7'h1b :
		RG_rl_101_t1 = TR_113 ;
	7'h1c :
		RG_rl_101_t1 = TR_113 ;
	7'h1d :
		RG_rl_101_t1 = TR_113 ;
	7'h1e :
		RG_rl_101_t1 = TR_113 ;
	7'h1f :
		RG_rl_101_t1 = TR_113 ;
	7'h20 :
		RG_rl_101_t1 = TR_113 ;
	7'h21 :
		RG_rl_101_t1 = TR_113 ;
	7'h22 :
		RG_rl_101_t1 = TR_113 ;
	7'h23 :
		RG_rl_101_t1 = TR_113 ;
	7'h24 :
		RG_rl_101_t1 = TR_113 ;
	7'h25 :
		RG_rl_101_t1 = TR_113 ;
	7'h26 :
		RG_rl_101_t1 = TR_113 ;
	7'h27 :
		RG_rl_101_t1 = TR_113 ;
	7'h28 :
		RG_rl_101_t1 = TR_113 ;
	7'h29 :
		RG_rl_101_t1 = TR_113 ;
	7'h2a :
		RG_rl_101_t1 = TR_113 ;
	7'h2b :
		RG_rl_101_t1 = TR_113 ;
	7'h2c :
		RG_rl_101_t1 = TR_113 ;
	7'h2d :
		RG_rl_101_t1 = TR_113 ;
	7'h2e :
		RG_rl_101_t1 = TR_113 ;
	7'h2f :
		RG_rl_101_t1 = TR_113 ;
	7'h30 :
		RG_rl_101_t1 = TR_113 ;
	7'h31 :
		RG_rl_101_t1 = TR_113 ;
	7'h32 :
		RG_rl_101_t1 = TR_113 ;
	7'h33 :
		RG_rl_101_t1 = TR_113 ;
	7'h34 :
		RG_rl_101_t1 = TR_113 ;
	7'h35 :
		RG_rl_101_t1 = TR_113 ;
	7'h36 :
		RG_rl_101_t1 = TR_113 ;
	7'h37 :
		RG_rl_101_t1 = TR_113 ;
	7'h38 :
		RG_rl_101_t1 = TR_113 ;
	7'h39 :
		RG_rl_101_t1 = TR_113 ;
	7'h3a :
		RG_rl_101_t1 = TR_113 ;
	7'h3b :
		RG_rl_101_t1 = TR_113 ;
	7'h3c :
		RG_rl_101_t1 = TR_113 ;
	7'h3d :
		RG_rl_101_t1 = TR_113 ;
	7'h3e :
		RG_rl_101_t1 = TR_113 ;
	7'h3f :
		RG_rl_101_t1 = TR_113 ;
	7'h40 :
		RG_rl_101_t1 = TR_113 ;
	7'h41 :
		RG_rl_101_t1 = TR_113 ;
	7'h42 :
		RG_rl_101_t1 = TR_113 ;
	7'h43 :
		RG_rl_101_t1 = TR_113 ;
	7'h44 :
		RG_rl_101_t1 = TR_113 ;
	7'h45 :
		RG_rl_101_t1 = TR_113 ;
	7'h46 :
		RG_rl_101_t1 = TR_113 ;
	7'h47 :
		RG_rl_101_t1 = TR_113 ;
	7'h48 :
		RG_rl_101_t1 = TR_113 ;
	7'h49 :
		RG_rl_101_t1 = TR_113 ;
	7'h4a :
		RG_rl_101_t1 = TR_113 ;
	7'h4b :
		RG_rl_101_t1 = TR_113 ;
	7'h4c :
		RG_rl_101_t1 = TR_113 ;
	7'h4d :
		RG_rl_101_t1 = TR_113 ;
	7'h4e :
		RG_rl_101_t1 = TR_113 ;
	7'h4f :
		RG_rl_101_t1 = TR_113 ;
	7'h50 :
		RG_rl_101_t1 = TR_113 ;
	7'h51 :
		RG_rl_101_t1 = TR_113 ;
	7'h52 :
		RG_rl_101_t1 = TR_113 ;
	7'h53 :
		RG_rl_101_t1 = TR_113 ;
	7'h54 :
		RG_rl_101_t1 = TR_113 ;
	7'h55 :
		RG_rl_101_t1 = TR_113 ;
	7'h56 :
		RG_rl_101_t1 = TR_113 ;
	7'h57 :
		RG_rl_101_t1 = TR_113 ;
	7'h58 :
		RG_rl_101_t1 = TR_113 ;
	7'h59 :
		RG_rl_101_t1 = TR_113 ;
	7'h5a :
		RG_rl_101_t1 = TR_113 ;
	7'h5b :
		RG_rl_101_t1 = TR_113 ;
	7'h5c :
		RG_rl_101_t1 = TR_113 ;
	7'h5d :
		RG_rl_101_t1 = TR_113 ;
	7'h5e :
		RG_rl_101_t1 = TR_113 ;
	7'h5f :
		RG_rl_101_t1 = TR_113 ;
	7'h60 :
		RG_rl_101_t1 = TR_113 ;
	7'h61 :
		RG_rl_101_t1 = TR_113 ;
	7'h62 :
		RG_rl_101_t1 = TR_113 ;
	7'h63 :
		RG_rl_101_t1 = TR_113 ;
	7'h64 :
		RG_rl_101_t1 = TR_113 ;
	7'h65 :
		RG_rl_101_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h66 :
		RG_rl_101_t1 = TR_113 ;
	7'h67 :
		RG_rl_101_t1 = TR_113 ;
	7'h68 :
		RG_rl_101_t1 = TR_113 ;
	7'h69 :
		RG_rl_101_t1 = TR_113 ;
	7'h6a :
		RG_rl_101_t1 = TR_113 ;
	7'h6b :
		RG_rl_101_t1 = TR_113 ;
	7'h6c :
		RG_rl_101_t1 = TR_113 ;
	7'h6d :
		RG_rl_101_t1 = TR_113 ;
	7'h6e :
		RG_rl_101_t1 = TR_113 ;
	7'h6f :
		RG_rl_101_t1 = TR_113 ;
	7'h70 :
		RG_rl_101_t1 = TR_113 ;
	7'h71 :
		RG_rl_101_t1 = TR_113 ;
	7'h72 :
		RG_rl_101_t1 = TR_113 ;
	7'h73 :
		RG_rl_101_t1 = TR_113 ;
	7'h74 :
		RG_rl_101_t1 = TR_113 ;
	7'h75 :
		RG_rl_101_t1 = TR_113 ;
	7'h76 :
		RG_rl_101_t1 = TR_113 ;
	7'h77 :
		RG_rl_101_t1 = TR_113 ;
	7'h78 :
		RG_rl_101_t1 = TR_113 ;
	7'h79 :
		RG_rl_101_t1 = TR_113 ;
	7'h7a :
		RG_rl_101_t1 = TR_113 ;
	7'h7b :
		RG_rl_101_t1 = TR_113 ;
	7'h7c :
		RG_rl_101_t1 = TR_113 ;
	7'h7d :
		RG_rl_101_t1 = TR_113 ;
	7'h7e :
		RG_rl_101_t1 = TR_113 ;
	7'h7f :
		RG_rl_101_t1 = TR_113 ;
	default :
		RG_rl_101_t1 = 9'hx ;
	endcase
always @ ( RG_rl_101_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_42 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_101_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h65 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_101_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_42 )
		| ( { 9{ U_569 } } & RG_rl_101_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_101_en = ( U_570 | RG_rl_101_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_101_en )
		RG_rl_101 <= RG_rl_101_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_114 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_102_t1 = TR_114 ;
	7'h01 :
		RG_rl_102_t1 = TR_114 ;
	7'h02 :
		RG_rl_102_t1 = TR_114 ;
	7'h03 :
		RG_rl_102_t1 = TR_114 ;
	7'h04 :
		RG_rl_102_t1 = TR_114 ;
	7'h05 :
		RG_rl_102_t1 = TR_114 ;
	7'h06 :
		RG_rl_102_t1 = TR_114 ;
	7'h07 :
		RG_rl_102_t1 = TR_114 ;
	7'h08 :
		RG_rl_102_t1 = TR_114 ;
	7'h09 :
		RG_rl_102_t1 = TR_114 ;
	7'h0a :
		RG_rl_102_t1 = TR_114 ;
	7'h0b :
		RG_rl_102_t1 = TR_114 ;
	7'h0c :
		RG_rl_102_t1 = TR_114 ;
	7'h0d :
		RG_rl_102_t1 = TR_114 ;
	7'h0e :
		RG_rl_102_t1 = TR_114 ;
	7'h0f :
		RG_rl_102_t1 = TR_114 ;
	7'h10 :
		RG_rl_102_t1 = TR_114 ;
	7'h11 :
		RG_rl_102_t1 = TR_114 ;
	7'h12 :
		RG_rl_102_t1 = TR_114 ;
	7'h13 :
		RG_rl_102_t1 = TR_114 ;
	7'h14 :
		RG_rl_102_t1 = TR_114 ;
	7'h15 :
		RG_rl_102_t1 = TR_114 ;
	7'h16 :
		RG_rl_102_t1 = TR_114 ;
	7'h17 :
		RG_rl_102_t1 = TR_114 ;
	7'h18 :
		RG_rl_102_t1 = TR_114 ;
	7'h19 :
		RG_rl_102_t1 = TR_114 ;
	7'h1a :
		RG_rl_102_t1 = TR_114 ;
	7'h1b :
		RG_rl_102_t1 = TR_114 ;
	7'h1c :
		RG_rl_102_t1 = TR_114 ;
	7'h1d :
		RG_rl_102_t1 = TR_114 ;
	7'h1e :
		RG_rl_102_t1 = TR_114 ;
	7'h1f :
		RG_rl_102_t1 = TR_114 ;
	7'h20 :
		RG_rl_102_t1 = TR_114 ;
	7'h21 :
		RG_rl_102_t1 = TR_114 ;
	7'h22 :
		RG_rl_102_t1 = TR_114 ;
	7'h23 :
		RG_rl_102_t1 = TR_114 ;
	7'h24 :
		RG_rl_102_t1 = TR_114 ;
	7'h25 :
		RG_rl_102_t1 = TR_114 ;
	7'h26 :
		RG_rl_102_t1 = TR_114 ;
	7'h27 :
		RG_rl_102_t1 = TR_114 ;
	7'h28 :
		RG_rl_102_t1 = TR_114 ;
	7'h29 :
		RG_rl_102_t1 = TR_114 ;
	7'h2a :
		RG_rl_102_t1 = TR_114 ;
	7'h2b :
		RG_rl_102_t1 = TR_114 ;
	7'h2c :
		RG_rl_102_t1 = TR_114 ;
	7'h2d :
		RG_rl_102_t1 = TR_114 ;
	7'h2e :
		RG_rl_102_t1 = TR_114 ;
	7'h2f :
		RG_rl_102_t1 = TR_114 ;
	7'h30 :
		RG_rl_102_t1 = TR_114 ;
	7'h31 :
		RG_rl_102_t1 = TR_114 ;
	7'h32 :
		RG_rl_102_t1 = TR_114 ;
	7'h33 :
		RG_rl_102_t1 = TR_114 ;
	7'h34 :
		RG_rl_102_t1 = TR_114 ;
	7'h35 :
		RG_rl_102_t1 = TR_114 ;
	7'h36 :
		RG_rl_102_t1 = TR_114 ;
	7'h37 :
		RG_rl_102_t1 = TR_114 ;
	7'h38 :
		RG_rl_102_t1 = TR_114 ;
	7'h39 :
		RG_rl_102_t1 = TR_114 ;
	7'h3a :
		RG_rl_102_t1 = TR_114 ;
	7'h3b :
		RG_rl_102_t1 = TR_114 ;
	7'h3c :
		RG_rl_102_t1 = TR_114 ;
	7'h3d :
		RG_rl_102_t1 = TR_114 ;
	7'h3e :
		RG_rl_102_t1 = TR_114 ;
	7'h3f :
		RG_rl_102_t1 = TR_114 ;
	7'h40 :
		RG_rl_102_t1 = TR_114 ;
	7'h41 :
		RG_rl_102_t1 = TR_114 ;
	7'h42 :
		RG_rl_102_t1 = TR_114 ;
	7'h43 :
		RG_rl_102_t1 = TR_114 ;
	7'h44 :
		RG_rl_102_t1 = TR_114 ;
	7'h45 :
		RG_rl_102_t1 = TR_114 ;
	7'h46 :
		RG_rl_102_t1 = TR_114 ;
	7'h47 :
		RG_rl_102_t1 = TR_114 ;
	7'h48 :
		RG_rl_102_t1 = TR_114 ;
	7'h49 :
		RG_rl_102_t1 = TR_114 ;
	7'h4a :
		RG_rl_102_t1 = TR_114 ;
	7'h4b :
		RG_rl_102_t1 = TR_114 ;
	7'h4c :
		RG_rl_102_t1 = TR_114 ;
	7'h4d :
		RG_rl_102_t1 = TR_114 ;
	7'h4e :
		RG_rl_102_t1 = TR_114 ;
	7'h4f :
		RG_rl_102_t1 = TR_114 ;
	7'h50 :
		RG_rl_102_t1 = TR_114 ;
	7'h51 :
		RG_rl_102_t1 = TR_114 ;
	7'h52 :
		RG_rl_102_t1 = TR_114 ;
	7'h53 :
		RG_rl_102_t1 = TR_114 ;
	7'h54 :
		RG_rl_102_t1 = TR_114 ;
	7'h55 :
		RG_rl_102_t1 = TR_114 ;
	7'h56 :
		RG_rl_102_t1 = TR_114 ;
	7'h57 :
		RG_rl_102_t1 = TR_114 ;
	7'h58 :
		RG_rl_102_t1 = TR_114 ;
	7'h59 :
		RG_rl_102_t1 = TR_114 ;
	7'h5a :
		RG_rl_102_t1 = TR_114 ;
	7'h5b :
		RG_rl_102_t1 = TR_114 ;
	7'h5c :
		RG_rl_102_t1 = TR_114 ;
	7'h5d :
		RG_rl_102_t1 = TR_114 ;
	7'h5e :
		RG_rl_102_t1 = TR_114 ;
	7'h5f :
		RG_rl_102_t1 = TR_114 ;
	7'h60 :
		RG_rl_102_t1 = TR_114 ;
	7'h61 :
		RG_rl_102_t1 = TR_114 ;
	7'h62 :
		RG_rl_102_t1 = TR_114 ;
	7'h63 :
		RG_rl_102_t1 = TR_114 ;
	7'h64 :
		RG_rl_102_t1 = TR_114 ;
	7'h65 :
		RG_rl_102_t1 = TR_114 ;
	7'h66 :
		RG_rl_102_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h67 :
		RG_rl_102_t1 = TR_114 ;
	7'h68 :
		RG_rl_102_t1 = TR_114 ;
	7'h69 :
		RG_rl_102_t1 = TR_114 ;
	7'h6a :
		RG_rl_102_t1 = TR_114 ;
	7'h6b :
		RG_rl_102_t1 = TR_114 ;
	7'h6c :
		RG_rl_102_t1 = TR_114 ;
	7'h6d :
		RG_rl_102_t1 = TR_114 ;
	7'h6e :
		RG_rl_102_t1 = TR_114 ;
	7'h6f :
		RG_rl_102_t1 = TR_114 ;
	7'h70 :
		RG_rl_102_t1 = TR_114 ;
	7'h71 :
		RG_rl_102_t1 = TR_114 ;
	7'h72 :
		RG_rl_102_t1 = TR_114 ;
	7'h73 :
		RG_rl_102_t1 = TR_114 ;
	7'h74 :
		RG_rl_102_t1 = TR_114 ;
	7'h75 :
		RG_rl_102_t1 = TR_114 ;
	7'h76 :
		RG_rl_102_t1 = TR_114 ;
	7'h77 :
		RG_rl_102_t1 = TR_114 ;
	7'h78 :
		RG_rl_102_t1 = TR_114 ;
	7'h79 :
		RG_rl_102_t1 = TR_114 ;
	7'h7a :
		RG_rl_102_t1 = TR_114 ;
	7'h7b :
		RG_rl_102_t1 = TR_114 ;
	7'h7c :
		RG_rl_102_t1 = TR_114 ;
	7'h7d :
		RG_rl_102_t1 = TR_114 ;
	7'h7e :
		RG_rl_102_t1 = TR_114 ;
	7'h7f :
		RG_rl_102_t1 = TR_114 ;
	default :
		RG_rl_102_t1 = 9'hx ;
	endcase
always @ ( RG_rl_102_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_43 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_102_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h66 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_102_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_43 )
		| ( { 9{ U_569 } } & RG_rl_102_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_102_en = ( U_570 | RG_rl_102_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_102_en )
		RG_rl_102 <= RG_rl_102_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_115 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_103_t1 = TR_115 ;
	7'h01 :
		RG_rl_103_t1 = TR_115 ;
	7'h02 :
		RG_rl_103_t1 = TR_115 ;
	7'h03 :
		RG_rl_103_t1 = TR_115 ;
	7'h04 :
		RG_rl_103_t1 = TR_115 ;
	7'h05 :
		RG_rl_103_t1 = TR_115 ;
	7'h06 :
		RG_rl_103_t1 = TR_115 ;
	7'h07 :
		RG_rl_103_t1 = TR_115 ;
	7'h08 :
		RG_rl_103_t1 = TR_115 ;
	7'h09 :
		RG_rl_103_t1 = TR_115 ;
	7'h0a :
		RG_rl_103_t1 = TR_115 ;
	7'h0b :
		RG_rl_103_t1 = TR_115 ;
	7'h0c :
		RG_rl_103_t1 = TR_115 ;
	7'h0d :
		RG_rl_103_t1 = TR_115 ;
	7'h0e :
		RG_rl_103_t1 = TR_115 ;
	7'h0f :
		RG_rl_103_t1 = TR_115 ;
	7'h10 :
		RG_rl_103_t1 = TR_115 ;
	7'h11 :
		RG_rl_103_t1 = TR_115 ;
	7'h12 :
		RG_rl_103_t1 = TR_115 ;
	7'h13 :
		RG_rl_103_t1 = TR_115 ;
	7'h14 :
		RG_rl_103_t1 = TR_115 ;
	7'h15 :
		RG_rl_103_t1 = TR_115 ;
	7'h16 :
		RG_rl_103_t1 = TR_115 ;
	7'h17 :
		RG_rl_103_t1 = TR_115 ;
	7'h18 :
		RG_rl_103_t1 = TR_115 ;
	7'h19 :
		RG_rl_103_t1 = TR_115 ;
	7'h1a :
		RG_rl_103_t1 = TR_115 ;
	7'h1b :
		RG_rl_103_t1 = TR_115 ;
	7'h1c :
		RG_rl_103_t1 = TR_115 ;
	7'h1d :
		RG_rl_103_t1 = TR_115 ;
	7'h1e :
		RG_rl_103_t1 = TR_115 ;
	7'h1f :
		RG_rl_103_t1 = TR_115 ;
	7'h20 :
		RG_rl_103_t1 = TR_115 ;
	7'h21 :
		RG_rl_103_t1 = TR_115 ;
	7'h22 :
		RG_rl_103_t1 = TR_115 ;
	7'h23 :
		RG_rl_103_t1 = TR_115 ;
	7'h24 :
		RG_rl_103_t1 = TR_115 ;
	7'h25 :
		RG_rl_103_t1 = TR_115 ;
	7'h26 :
		RG_rl_103_t1 = TR_115 ;
	7'h27 :
		RG_rl_103_t1 = TR_115 ;
	7'h28 :
		RG_rl_103_t1 = TR_115 ;
	7'h29 :
		RG_rl_103_t1 = TR_115 ;
	7'h2a :
		RG_rl_103_t1 = TR_115 ;
	7'h2b :
		RG_rl_103_t1 = TR_115 ;
	7'h2c :
		RG_rl_103_t1 = TR_115 ;
	7'h2d :
		RG_rl_103_t1 = TR_115 ;
	7'h2e :
		RG_rl_103_t1 = TR_115 ;
	7'h2f :
		RG_rl_103_t1 = TR_115 ;
	7'h30 :
		RG_rl_103_t1 = TR_115 ;
	7'h31 :
		RG_rl_103_t1 = TR_115 ;
	7'h32 :
		RG_rl_103_t1 = TR_115 ;
	7'h33 :
		RG_rl_103_t1 = TR_115 ;
	7'h34 :
		RG_rl_103_t1 = TR_115 ;
	7'h35 :
		RG_rl_103_t1 = TR_115 ;
	7'h36 :
		RG_rl_103_t1 = TR_115 ;
	7'h37 :
		RG_rl_103_t1 = TR_115 ;
	7'h38 :
		RG_rl_103_t1 = TR_115 ;
	7'h39 :
		RG_rl_103_t1 = TR_115 ;
	7'h3a :
		RG_rl_103_t1 = TR_115 ;
	7'h3b :
		RG_rl_103_t1 = TR_115 ;
	7'h3c :
		RG_rl_103_t1 = TR_115 ;
	7'h3d :
		RG_rl_103_t1 = TR_115 ;
	7'h3e :
		RG_rl_103_t1 = TR_115 ;
	7'h3f :
		RG_rl_103_t1 = TR_115 ;
	7'h40 :
		RG_rl_103_t1 = TR_115 ;
	7'h41 :
		RG_rl_103_t1 = TR_115 ;
	7'h42 :
		RG_rl_103_t1 = TR_115 ;
	7'h43 :
		RG_rl_103_t1 = TR_115 ;
	7'h44 :
		RG_rl_103_t1 = TR_115 ;
	7'h45 :
		RG_rl_103_t1 = TR_115 ;
	7'h46 :
		RG_rl_103_t1 = TR_115 ;
	7'h47 :
		RG_rl_103_t1 = TR_115 ;
	7'h48 :
		RG_rl_103_t1 = TR_115 ;
	7'h49 :
		RG_rl_103_t1 = TR_115 ;
	7'h4a :
		RG_rl_103_t1 = TR_115 ;
	7'h4b :
		RG_rl_103_t1 = TR_115 ;
	7'h4c :
		RG_rl_103_t1 = TR_115 ;
	7'h4d :
		RG_rl_103_t1 = TR_115 ;
	7'h4e :
		RG_rl_103_t1 = TR_115 ;
	7'h4f :
		RG_rl_103_t1 = TR_115 ;
	7'h50 :
		RG_rl_103_t1 = TR_115 ;
	7'h51 :
		RG_rl_103_t1 = TR_115 ;
	7'h52 :
		RG_rl_103_t1 = TR_115 ;
	7'h53 :
		RG_rl_103_t1 = TR_115 ;
	7'h54 :
		RG_rl_103_t1 = TR_115 ;
	7'h55 :
		RG_rl_103_t1 = TR_115 ;
	7'h56 :
		RG_rl_103_t1 = TR_115 ;
	7'h57 :
		RG_rl_103_t1 = TR_115 ;
	7'h58 :
		RG_rl_103_t1 = TR_115 ;
	7'h59 :
		RG_rl_103_t1 = TR_115 ;
	7'h5a :
		RG_rl_103_t1 = TR_115 ;
	7'h5b :
		RG_rl_103_t1 = TR_115 ;
	7'h5c :
		RG_rl_103_t1 = TR_115 ;
	7'h5d :
		RG_rl_103_t1 = TR_115 ;
	7'h5e :
		RG_rl_103_t1 = TR_115 ;
	7'h5f :
		RG_rl_103_t1 = TR_115 ;
	7'h60 :
		RG_rl_103_t1 = TR_115 ;
	7'h61 :
		RG_rl_103_t1 = TR_115 ;
	7'h62 :
		RG_rl_103_t1 = TR_115 ;
	7'h63 :
		RG_rl_103_t1 = TR_115 ;
	7'h64 :
		RG_rl_103_t1 = TR_115 ;
	7'h65 :
		RG_rl_103_t1 = TR_115 ;
	7'h66 :
		RG_rl_103_t1 = TR_115 ;
	7'h67 :
		RG_rl_103_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h68 :
		RG_rl_103_t1 = TR_115 ;
	7'h69 :
		RG_rl_103_t1 = TR_115 ;
	7'h6a :
		RG_rl_103_t1 = TR_115 ;
	7'h6b :
		RG_rl_103_t1 = TR_115 ;
	7'h6c :
		RG_rl_103_t1 = TR_115 ;
	7'h6d :
		RG_rl_103_t1 = TR_115 ;
	7'h6e :
		RG_rl_103_t1 = TR_115 ;
	7'h6f :
		RG_rl_103_t1 = TR_115 ;
	7'h70 :
		RG_rl_103_t1 = TR_115 ;
	7'h71 :
		RG_rl_103_t1 = TR_115 ;
	7'h72 :
		RG_rl_103_t1 = TR_115 ;
	7'h73 :
		RG_rl_103_t1 = TR_115 ;
	7'h74 :
		RG_rl_103_t1 = TR_115 ;
	7'h75 :
		RG_rl_103_t1 = TR_115 ;
	7'h76 :
		RG_rl_103_t1 = TR_115 ;
	7'h77 :
		RG_rl_103_t1 = TR_115 ;
	7'h78 :
		RG_rl_103_t1 = TR_115 ;
	7'h79 :
		RG_rl_103_t1 = TR_115 ;
	7'h7a :
		RG_rl_103_t1 = TR_115 ;
	7'h7b :
		RG_rl_103_t1 = TR_115 ;
	7'h7c :
		RG_rl_103_t1 = TR_115 ;
	7'h7d :
		RG_rl_103_t1 = TR_115 ;
	7'h7e :
		RG_rl_103_t1 = TR_115 ;
	7'h7f :
		RG_rl_103_t1 = TR_115 ;
	default :
		RG_rl_103_t1 = 9'hx ;
	endcase
always @ ( RG_rl_103_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_44 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_103_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h67 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_103_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_44 )
		| ( { 9{ U_569 } } & RG_rl_103_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_103_en = ( U_570 | RG_rl_103_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_103_en )
		RG_rl_103 <= RG_rl_103_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_116 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_104_t1 = TR_116 ;
	7'h01 :
		RG_rl_104_t1 = TR_116 ;
	7'h02 :
		RG_rl_104_t1 = TR_116 ;
	7'h03 :
		RG_rl_104_t1 = TR_116 ;
	7'h04 :
		RG_rl_104_t1 = TR_116 ;
	7'h05 :
		RG_rl_104_t1 = TR_116 ;
	7'h06 :
		RG_rl_104_t1 = TR_116 ;
	7'h07 :
		RG_rl_104_t1 = TR_116 ;
	7'h08 :
		RG_rl_104_t1 = TR_116 ;
	7'h09 :
		RG_rl_104_t1 = TR_116 ;
	7'h0a :
		RG_rl_104_t1 = TR_116 ;
	7'h0b :
		RG_rl_104_t1 = TR_116 ;
	7'h0c :
		RG_rl_104_t1 = TR_116 ;
	7'h0d :
		RG_rl_104_t1 = TR_116 ;
	7'h0e :
		RG_rl_104_t1 = TR_116 ;
	7'h0f :
		RG_rl_104_t1 = TR_116 ;
	7'h10 :
		RG_rl_104_t1 = TR_116 ;
	7'h11 :
		RG_rl_104_t1 = TR_116 ;
	7'h12 :
		RG_rl_104_t1 = TR_116 ;
	7'h13 :
		RG_rl_104_t1 = TR_116 ;
	7'h14 :
		RG_rl_104_t1 = TR_116 ;
	7'h15 :
		RG_rl_104_t1 = TR_116 ;
	7'h16 :
		RG_rl_104_t1 = TR_116 ;
	7'h17 :
		RG_rl_104_t1 = TR_116 ;
	7'h18 :
		RG_rl_104_t1 = TR_116 ;
	7'h19 :
		RG_rl_104_t1 = TR_116 ;
	7'h1a :
		RG_rl_104_t1 = TR_116 ;
	7'h1b :
		RG_rl_104_t1 = TR_116 ;
	7'h1c :
		RG_rl_104_t1 = TR_116 ;
	7'h1d :
		RG_rl_104_t1 = TR_116 ;
	7'h1e :
		RG_rl_104_t1 = TR_116 ;
	7'h1f :
		RG_rl_104_t1 = TR_116 ;
	7'h20 :
		RG_rl_104_t1 = TR_116 ;
	7'h21 :
		RG_rl_104_t1 = TR_116 ;
	7'h22 :
		RG_rl_104_t1 = TR_116 ;
	7'h23 :
		RG_rl_104_t1 = TR_116 ;
	7'h24 :
		RG_rl_104_t1 = TR_116 ;
	7'h25 :
		RG_rl_104_t1 = TR_116 ;
	7'h26 :
		RG_rl_104_t1 = TR_116 ;
	7'h27 :
		RG_rl_104_t1 = TR_116 ;
	7'h28 :
		RG_rl_104_t1 = TR_116 ;
	7'h29 :
		RG_rl_104_t1 = TR_116 ;
	7'h2a :
		RG_rl_104_t1 = TR_116 ;
	7'h2b :
		RG_rl_104_t1 = TR_116 ;
	7'h2c :
		RG_rl_104_t1 = TR_116 ;
	7'h2d :
		RG_rl_104_t1 = TR_116 ;
	7'h2e :
		RG_rl_104_t1 = TR_116 ;
	7'h2f :
		RG_rl_104_t1 = TR_116 ;
	7'h30 :
		RG_rl_104_t1 = TR_116 ;
	7'h31 :
		RG_rl_104_t1 = TR_116 ;
	7'h32 :
		RG_rl_104_t1 = TR_116 ;
	7'h33 :
		RG_rl_104_t1 = TR_116 ;
	7'h34 :
		RG_rl_104_t1 = TR_116 ;
	7'h35 :
		RG_rl_104_t1 = TR_116 ;
	7'h36 :
		RG_rl_104_t1 = TR_116 ;
	7'h37 :
		RG_rl_104_t1 = TR_116 ;
	7'h38 :
		RG_rl_104_t1 = TR_116 ;
	7'h39 :
		RG_rl_104_t1 = TR_116 ;
	7'h3a :
		RG_rl_104_t1 = TR_116 ;
	7'h3b :
		RG_rl_104_t1 = TR_116 ;
	7'h3c :
		RG_rl_104_t1 = TR_116 ;
	7'h3d :
		RG_rl_104_t1 = TR_116 ;
	7'h3e :
		RG_rl_104_t1 = TR_116 ;
	7'h3f :
		RG_rl_104_t1 = TR_116 ;
	7'h40 :
		RG_rl_104_t1 = TR_116 ;
	7'h41 :
		RG_rl_104_t1 = TR_116 ;
	7'h42 :
		RG_rl_104_t1 = TR_116 ;
	7'h43 :
		RG_rl_104_t1 = TR_116 ;
	7'h44 :
		RG_rl_104_t1 = TR_116 ;
	7'h45 :
		RG_rl_104_t1 = TR_116 ;
	7'h46 :
		RG_rl_104_t1 = TR_116 ;
	7'h47 :
		RG_rl_104_t1 = TR_116 ;
	7'h48 :
		RG_rl_104_t1 = TR_116 ;
	7'h49 :
		RG_rl_104_t1 = TR_116 ;
	7'h4a :
		RG_rl_104_t1 = TR_116 ;
	7'h4b :
		RG_rl_104_t1 = TR_116 ;
	7'h4c :
		RG_rl_104_t1 = TR_116 ;
	7'h4d :
		RG_rl_104_t1 = TR_116 ;
	7'h4e :
		RG_rl_104_t1 = TR_116 ;
	7'h4f :
		RG_rl_104_t1 = TR_116 ;
	7'h50 :
		RG_rl_104_t1 = TR_116 ;
	7'h51 :
		RG_rl_104_t1 = TR_116 ;
	7'h52 :
		RG_rl_104_t1 = TR_116 ;
	7'h53 :
		RG_rl_104_t1 = TR_116 ;
	7'h54 :
		RG_rl_104_t1 = TR_116 ;
	7'h55 :
		RG_rl_104_t1 = TR_116 ;
	7'h56 :
		RG_rl_104_t1 = TR_116 ;
	7'h57 :
		RG_rl_104_t1 = TR_116 ;
	7'h58 :
		RG_rl_104_t1 = TR_116 ;
	7'h59 :
		RG_rl_104_t1 = TR_116 ;
	7'h5a :
		RG_rl_104_t1 = TR_116 ;
	7'h5b :
		RG_rl_104_t1 = TR_116 ;
	7'h5c :
		RG_rl_104_t1 = TR_116 ;
	7'h5d :
		RG_rl_104_t1 = TR_116 ;
	7'h5e :
		RG_rl_104_t1 = TR_116 ;
	7'h5f :
		RG_rl_104_t1 = TR_116 ;
	7'h60 :
		RG_rl_104_t1 = TR_116 ;
	7'h61 :
		RG_rl_104_t1 = TR_116 ;
	7'h62 :
		RG_rl_104_t1 = TR_116 ;
	7'h63 :
		RG_rl_104_t1 = TR_116 ;
	7'h64 :
		RG_rl_104_t1 = TR_116 ;
	7'h65 :
		RG_rl_104_t1 = TR_116 ;
	7'h66 :
		RG_rl_104_t1 = TR_116 ;
	7'h67 :
		RG_rl_104_t1 = TR_116 ;
	7'h68 :
		RG_rl_104_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h69 :
		RG_rl_104_t1 = TR_116 ;
	7'h6a :
		RG_rl_104_t1 = TR_116 ;
	7'h6b :
		RG_rl_104_t1 = TR_116 ;
	7'h6c :
		RG_rl_104_t1 = TR_116 ;
	7'h6d :
		RG_rl_104_t1 = TR_116 ;
	7'h6e :
		RG_rl_104_t1 = TR_116 ;
	7'h6f :
		RG_rl_104_t1 = TR_116 ;
	7'h70 :
		RG_rl_104_t1 = TR_116 ;
	7'h71 :
		RG_rl_104_t1 = TR_116 ;
	7'h72 :
		RG_rl_104_t1 = TR_116 ;
	7'h73 :
		RG_rl_104_t1 = TR_116 ;
	7'h74 :
		RG_rl_104_t1 = TR_116 ;
	7'h75 :
		RG_rl_104_t1 = TR_116 ;
	7'h76 :
		RG_rl_104_t1 = TR_116 ;
	7'h77 :
		RG_rl_104_t1 = TR_116 ;
	7'h78 :
		RG_rl_104_t1 = TR_116 ;
	7'h79 :
		RG_rl_104_t1 = TR_116 ;
	7'h7a :
		RG_rl_104_t1 = TR_116 ;
	7'h7b :
		RG_rl_104_t1 = TR_116 ;
	7'h7c :
		RG_rl_104_t1 = TR_116 ;
	7'h7d :
		RG_rl_104_t1 = TR_116 ;
	7'h7e :
		RG_rl_104_t1 = TR_116 ;
	7'h7f :
		RG_rl_104_t1 = TR_116 ;
	default :
		RG_rl_104_t1 = 9'hx ;
	endcase
always @ ( RG_rl_104_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_45 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_104_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h68 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_104_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_45 )
		| ( { 9{ U_569 } } & RG_rl_104_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_104_en = ( U_570 | RG_rl_104_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_104_en )
		RG_rl_104 <= RG_rl_104_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_117 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_105_t1 = TR_117 ;
	7'h01 :
		RG_rl_105_t1 = TR_117 ;
	7'h02 :
		RG_rl_105_t1 = TR_117 ;
	7'h03 :
		RG_rl_105_t1 = TR_117 ;
	7'h04 :
		RG_rl_105_t1 = TR_117 ;
	7'h05 :
		RG_rl_105_t1 = TR_117 ;
	7'h06 :
		RG_rl_105_t1 = TR_117 ;
	7'h07 :
		RG_rl_105_t1 = TR_117 ;
	7'h08 :
		RG_rl_105_t1 = TR_117 ;
	7'h09 :
		RG_rl_105_t1 = TR_117 ;
	7'h0a :
		RG_rl_105_t1 = TR_117 ;
	7'h0b :
		RG_rl_105_t1 = TR_117 ;
	7'h0c :
		RG_rl_105_t1 = TR_117 ;
	7'h0d :
		RG_rl_105_t1 = TR_117 ;
	7'h0e :
		RG_rl_105_t1 = TR_117 ;
	7'h0f :
		RG_rl_105_t1 = TR_117 ;
	7'h10 :
		RG_rl_105_t1 = TR_117 ;
	7'h11 :
		RG_rl_105_t1 = TR_117 ;
	7'h12 :
		RG_rl_105_t1 = TR_117 ;
	7'h13 :
		RG_rl_105_t1 = TR_117 ;
	7'h14 :
		RG_rl_105_t1 = TR_117 ;
	7'h15 :
		RG_rl_105_t1 = TR_117 ;
	7'h16 :
		RG_rl_105_t1 = TR_117 ;
	7'h17 :
		RG_rl_105_t1 = TR_117 ;
	7'h18 :
		RG_rl_105_t1 = TR_117 ;
	7'h19 :
		RG_rl_105_t1 = TR_117 ;
	7'h1a :
		RG_rl_105_t1 = TR_117 ;
	7'h1b :
		RG_rl_105_t1 = TR_117 ;
	7'h1c :
		RG_rl_105_t1 = TR_117 ;
	7'h1d :
		RG_rl_105_t1 = TR_117 ;
	7'h1e :
		RG_rl_105_t1 = TR_117 ;
	7'h1f :
		RG_rl_105_t1 = TR_117 ;
	7'h20 :
		RG_rl_105_t1 = TR_117 ;
	7'h21 :
		RG_rl_105_t1 = TR_117 ;
	7'h22 :
		RG_rl_105_t1 = TR_117 ;
	7'h23 :
		RG_rl_105_t1 = TR_117 ;
	7'h24 :
		RG_rl_105_t1 = TR_117 ;
	7'h25 :
		RG_rl_105_t1 = TR_117 ;
	7'h26 :
		RG_rl_105_t1 = TR_117 ;
	7'h27 :
		RG_rl_105_t1 = TR_117 ;
	7'h28 :
		RG_rl_105_t1 = TR_117 ;
	7'h29 :
		RG_rl_105_t1 = TR_117 ;
	7'h2a :
		RG_rl_105_t1 = TR_117 ;
	7'h2b :
		RG_rl_105_t1 = TR_117 ;
	7'h2c :
		RG_rl_105_t1 = TR_117 ;
	7'h2d :
		RG_rl_105_t1 = TR_117 ;
	7'h2e :
		RG_rl_105_t1 = TR_117 ;
	7'h2f :
		RG_rl_105_t1 = TR_117 ;
	7'h30 :
		RG_rl_105_t1 = TR_117 ;
	7'h31 :
		RG_rl_105_t1 = TR_117 ;
	7'h32 :
		RG_rl_105_t1 = TR_117 ;
	7'h33 :
		RG_rl_105_t1 = TR_117 ;
	7'h34 :
		RG_rl_105_t1 = TR_117 ;
	7'h35 :
		RG_rl_105_t1 = TR_117 ;
	7'h36 :
		RG_rl_105_t1 = TR_117 ;
	7'h37 :
		RG_rl_105_t1 = TR_117 ;
	7'h38 :
		RG_rl_105_t1 = TR_117 ;
	7'h39 :
		RG_rl_105_t1 = TR_117 ;
	7'h3a :
		RG_rl_105_t1 = TR_117 ;
	7'h3b :
		RG_rl_105_t1 = TR_117 ;
	7'h3c :
		RG_rl_105_t1 = TR_117 ;
	7'h3d :
		RG_rl_105_t1 = TR_117 ;
	7'h3e :
		RG_rl_105_t1 = TR_117 ;
	7'h3f :
		RG_rl_105_t1 = TR_117 ;
	7'h40 :
		RG_rl_105_t1 = TR_117 ;
	7'h41 :
		RG_rl_105_t1 = TR_117 ;
	7'h42 :
		RG_rl_105_t1 = TR_117 ;
	7'h43 :
		RG_rl_105_t1 = TR_117 ;
	7'h44 :
		RG_rl_105_t1 = TR_117 ;
	7'h45 :
		RG_rl_105_t1 = TR_117 ;
	7'h46 :
		RG_rl_105_t1 = TR_117 ;
	7'h47 :
		RG_rl_105_t1 = TR_117 ;
	7'h48 :
		RG_rl_105_t1 = TR_117 ;
	7'h49 :
		RG_rl_105_t1 = TR_117 ;
	7'h4a :
		RG_rl_105_t1 = TR_117 ;
	7'h4b :
		RG_rl_105_t1 = TR_117 ;
	7'h4c :
		RG_rl_105_t1 = TR_117 ;
	7'h4d :
		RG_rl_105_t1 = TR_117 ;
	7'h4e :
		RG_rl_105_t1 = TR_117 ;
	7'h4f :
		RG_rl_105_t1 = TR_117 ;
	7'h50 :
		RG_rl_105_t1 = TR_117 ;
	7'h51 :
		RG_rl_105_t1 = TR_117 ;
	7'h52 :
		RG_rl_105_t1 = TR_117 ;
	7'h53 :
		RG_rl_105_t1 = TR_117 ;
	7'h54 :
		RG_rl_105_t1 = TR_117 ;
	7'h55 :
		RG_rl_105_t1 = TR_117 ;
	7'h56 :
		RG_rl_105_t1 = TR_117 ;
	7'h57 :
		RG_rl_105_t1 = TR_117 ;
	7'h58 :
		RG_rl_105_t1 = TR_117 ;
	7'h59 :
		RG_rl_105_t1 = TR_117 ;
	7'h5a :
		RG_rl_105_t1 = TR_117 ;
	7'h5b :
		RG_rl_105_t1 = TR_117 ;
	7'h5c :
		RG_rl_105_t1 = TR_117 ;
	7'h5d :
		RG_rl_105_t1 = TR_117 ;
	7'h5e :
		RG_rl_105_t1 = TR_117 ;
	7'h5f :
		RG_rl_105_t1 = TR_117 ;
	7'h60 :
		RG_rl_105_t1 = TR_117 ;
	7'h61 :
		RG_rl_105_t1 = TR_117 ;
	7'h62 :
		RG_rl_105_t1 = TR_117 ;
	7'h63 :
		RG_rl_105_t1 = TR_117 ;
	7'h64 :
		RG_rl_105_t1 = TR_117 ;
	7'h65 :
		RG_rl_105_t1 = TR_117 ;
	7'h66 :
		RG_rl_105_t1 = TR_117 ;
	7'h67 :
		RG_rl_105_t1 = TR_117 ;
	7'h68 :
		RG_rl_105_t1 = TR_117 ;
	7'h69 :
		RG_rl_105_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6a :
		RG_rl_105_t1 = TR_117 ;
	7'h6b :
		RG_rl_105_t1 = TR_117 ;
	7'h6c :
		RG_rl_105_t1 = TR_117 ;
	7'h6d :
		RG_rl_105_t1 = TR_117 ;
	7'h6e :
		RG_rl_105_t1 = TR_117 ;
	7'h6f :
		RG_rl_105_t1 = TR_117 ;
	7'h70 :
		RG_rl_105_t1 = TR_117 ;
	7'h71 :
		RG_rl_105_t1 = TR_117 ;
	7'h72 :
		RG_rl_105_t1 = TR_117 ;
	7'h73 :
		RG_rl_105_t1 = TR_117 ;
	7'h74 :
		RG_rl_105_t1 = TR_117 ;
	7'h75 :
		RG_rl_105_t1 = TR_117 ;
	7'h76 :
		RG_rl_105_t1 = TR_117 ;
	7'h77 :
		RG_rl_105_t1 = TR_117 ;
	7'h78 :
		RG_rl_105_t1 = TR_117 ;
	7'h79 :
		RG_rl_105_t1 = TR_117 ;
	7'h7a :
		RG_rl_105_t1 = TR_117 ;
	7'h7b :
		RG_rl_105_t1 = TR_117 ;
	7'h7c :
		RG_rl_105_t1 = TR_117 ;
	7'h7d :
		RG_rl_105_t1 = TR_117 ;
	7'h7e :
		RG_rl_105_t1 = TR_117 ;
	7'h7f :
		RG_rl_105_t1 = TR_117 ;
	default :
		RG_rl_105_t1 = 9'hx ;
	endcase
always @ ( RG_rl_105_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_46 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_105_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h69 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_105_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_46 )
		| ( { 9{ U_569 } } & RG_rl_105_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_105_en = ( U_570 | RG_rl_105_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_105_en )
		RG_rl_105 <= RG_rl_105_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_118 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_106_t1 = TR_118 ;
	7'h01 :
		RG_rl_106_t1 = TR_118 ;
	7'h02 :
		RG_rl_106_t1 = TR_118 ;
	7'h03 :
		RG_rl_106_t1 = TR_118 ;
	7'h04 :
		RG_rl_106_t1 = TR_118 ;
	7'h05 :
		RG_rl_106_t1 = TR_118 ;
	7'h06 :
		RG_rl_106_t1 = TR_118 ;
	7'h07 :
		RG_rl_106_t1 = TR_118 ;
	7'h08 :
		RG_rl_106_t1 = TR_118 ;
	7'h09 :
		RG_rl_106_t1 = TR_118 ;
	7'h0a :
		RG_rl_106_t1 = TR_118 ;
	7'h0b :
		RG_rl_106_t1 = TR_118 ;
	7'h0c :
		RG_rl_106_t1 = TR_118 ;
	7'h0d :
		RG_rl_106_t1 = TR_118 ;
	7'h0e :
		RG_rl_106_t1 = TR_118 ;
	7'h0f :
		RG_rl_106_t1 = TR_118 ;
	7'h10 :
		RG_rl_106_t1 = TR_118 ;
	7'h11 :
		RG_rl_106_t1 = TR_118 ;
	7'h12 :
		RG_rl_106_t1 = TR_118 ;
	7'h13 :
		RG_rl_106_t1 = TR_118 ;
	7'h14 :
		RG_rl_106_t1 = TR_118 ;
	7'h15 :
		RG_rl_106_t1 = TR_118 ;
	7'h16 :
		RG_rl_106_t1 = TR_118 ;
	7'h17 :
		RG_rl_106_t1 = TR_118 ;
	7'h18 :
		RG_rl_106_t1 = TR_118 ;
	7'h19 :
		RG_rl_106_t1 = TR_118 ;
	7'h1a :
		RG_rl_106_t1 = TR_118 ;
	7'h1b :
		RG_rl_106_t1 = TR_118 ;
	7'h1c :
		RG_rl_106_t1 = TR_118 ;
	7'h1d :
		RG_rl_106_t1 = TR_118 ;
	7'h1e :
		RG_rl_106_t1 = TR_118 ;
	7'h1f :
		RG_rl_106_t1 = TR_118 ;
	7'h20 :
		RG_rl_106_t1 = TR_118 ;
	7'h21 :
		RG_rl_106_t1 = TR_118 ;
	7'h22 :
		RG_rl_106_t1 = TR_118 ;
	7'h23 :
		RG_rl_106_t1 = TR_118 ;
	7'h24 :
		RG_rl_106_t1 = TR_118 ;
	7'h25 :
		RG_rl_106_t1 = TR_118 ;
	7'h26 :
		RG_rl_106_t1 = TR_118 ;
	7'h27 :
		RG_rl_106_t1 = TR_118 ;
	7'h28 :
		RG_rl_106_t1 = TR_118 ;
	7'h29 :
		RG_rl_106_t1 = TR_118 ;
	7'h2a :
		RG_rl_106_t1 = TR_118 ;
	7'h2b :
		RG_rl_106_t1 = TR_118 ;
	7'h2c :
		RG_rl_106_t1 = TR_118 ;
	7'h2d :
		RG_rl_106_t1 = TR_118 ;
	7'h2e :
		RG_rl_106_t1 = TR_118 ;
	7'h2f :
		RG_rl_106_t1 = TR_118 ;
	7'h30 :
		RG_rl_106_t1 = TR_118 ;
	7'h31 :
		RG_rl_106_t1 = TR_118 ;
	7'h32 :
		RG_rl_106_t1 = TR_118 ;
	7'h33 :
		RG_rl_106_t1 = TR_118 ;
	7'h34 :
		RG_rl_106_t1 = TR_118 ;
	7'h35 :
		RG_rl_106_t1 = TR_118 ;
	7'h36 :
		RG_rl_106_t1 = TR_118 ;
	7'h37 :
		RG_rl_106_t1 = TR_118 ;
	7'h38 :
		RG_rl_106_t1 = TR_118 ;
	7'h39 :
		RG_rl_106_t1 = TR_118 ;
	7'h3a :
		RG_rl_106_t1 = TR_118 ;
	7'h3b :
		RG_rl_106_t1 = TR_118 ;
	7'h3c :
		RG_rl_106_t1 = TR_118 ;
	7'h3d :
		RG_rl_106_t1 = TR_118 ;
	7'h3e :
		RG_rl_106_t1 = TR_118 ;
	7'h3f :
		RG_rl_106_t1 = TR_118 ;
	7'h40 :
		RG_rl_106_t1 = TR_118 ;
	7'h41 :
		RG_rl_106_t1 = TR_118 ;
	7'h42 :
		RG_rl_106_t1 = TR_118 ;
	7'h43 :
		RG_rl_106_t1 = TR_118 ;
	7'h44 :
		RG_rl_106_t1 = TR_118 ;
	7'h45 :
		RG_rl_106_t1 = TR_118 ;
	7'h46 :
		RG_rl_106_t1 = TR_118 ;
	7'h47 :
		RG_rl_106_t1 = TR_118 ;
	7'h48 :
		RG_rl_106_t1 = TR_118 ;
	7'h49 :
		RG_rl_106_t1 = TR_118 ;
	7'h4a :
		RG_rl_106_t1 = TR_118 ;
	7'h4b :
		RG_rl_106_t1 = TR_118 ;
	7'h4c :
		RG_rl_106_t1 = TR_118 ;
	7'h4d :
		RG_rl_106_t1 = TR_118 ;
	7'h4e :
		RG_rl_106_t1 = TR_118 ;
	7'h4f :
		RG_rl_106_t1 = TR_118 ;
	7'h50 :
		RG_rl_106_t1 = TR_118 ;
	7'h51 :
		RG_rl_106_t1 = TR_118 ;
	7'h52 :
		RG_rl_106_t1 = TR_118 ;
	7'h53 :
		RG_rl_106_t1 = TR_118 ;
	7'h54 :
		RG_rl_106_t1 = TR_118 ;
	7'h55 :
		RG_rl_106_t1 = TR_118 ;
	7'h56 :
		RG_rl_106_t1 = TR_118 ;
	7'h57 :
		RG_rl_106_t1 = TR_118 ;
	7'h58 :
		RG_rl_106_t1 = TR_118 ;
	7'h59 :
		RG_rl_106_t1 = TR_118 ;
	7'h5a :
		RG_rl_106_t1 = TR_118 ;
	7'h5b :
		RG_rl_106_t1 = TR_118 ;
	7'h5c :
		RG_rl_106_t1 = TR_118 ;
	7'h5d :
		RG_rl_106_t1 = TR_118 ;
	7'h5e :
		RG_rl_106_t1 = TR_118 ;
	7'h5f :
		RG_rl_106_t1 = TR_118 ;
	7'h60 :
		RG_rl_106_t1 = TR_118 ;
	7'h61 :
		RG_rl_106_t1 = TR_118 ;
	7'h62 :
		RG_rl_106_t1 = TR_118 ;
	7'h63 :
		RG_rl_106_t1 = TR_118 ;
	7'h64 :
		RG_rl_106_t1 = TR_118 ;
	7'h65 :
		RG_rl_106_t1 = TR_118 ;
	7'h66 :
		RG_rl_106_t1 = TR_118 ;
	7'h67 :
		RG_rl_106_t1 = TR_118 ;
	7'h68 :
		RG_rl_106_t1 = TR_118 ;
	7'h69 :
		RG_rl_106_t1 = TR_118 ;
	7'h6a :
		RG_rl_106_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6b :
		RG_rl_106_t1 = TR_118 ;
	7'h6c :
		RG_rl_106_t1 = TR_118 ;
	7'h6d :
		RG_rl_106_t1 = TR_118 ;
	7'h6e :
		RG_rl_106_t1 = TR_118 ;
	7'h6f :
		RG_rl_106_t1 = TR_118 ;
	7'h70 :
		RG_rl_106_t1 = TR_118 ;
	7'h71 :
		RG_rl_106_t1 = TR_118 ;
	7'h72 :
		RG_rl_106_t1 = TR_118 ;
	7'h73 :
		RG_rl_106_t1 = TR_118 ;
	7'h74 :
		RG_rl_106_t1 = TR_118 ;
	7'h75 :
		RG_rl_106_t1 = TR_118 ;
	7'h76 :
		RG_rl_106_t1 = TR_118 ;
	7'h77 :
		RG_rl_106_t1 = TR_118 ;
	7'h78 :
		RG_rl_106_t1 = TR_118 ;
	7'h79 :
		RG_rl_106_t1 = TR_118 ;
	7'h7a :
		RG_rl_106_t1 = TR_118 ;
	7'h7b :
		RG_rl_106_t1 = TR_118 ;
	7'h7c :
		RG_rl_106_t1 = TR_118 ;
	7'h7d :
		RG_rl_106_t1 = TR_118 ;
	7'h7e :
		RG_rl_106_t1 = TR_118 ;
	7'h7f :
		RG_rl_106_t1 = TR_118 ;
	default :
		RG_rl_106_t1 = 9'hx ;
	endcase
always @ ( RG_rl_106_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_47 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_106_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h6a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_106_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_47 )
		| ( { 9{ U_569 } } & RG_rl_106_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_106_en = ( U_570 | RG_rl_106_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_106_en )
		RG_rl_106 <= RG_rl_106_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_119 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_107_t1 = TR_119 ;
	7'h01 :
		RG_rl_107_t1 = TR_119 ;
	7'h02 :
		RG_rl_107_t1 = TR_119 ;
	7'h03 :
		RG_rl_107_t1 = TR_119 ;
	7'h04 :
		RG_rl_107_t1 = TR_119 ;
	7'h05 :
		RG_rl_107_t1 = TR_119 ;
	7'h06 :
		RG_rl_107_t1 = TR_119 ;
	7'h07 :
		RG_rl_107_t1 = TR_119 ;
	7'h08 :
		RG_rl_107_t1 = TR_119 ;
	7'h09 :
		RG_rl_107_t1 = TR_119 ;
	7'h0a :
		RG_rl_107_t1 = TR_119 ;
	7'h0b :
		RG_rl_107_t1 = TR_119 ;
	7'h0c :
		RG_rl_107_t1 = TR_119 ;
	7'h0d :
		RG_rl_107_t1 = TR_119 ;
	7'h0e :
		RG_rl_107_t1 = TR_119 ;
	7'h0f :
		RG_rl_107_t1 = TR_119 ;
	7'h10 :
		RG_rl_107_t1 = TR_119 ;
	7'h11 :
		RG_rl_107_t1 = TR_119 ;
	7'h12 :
		RG_rl_107_t1 = TR_119 ;
	7'h13 :
		RG_rl_107_t1 = TR_119 ;
	7'h14 :
		RG_rl_107_t1 = TR_119 ;
	7'h15 :
		RG_rl_107_t1 = TR_119 ;
	7'h16 :
		RG_rl_107_t1 = TR_119 ;
	7'h17 :
		RG_rl_107_t1 = TR_119 ;
	7'h18 :
		RG_rl_107_t1 = TR_119 ;
	7'h19 :
		RG_rl_107_t1 = TR_119 ;
	7'h1a :
		RG_rl_107_t1 = TR_119 ;
	7'h1b :
		RG_rl_107_t1 = TR_119 ;
	7'h1c :
		RG_rl_107_t1 = TR_119 ;
	7'h1d :
		RG_rl_107_t1 = TR_119 ;
	7'h1e :
		RG_rl_107_t1 = TR_119 ;
	7'h1f :
		RG_rl_107_t1 = TR_119 ;
	7'h20 :
		RG_rl_107_t1 = TR_119 ;
	7'h21 :
		RG_rl_107_t1 = TR_119 ;
	7'h22 :
		RG_rl_107_t1 = TR_119 ;
	7'h23 :
		RG_rl_107_t1 = TR_119 ;
	7'h24 :
		RG_rl_107_t1 = TR_119 ;
	7'h25 :
		RG_rl_107_t1 = TR_119 ;
	7'h26 :
		RG_rl_107_t1 = TR_119 ;
	7'h27 :
		RG_rl_107_t1 = TR_119 ;
	7'h28 :
		RG_rl_107_t1 = TR_119 ;
	7'h29 :
		RG_rl_107_t1 = TR_119 ;
	7'h2a :
		RG_rl_107_t1 = TR_119 ;
	7'h2b :
		RG_rl_107_t1 = TR_119 ;
	7'h2c :
		RG_rl_107_t1 = TR_119 ;
	7'h2d :
		RG_rl_107_t1 = TR_119 ;
	7'h2e :
		RG_rl_107_t1 = TR_119 ;
	7'h2f :
		RG_rl_107_t1 = TR_119 ;
	7'h30 :
		RG_rl_107_t1 = TR_119 ;
	7'h31 :
		RG_rl_107_t1 = TR_119 ;
	7'h32 :
		RG_rl_107_t1 = TR_119 ;
	7'h33 :
		RG_rl_107_t1 = TR_119 ;
	7'h34 :
		RG_rl_107_t1 = TR_119 ;
	7'h35 :
		RG_rl_107_t1 = TR_119 ;
	7'h36 :
		RG_rl_107_t1 = TR_119 ;
	7'h37 :
		RG_rl_107_t1 = TR_119 ;
	7'h38 :
		RG_rl_107_t1 = TR_119 ;
	7'h39 :
		RG_rl_107_t1 = TR_119 ;
	7'h3a :
		RG_rl_107_t1 = TR_119 ;
	7'h3b :
		RG_rl_107_t1 = TR_119 ;
	7'h3c :
		RG_rl_107_t1 = TR_119 ;
	7'h3d :
		RG_rl_107_t1 = TR_119 ;
	7'h3e :
		RG_rl_107_t1 = TR_119 ;
	7'h3f :
		RG_rl_107_t1 = TR_119 ;
	7'h40 :
		RG_rl_107_t1 = TR_119 ;
	7'h41 :
		RG_rl_107_t1 = TR_119 ;
	7'h42 :
		RG_rl_107_t1 = TR_119 ;
	7'h43 :
		RG_rl_107_t1 = TR_119 ;
	7'h44 :
		RG_rl_107_t1 = TR_119 ;
	7'h45 :
		RG_rl_107_t1 = TR_119 ;
	7'h46 :
		RG_rl_107_t1 = TR_119 ;
	7'h47 :
		RG_rl_107_t1 = TR_119 ;
	7'h48 :
		RG_rl_107_t1 = TR_119 ;
	7'h49 :
		RG_rl_107_t1 = TR_119 ;
	7'h4a :
		RG_rl_107_t1 = TR_119 ;
	7'h4b :
		RG_rl_107_t1 = TR_119 ;
	7'h4c :
		RG_rl_107_t1 = TR_119 ;
	7'h4d :
		RG_rl_107_t1 = TR_119 ;
	7'h4e :
		RG_rl_107_t1 = TR_119 ;
	7'h4f :
		RG_rl_107_t1 = TR_119 ;
	7'h50 :
		RG_rl_107_t1 = TR_119 ;
	7'h51 :
		RG_rl_107_t1 = TR_119 ;
	7'h52 :
		RG_rl_107_t1 = TR_119 ;
	7'h53 :
		RG_rl_107_t1 = TR_119 ;
	7'h54 :
		RG_rl_107_t1 = TR_119 ;
	7'h55 :
		RG_rl_107_t1 = TR_119 ;
	7'h56 :
		RG_rl_107_t1 = TR_119 ;
	7'h57 :
		RG_rl_107_t1 = TR_119 ;
	7'h58 :
		RG_rl_107_t1 = TR_119 ;
	7'h59 :
		RG_rl_107_t1 = TR_119 ;
	7'h5a :
		RG_rl_107_t1 = TR_119 ;
	7'h5b :
		RG_rl_107_t1 = TR_119 ;
	7'h5c :
		RG_rl_107_t1 = TR_119 ;
	7'h5d :
		RG_rl_107_t1 = TR_119 ;
	7'h5e :
		RG_rl_107_t1 = TR_119 ;
	7'h5f :
		RG_rl_107_t1 = TR_119 ;
	7'h60 :
		RG_rl_107_t1 = TR_119 ;
	7'h61 :
		RG_rl_107_t1 = TR_119 ;
	7'h62 :
		RG_rl_107_t1 = TR_119 ;
	7'h63 :
		RG_rl_107_t1 = TR_119 ;
	7'h64 :
		RG_rl_107_t1 = TR_119 ;
	7'h65 :
		RG_rl_107_t1 = TR_119 ;
	7'h66 :
		RG_rl_107_t1 = TR_119 ;
	7'h67 :
		RG_rl_107_t1 = TR_119 ;
	7'h68 :
		RG_rl_107_t1 = TR_119 ;
	7'h69 :
		RG_rl_107_t1 = TR_119 ;
	7'h6a :
		RG_rl_107_t1 = TR_119 ;
	7'h6b :
		RG_rl_107_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6c :
		RG_rl_107_t1 = TR_119 ;
	7'h6d :
		RG_rl_107_t1 = TR_119 ;
	7'h6e :
		RG_rl_107_t1 = TR_119 ;
	7'h6f :
		RG_rl_107_t1 = TR_119 ;
	7'h70 :
		RG_rl_107_t1 = TR_119 ;
	7'h71 :
		RG_rl_107_t1 = TR_119 ;
	7'h72 :
		RG_rl_107_t1 = TR_119 ;
	7'h73 :
		RG_rl_107_t1 = TR_119 ;
	7'h74 :
		RG_rl_107_t1 = TR_119 ;
	7'h75 :
		RG_rl_107_t1 = TR_119 ;
	7'h76 :
		RG_rl_107_t1 = TR_119 ;
	7'h77 :
		RG_rl_107_t1 = TR_119 ;
	7'h78 :
		RG_rl_107_t1 = TR_119 ;
	7'h79 :
		RG_rl_107_t1 = TR_119 ;
	7'h7a :
		RG_rl_107_t1 = TR_119 ;
	7'h7b :
		RG_rl_107_t1 = TR_119 ;
	7'h7c :
		RG_rl_107_t1 = TR_119 ;
	7'h7d :
		RG_rl_107_t1 = TR_119 ;
	7'h7e :
		RG_rl_107_t1 = TR_119 ;
	7'h7f :
		RG_rl_107_t1 = TR_119 ;
	default :
		RG_rl_107_t1 = 9'hx ;
	endcase
always @ ( RG_rl_107_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_48 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_107_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h6b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_107_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_48 )
		| ( { 9{ U_569 } } & RG_rl_107_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_107_en = ( U_570 | RG_rl_107_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_107_en )
		RG_rl_107 <= RG_rl_107_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_120 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_108_t1 = TR_120 ;
	7'h01 :
		RG_rl_108_t1 = TR_120 ;
	7'h02 :
		RG_rl_108_t1 = TR_120 ;
	7'h03 :
		RG_rl_108_t1 = TR_120 ;
	7'h04 :
		RG_rl_108_t1 = TR_120 ;
	7'h05 :
		RG_rl_108_t1 = TR_120 ;
	7'h06 :
		RG_rl_108_t1 = TR_120 ;
	7'h07 :
		RG_rl_108_t1 = TR_120 ;
	7'h08 :
		RG_rl_108_t1 = TR_120 ;
	7'h09 :
		RG_rl_108_t1 = TR_120 ;
	7'h0a :
		RG_rl_108_t1 = TR_120 ;
	7'h0b :
		RG_rl_108_t1 = TR_120 ;
	7'h0c :
		RG_rl_108_t1 = TR_120 ;
	7'h0d :
		RG_rl_108_t1 = TR_120 ;
	7'h0e :
		RG_rl_108_t1 = TR_120 ;
	7'h0f :
		RG_rl_108_t1 = TR_120 ;
	7'h10 :
		RG_rl_108_t1 = TR_120 ;
	7'h11 :
		RG_rl_108_t1 = TR_120 ;
	7'h12 :
		RG_rl_108_t1 = TR_120 ;
	7'h13 :
		RG_rl_108_t1 = TR_120 ;
	7'h14 :
		RG_rl_108_t1 = TR_120 ;
	7'h15 :
		RG_rl_108_t1 = TR_120 ;
	7'h16 :
		RG_rl_108_t1 = TR_120 ;
	7'h17 :
		RG_rl_108_t1 = TR_120 ;
	7'h18 :
		RG_rl_108_t1 = TR_120 ;
	7'h19 :
		RG_rl_108_t1 = TR_120 ;
	7'h1a :
		RG_rl_108_t1 = TR_120 ;
	7'h1b :
		RG_rl_108_t1 = TR_120 ;
	7'h1c :
		RG_rl_108_t1 = TR_120 ;
	7'h1d :
		RG_rl_108_t1 = TR_120 ;
	7'h1e :
		RG_rl_108_t1 = TR_120 ;
	7'h1f :
		RG_rl_108_t1 = TR_120 ;
	7'h20 :
		RG_rl_108_t1 = TR_120 ;
	7'h21 :
		RG_rl_108_t1 = TR_120 ;
	7'h22 :
		RG_rl_108_t1 = TR_120 ;
	7'h23 :
		RG_rl_108_t1 = TR_120 ;
	7'h24 :
		RG_rl_108_t1 = TR_120 ;
	7'h25 :
		RG_rl_108_t1 = TR_120 ;
	7'h26 :
		RG_rl_108_t1 = TR_120 ;
	7'h27 :
		RG_rl_108_t1 = TR_120 ;
	7'h28 :
		RG_rl_108_t1 = TR_120 ;
	7'h29 :
		RG_rl_108_t1 = TR_120 ;
	7'h2a :
		RG_rl_108_t1 = TR_120 ;
	7'h2b :
		RG_rl_108_t1 = TR_120 ;
	7'h2c :
		RG_rl_108_t1 = TR_120 ;
	7'h2d :
		RG_rl_108_t1 = TR_120 ;
	7'h2e :
		RG_rl_108_t1 = TR_120 ;
	7'h2f :
		RG_rl_108_t1 = TR_120 ;
	7'h30 :
		RG_rl_108_t1 = TR_120 ;
	7'h31 :
		RG_rl_108_t1 = TR_120 ;
	7'h32 :
		RG_rl_108_t1 = TR_120 ;
	7'h33 :
		RG_rl_108_t1 = TR_120 ;
	7'h34 :
		RG_rl_108_t1 = TR_120 ;
	7'h35 :
		RG_rl_108_t1 = TR_120 ;
	7'h36 :
		RG_rl_108_t1 = TR_120 ;
	7'h37 :
		RG_rl_108_t1 = TR_120 ;
	7'h38 :
		RG_rl_108_t1 = TR_120 ;
	7'h39 :
		RG_rl_108_t1 = TR_120 ;
	7'h3a :
		RG_rl_108_t1 = TR_120 ;
	7'h3b :
		RG_rl_108_t1 = TR_120 ;
	7'h3c :
		RG_rl_108_t1 = TR_120 ;
	7'h3d :
		RG_rl_108_t1 = TR_120 ;
	7'h3e :
		RG_rl_108_t1 = TR_120 ;
	7'h3f :
		RG_rl_108_t1 = TR_120 ;
	7'h40 :
		RG_rl_108_t1 = TR_120 ;
	7'h41 :
		RG_rl_108_t1 = TR_120 ;
	7'h42 :
		RG_rl_108_t1 = TR_120 ;
	7'h43 :
		RG_rl_108_t1 = TR_120 ;
	7'h44 :
		RG_rl_108_t1 = TR_120 ;
	7'h45 :
		RG_rl_108_t1 = TR_120 ;
	7'h46 :
		RG_rl_108_t1 = TR_120 ;
	7'h47 :
		RG_rl_108_t1 = TR_120 ;
	7'h48 :
		RG_rl_108_t1 = TR_120 ;
	7'h49 :
		RG_rl_108_t1 = TR_120 ;
	7'h4a :
		RG_rl_108_t1 = TR_120 ;
	7'h4b :
		RG_rl_108_t1 = TR_120 ;
	7'h4c :
		RG_rl_108_t1 = TR_120 ;
	7'h4d :
		RG_rl_108_t1 = TR_120 ;
	7'h4e :
		RG_rl_108_t1 = TR_120 ;
	7'h4f :
		RG_rl_108_t1 = TR_120 ;
	7'h50 :
		RG_rl_108_t1 = TR_120 ;
	7'h51 :
		RG_rl_108_t1 = TR_120 ;
	7'h52 :
		RG_rl_108_t1 = TR_120 ;
	7'h53 :
		RG_rl_108_t1 = TR_120 ;
	7'h54 :
		RG_rl_108_t1 = TR_120 ;
	7'h55 :
		RG_rl_108_t1 = TR_120 ;
	7'h56 :
		RG_rl_108_t1 = TR_120 ;
	7'h57 :
		RG_rl_108_t1 = TR_120 ;
	7'h58 :
		RG_rl_108_t1 = TR_120 ;
	7'h59 :
		RG_rl_108_t1 = TR_120 ;
	7'h5a :
		RG_rl_108_t1 = TR_120 ;
	7'h5b :
		RG_rl_108_t1 = TR_120 ;
	7'h5c :
		RG_rl_108_t1 = TR_120 ;
	7'h5d :
		RG_rl_108_t1 = TR_120 ;
	7'h5e :
		RG_rl_108_t1 = TR_120 ;
	7'h5f :
		RG_rl_108_t1 = TR_120 ;
	7'h60 :
		RG_rl_108_t1 = TR_120 ;
	7'h61 :
		RG_rl_108_t1 = TR_120 ;
	7'h62 :
		RG_rl_108_t1 = TR_120 ;
	7'h63 :
		RG_rl_108_t1 = TR_120 ;
	7'h64 :
		RG_rl_108_t1 = TR_120 ;
	7'h65 :
		RG_rl_108_t1 = TR_120 ;
	7'h66 :
		RG_rl_108_t1 = TR_120 ;
	7'h67 :
		RG_rl_108_t1 = TR_120 ;
	7'h68 :
		RG_rl_108_t1 = TR_120 ;
	7'h69 :
		RG_rl_108_t1 = TR_120 ;
	7'h6a :
		RG_rl_108_t1 = TR_120 ;
	7'h6b :
		RG_rl_108_t1 = TR_120 ;
	7'h6c :
		RG_rl_108_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6d :
		RG_rl_108_t1 = TR_120 ;
	7'h6e :
		RG_rl_108_t1 = TR_120 ;
	7'h6f :
		RG_rl_108_t1 = TR_120 ;
	7'h70 :
		RG_rl_108_t1 = TR_120 ;
	7'h71 :
		RG_rl_108_t1 = TR_120 ;
	7'h72 :
		RG_rl_108_t1 = TR_120 ;
	7'h73 :
		RG_rl_108_t1 = TR_120 ;
	7'h74 :
		RG_rl_108_t1 = TR_120 ;
	7'h75 :
		RG_rl_108_t1 = TR_120 ;
	7'h76 :
		RG_rl_108_t1 = TR_120 ;
	7'h77 :
		RG_rl_108_t1 = TR_120 ;
	7'h78 :
		RG_rl_108_t1 = TR_120 ;
	7'h79 :
		RG_rl_108_t1 = TR_120 ;
	7'h7a :
		RG_rl_108_t1 = TR_120 ;
	7'h7b :
		RG_rl_108_t1 = TR_120 ;
	7'h7c :
		RG_rl_108_t1 = TR_120 ;
	7'h7d :
		RG_rl_108_t1 = TR_120 ;
	7'h7e :
		RG_rl_108_t1 = TR_120 ;
	7'h7f :
		RG_rl_108_t1 = TR_120 ;
	default :
		RG_rl_108_t1 = 9'hx ;
	endcase
always @ ( RG_rl_108_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_49 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_108_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h6c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_108_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_49 )
		| ( { 9{ U_569 } } & RG_rl_108_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_108_en = ( U_570 | RG_rl_108_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_108_en )
		RG_rl_108 <= RG_rl_108_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_121 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_109_t1 = TR_121 ;
	7'h01 :
		RG_rl_109_t1 = TR_121 ;
	7'h02 :
		RG_rl_109_t1 = TR_121 ;
	7'h03 :
		RG_rl_109_t1 = TR_121 ;
	7'h04 :
		RG_rl_109_t1 = TR_121 ;
	7'h05 :
		RG_rl_109_t1 = TR_121 ;
	7'h06 :
		RG_rl_109_t1 = TR_121 ;
	7'h07 :
		RG_rl_109_t1 = TR_121 ;
	7'h08 :
		RG_rl_109_t1 = TR_121 ;
	7'h09 :
		RG_rl_109_t1 = TR_121 ;
	7'h0a :
		RG_rl_109_t1 = TR_121 ;
	7'h0b :
		RG_rl_109_t1 = TR_121 ;
	7'h0c :
		RG_rl_109_t1 = TR_121 ;
	7'h0d :
		RG_rl_109_t1 = TR_121 ;
	7'h0e :
		RG_rl_109_t1 = TR_121 ;
	7'h0f :
		RG_rl_109_t1 = TR_121 ;
	7'h10 :
		RG_rl_109_t1 = TR_121 ;
	7'h11 :
		RG_rl_109_t1 = TR_121 ;
	7'h12 :
		RG_rl_109_t1 = TR_121 ;
	7'h13 :
		RG_rl_109_t1 = TR_121 ;
	7'h14 :
		RG_rl_109_t1 = TR_121 ;
	7'h15 :
		RG_rl_109_t1 = TR_121 ;
	7'h16 :
		RG_rl_109_t1 = TR_121 ;
	7'h17 :
		RG_rl_109_t1 = TR_121 ;
	7'h18 :
		RG_rl_109_t1 = TR_121 ;
	7'h19 :
		RG_rl_109_t1 = TR_121 ;
	7'h1a :
		RG_rl_109_t1 = TR_121 ;
	7'h1b :
		RG_rl_109_t1 = TR_121 ;
	7'h1c :
		RG_rl_109_t1 = TR_121 ;
	7'h1d :
		RG_rl_109_t1 = TR_121 ;
	7'h1e :
		RG_rl_109_t1 = TR_121 ;
	7'h1f :
		RG_rl_109_t1 = TR_121 ;
	7'h20 :
		RG_rl_109_t1 = TR_121 ;
	7'h21 :
		RG_rl_109_t1 = TR_121 ;
	7'h22 :
		RG_rl_109_t1 = TR_121 ;
	7'h23 :
		RG_rl_109_t1 = TR_121 ;
	7'h24 :
		RG_rl_109_t1 = TR_121 ;
	7'h25 :
		RG_rl_109_t1 = TR_121 ;
	7'h26 :
		RG_rl_109_t1 = TR_121 ;
	7'h27 :
		RG_rl_109_t1 = TR_121 ;
	7'h28 :
		RG_rl_109_t1 = TR_121 ;
	7'h29 :
		RG_rl_109_t1 = TR_121 ;
	7'h2a :
		RG_rl_109_t1 = TR_121 ;
	7'h2b :
		RG_rl_109_t1 = TR_121 ;
	7'h2c :
		RG_rl_109_t1 = TR_121 ;
	7'h2d :
		RG_rl_109_t1 = TR_121 ;
	7'h2e :
		RG_rl_109_t1 = TR_121 ;
	7'h2f :
		RG_rl_109_t1 = TR_121 ;
	7'h30 :
		RG_rl_109_t1 = TR_121 ;
	7'h31 :
		RG_rl_109_t1 = TR_121 ;
	7'h32 :
		RG_rl_109_t1 = TR_121 ;
	7'h33 :
		RG_rl_109_t1 = TR_121 ;
	7'h34 :
		RG_rl_109_t1 = TR_121 ;
	7'h35 :
		RG_rl_109_t1 = TR_121 ;
	7'h36 :
		RG_rl_109_t1 = TR_121 ;
	7'h37 :
		RG_rl_109_t1 = TR_121 ;
	7'h38 :
		RG_rl_109_t1 = TR_121 ;
	7'h39 :
		RG_rl_109_t1 = TR_121 ;
	7'h3a :
		RG_rl_109_t1 = TR_121 ;
	7'h3b :
		RG_rl_109_t1 = TR_121 ;
	7'h3c :
		RG_rl_109_t1 = TR_121 ;
	7'h3d :
		RG_rl_109_t1 = TR_121 ;
	7'h3e :
		RG_rl_109_t1 = TR_121 ;
	7'h3f :
		RG_rl_109_t1 = TR_121 ;
	7'h40 :
		RG_rl_109_t1 = TR_121 ;
	7'h41 :
		RG_rl_109_t1 = TR_121 ;
	7'h42 :
		RG_rl_109_t1 = TR_121 ;
	7'h43 :
		RG_rl_109_t1 = TR_121 ;
	7'h44 :
		RG_rl_109_t1 = TR_121 ;
	7'h45 :
		RG_rl_109_t1 = TR_121 ;
	7'h46 :
		RG_rl_109_t1 = TR_121 ;
	7'h47 :
		RG_rl_109_t1 = TR_121 ;
	7'h48 :
		RG_rl_109_t1 = TR_121 ;
	7'h49 :
		RG_rl_109_t1 = TR_121 ;
	7'h4a :
		RG_rl_109_t1 = TR_121 ;
	7'h4b :
		RG_rl_109_t1 = TR_121 ;
	7'h4c :
		RG_rl_109_t1 = TR_121 ;
	7'h4d :
		RG_rl_109_t1 = TR_121 ;
	7'h4e :
		RG_rl_109_t1 = TR_121 ;
	7'h4f :
		RG_rl_109_t1 = TR_121 ;
	7'h50 :
		RG_rl_109_t1 = TR_121 ;
	7'h51 :
		RG_rl_109_t1 = TR_121 ;
	7'h52 :
		RG_rl_109_t1 = TR_121 ;
	7'h53 :
		RG_rl_109_t1 = TR_121 ;
	7'h54 :
		RG_rl_109_t1 = TR_121 ;
	7'h55 :
		RG_rl_109_t1 = TR_121 ;
	7'h56 :
		RG_rl_109_t1 = TR_121 ;
	7'h57 :
		RG_rl_109_t1 = TR_121 ;
	7'h58 :
		RG_rl_109_t1 = TR_121 ;
	7'h59 :
		RG_rl_109_t1 = TR_121 ;
	7'h5a :
		RG_rl_109_t1 = TR_121 ;
	7'h5b :
		RG_rl_109_t1 = TR_121 ;
	7'h5c :
		RG_rl_109_t1 = TR_121 ;
	7'h5d :
		RG_rl_109_t1 = TR_121 ;
	7'h5e :
		RG_rl_109_t1 = TR_121 ;
	7'h5f :
		RG_rl_109_t1 = TR_121 ;
	7'h60 :
		RG_rl_109_t1 = TR_121 ;
	7'h61 :
		RG_rl_109_t1 = TR_121 ;
	7'h62 :
		RG_rl_109_t1 = TR_121 ;
	7'h63 :
		RG_rl_109_t1 = TR_121 ;
	7'h64 :
		RG_rl_109_t1 = TR_121 ;
	7'h65 :
		RG_rl_109_t1 = TR_121 ;
	7'h66 :
		RG_rl_109_t1 = TR_121 ;
	7'h67 :
		RG_rl_109_t1 = TR_121 ;
	7'h68 :
		RG_rl_109_t1 = TR_121 ;
	7'h69 :
		RG_rl_109_t1 = TR_121 ;
	7'h6a :
		RG_rl_109_t1 = TR_121 ;
	7'h6b :
		RG_rl_109_t1 = TR_121 ;
	7'h6c :
		RG_rl_109_t1 = TR_121 ;
	7'h6d :
		RG_rl_109_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6e :
		RG_rl_109_t1 = TR_121 ;
	7'h6f :
		RG_rl_109_t1 = TR_121 ;
	7'h70 :
		RG_rl_109_t1 = TR_121 ;
	7'h71 :
		RG_rl_109_t1 = TR_121 ;
	7'h72 :
		RG_rl_109_t1 = TR_121 ;
	7'h73 :
		RG_rl_109_t1 = TR_121 ;
	7'h74 :
		RG_rl_109_t1 = TR_121 ;
	7'h75 :
		RG_rl_109_t1 = TR_121 ;
	7'h76 :
		RG_rl_109_t1 = TR_121 ;
	7'h77 :
		RG_rl_109_t1 = TR_121 ;
	7'h78 :
		RG_rl_109_t1 = TR_121 ;
	7'h79 :
		RG_rl_109_t1 = TR_121 ;
	7'h7a :
		RG_rl_109_t1 = TR_121 ;
	7'h7b :
		RG_rl_109_t1 = TR_121 ;
	7'h7c :
		RG_rl_109_t1 = TR_121 ;
	7'h7d :
		RG_rl_109_t1 = TR_121 ;
	7'h7e :
		RG_rl_109_t1 = TR_121 ;
	7'h7f :
		RG_rl_109_t1 = TR_121 ;
	default :
		RG_rl_109_t1 = 9'hx ;
	endcase
always @ ( RG_rl_109_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_50 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_109_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h6d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_109_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_50 )
		| ( { 9{ U_569 } } & RG_rl_109_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_109_en = ( U_570 | RG_rl_109_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_109_en )
		RG_rl_109 <= RG_rl_109_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_122 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_110_t1 = TR_122 ;
	7'h01 :
		RG_rl_110_t1 = TR_122 ;
	7'h02 :
		RG_rl_110_t1 = TR_122 ;
	7'h03 :
		RG_rl_110_t1 = TR_122 ;
	7'h04 :
		RG_rl_110_t1 = TR_122 ;
	7'h05 :
		RG_rl_110_t1 = TR_122 ;
	7'h06 :
		RG_rl_110_t1 = TR_122 ;
	7'h07 :
		RG_rl_110_t1 = TR_122 ;
	7'h08 :
		RG_rl_110_t1 = TR_122 ;
	7'h09 :
		RG_rl_110_t1 = TR_122 ;
	7'h0a :
		RG_rl_110_t1 = TR_122 ;
	7'h0b :
		RG_rl_110_t1 = TR_122 ;
	7'h0c :
		RG_rl_110_t1 = TR_122 ;
	7'h0d :
		RG_rl_110_t1 = TR_122 ;
	7'h0e :
		RG_rl_110_t1 = TR_122 ;
	7'h0f :
		RG_rl_110_t1 = TR_122 ;
	7'h10 :
		RG_rl_110_t1 = TR_122 ;
	7'h11 :
		RG_rl_110_t1 = TR_122 ;
	7'h12 :
		RG_rl_110_t1 = TR_122 ;
	7'h13 :
		RG_rl_110_t1 = TR_122 ;
	7'h14 :
		RG_rl_110_t1 = TR_122 ;
	7'h15 :
		RG_rl_110_t1 = TR_122 ;
	7'h16 :
		RG_rl_110_t1 = TR_122 ;
	7'h17 :
		RG_rl_110_t1 = TR_122 ;
	7'h18 :
		RG_rl_110_t1 = TR_122 ;
	7'h19 :
		RG_rl_110_t1 = TR_122 ;
	7'h1a :
		RG_rl_110_t1 = TR_122 ;
	7'h1b :
		RG_rl_110_t1 = TR_122 ;
	7'h1c :
		RG_rl_110_t1 = TR_122 ;
	7'h1d :
		RG_rl_110_t1 = TR_122 ;
	7'h1e :
		RG_rl_110_t1 = TR_122 ;
	7'h1f :
		RG_rl_110_t1 = TR_122 ;
	7'h20 :
		RG_rl_110_t1 = TR_122 ;
	7'h21 :
		RG_rl_110_t1 = TR_122 ;
	7'h22 :
		RG_rl_110_t1 = TR_122 ;
	7'h23 :
		RG_rl_110_t1 = TR_122 ;
	7'h24 :
		RG_rl_110_t1 = TR_122 ;
	7'h25 :
		RG_rl_110_t1 = TR_122 ;
	7'h26 :
		RG_rl_110_t1 = TR_122 ;
	7'h27 :
		RG_rl_110_t1 = TR_122 ;
	7'h28 :
		RG_rl_110_t1 = TR_122 ;
	7'h29 :
		RG_rl_110_t1 = TR_122 ;
	7'h2a :
		RG_rl_110_t1 = TR_122 ;
	7'h2b :
		RG_rl_110_t1 = TR_122 ;
	7'h2c :
		RG_rl_110_t1 = TR_122 ;
	7'h2d :
		RG_rl_110_t1 = TR_122 ;
	7'h2e :
		RG_rl_110_t1 = TR_122 ;
	7'h2f :
		RG_rl_110_t1 = TR_122 ;
	7'h30 :
		RG_rl_110_t1 = TR_122 ;
	7'h31 :
		RG_rl_110_t1 = TR_122 ;
	7'h32 :
		RG_rl_110_t1 = TR_122 ;
	7'h33 :
		RG_rl_110_t1 = TR_122 ;
	7'h34 :
		RG_rl_110_t1 = TR_122 ;
	7'h35 :
		RG_rl_110_t1 = TR_122 ;
	7'h36 :
		RG_rl_110_t1 = TR_122 ;
	7'h37 :
		RG_rl_110_t1 = TR_122 ;
	7'h38 :
		RG_rl_110_t1 = TR_122 ;
	7'h39 :
		RG_rl_110_t1 = TR_122 ;
	7'h3a :
		RG_rl_110_t1 = TR_122 ;
	7'h3b :
		RG_rl_110_t1 = TR_122 ;
	7'h3c :
		RG_rl_110_t1 = TR_122 ;
	7'h3d :
		RG_rl_110_t1 = TR_122 ;
	7'h3e :
		RG_rl_110_t1 = TR_122 ;
	7'h3f :
		RG_rl_110_t1 = TR_122 ;
	7'h40 :
		RG_rl_110_t1 = TR_122 ;
	7'h41 :
		RG_rl_110_t1 = TR_122 ;
	7'h42 :
		RG_rl_110_t1 = TR_122 ;
	7'h43 :
		RG_rl_110_t1 = TR_122 ;
	7'h44 :
		RG_rl_110_t1 = TR_122 ;
	7'h45 :
		RG_rl_110_t1 = TR_122 ;
	7'h46 :
		RG_rl_110_t1 = TR_122 ;
	7'h47 :
		RG_rl_110_t1 = TR_122 ;
	7'h48 :
		RG_rl_110_t1 = TR_122 ;
	7'h49 :
		RG_rl_110_t1 = TR_122 ;
	7'h4a :
		RG_rl_110_t1 = TR_122 ;
	7'h4b :
		RG_rl_110_t1 = TR_122 ;
	7'h4c :
		RG_rl_110_t1 = TR_122 ;
	7'h4d :
		RG_rl_110_t1 = TR_122 ;
	7'h4e :
		RG_rl_110_t1 = TR_122 ;
	7'h4f :
		RG_rl_110_t1 = TR_122 ;
	7'h50 :
		RG_rl_110_t1 = TR_122 ;
	7'h51 :
		RG_rl_110_t1 = TR_122 ;
	7'h52 :
		RG_rl_110_t1 = TR_122 ;
	7'h53 :
		RG_rl_110_t1 = TR_122 ;
	7'h54 :
		RG_rl_110_t1 = TR_122 ;
	7'h55 :
		RG_rl_110_t1 = TR_122 ;
	7'h56 :
		RG_rl_110_t1 = TR_122 ;
	7'h57 :
		RG_rl_110_t1 = TR_122 ;
	7'h58 :
		RG_rl_110_t1 = TR_122 ;
	7'h59 :
		RG_rl_110_t1 = TR_122 ;
	7'h5a :
		RG_rl_110_t1 = TR_122 ;
	7'h5b :
		RG_rl_110_t1 = TR_122 ;
	7'h5c :
		RG_rl_110_t1 = TR_122 ;
	7'h5d :
		RG_rl_110_t1 = TR_122 ;
	7'h5e :
		RG_rl_110_t1 = TR_122 ;
	7'h5f :
		RG_rl_110_t1 = TR_122 ;
	7'h60 :
		RG_rl_110_t1 = TR_122 ;
	7'h61 :
		RG_rl_110_t1 = TR_122 ;
	7'h62 :
		RG_rl_110_t1 = TR_122 ;
	7'h63 :
		RG_rl_110_t1 = TR_122 ;
	7'h64 :
		RG_rl_110_t1 = TR_122 ;
	7'h65 :
		RG_rl_110_t1 = TR_122 ;
	7'h66 :
		RG_rl_110_t1 = TR_122 ;
	7'h67 :
		RG_rl_110_t1 = TR_122 ;
	7'h68 :
		RG_rl_110_t1 = TR_122 ;
	7'h69 :
		RG_rl_110_t1 = TR_122 ;
	7'h6a :
		RG_rl_110_t1 = TR_122 ;
	7'h6b :
		RG_rl_110_t1 = TR_122 ;
	7'h6c :
		RG_rl_110_t1 = TR_122 ;
	7'h6d :
		RG_rl_110_t1 = TR_122 ;
	7'h6e :
		RG_rl_110_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h6f :
		RG_rl_110_t1 = TR_122 ;
	7'h70 :
		RG_rl_110_t1 = TR_122 ;
	7'h71 :
		RG_rl_110_t1 = TR_122 ;
	7'h72 :
		RG_rl_110_t1 = TR_122 ;
	7'h73 :
		RG_rl_110_t1 = TR_122 ;
	7'h74 :
		RG_rl_110_t1 = TR_122 ;
	7'h75 :
		RG_rl_110_t1 = TR_122 ;
	7'h76 :
		RG_rl_110_t1 = TR_122 ;
	7'h77 :
		RG_rl_110_t1 = TR_122 ;
	7'h78 :
		RG_rl_110_t1 = TR_122 ;
	7'h79 :
		RG_rl_110_t1 = TR_122 ;
	7'h7a :
		RG_rl_110_t1 = TR_122 ;
	7'h7b :
		RG_rl_110_t1 = TR_122 ;
	7'h7c :
		RG_rl_110_t1 = TR_122 ;
	7'h7d :
		RG_rl_110_t1 = TR_122 ;
	7'h7e :
		RG_rl_110_t1 = TR_122 ;
	7'h7f :
		RG_rl_110_t1 = TR_122 ;
	default :
		RG_rl_110_t1 = 9'hx ;
	endcase
always @ ( RG_rl_110_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_51 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_110_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h6e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_110_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_51 )
		| ( { 9{ U_569 } } & RG_rl_110_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_110_en = ( U_570 | RG_rl_110_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_110_en )
		RG_rl_110 <= RG_rl_110_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_123 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_111_t1 = TR_123 ;
	7'h01 :
		RG_rl_111_t1 = TR_123 ;
	7'h02 :
		RG_rl_111_t1 = TR_123 ;
	7'h03 :
		RG_rl_111_t1 = TR_123 ;
	7'h04 :
		RG_rl_111_t1 = TR_123 ;
	7'h05 :
		RG_rl_111_t1 = TR_123 ;
	7'h06 :
		RG_rl_111_t1 = TR_123 ;
	7'h07 :
		RG_rl_111_t1 = TR_123 ;
	7'h08 :
		RG_rl_111_t1 = TR_123 ;
	7'h09 :
		RG_rl_111_t1 = TR_123 ;
	7'h0a :
		RG_rl_111_t1 = TR_123 ;
	7'h0b :
		RG_rl_111_t1 = TR_123 ;
	7'h0c :
		RG_rl_111_t1 = TR_123 ;
	7'h0d :
		RG_rl_111_t1 = TR_123 ;
	7'h0e :
		RG_rl_111_t1 = TR_123 ;
	7'h0f :
		RG_rl_111_t1 = TR_123 ;
	7'h10 :
		RG_rl_111_t1 = TR_123 ;
	7'h11 :
		RG_rl_111_t1 = TR_123 ;
	7'h12 :
		RG_rl_111_t1 = TR_123 ;
	7'h13 :
		RG_rl_111_t1 = TR_123 ;
	7'h14 :
		RG_rl_111_t1 = TR_123 ;
	7'h15 :
		RG_rl_111_t1 = TR_123 ;
	7'h16 :
		RG_rl_111_t1 = TR_123 ;
	7'h17 :
		RG_rl_111_t1 = TR_123 ;
	7'h18 :
		RG_rl_111_t1 = TR_123 ;
	7'h19 :
		RG_rl_111_t1 = TR_123 ;
	7'h1a :
		RG_rl_111_t1 = TR_123 ;
	7'h1b :
		RG_rl_111_t1 = TR_123 ;
	7'h1c :
		RG_rl_111_t1 = TR_123 ;
	7'h1d :
		RG_rl_111_t1 = TR_123 ;
	7'h1e :
		RG_rl_111_t1 = TR_123 ;
	7'h1f :
		RG_rl_111_t1 = TR_123 ;
	7'h20 :
		RG_rl_111_t1 = TR_123 ;
	7'h21 :
		RG_rl_111_t1 = TR_123 ;
	7'h22 :
		RG_rl_111_t1 = TR_123 ;
	7'h23 :
		RG_rl_111_t1 = TR_123 ;
	7'h24 :
		RG_rl_111_t1 = TR_123 ;
	7'h25 :
		RG_rl_111_t1 = TR_123 ;
	7'h26 :
		RG_rl_111_t1 = TR_123 ;
	7'h27 :
		RG_rl_111_t1 = TR_123 ;
	7'h28 :
		RG_rl_111_t1 = TR_123 ;
	7'h29 :
		RG_rl_111_t1 = TR_123 ;
	7'h2a :
		RG_rl_111_t1 = TR_123 ;
	7'h2b :
		RG_rl_111_t1 = TR_123 ;
	7'h2c :
		RG_rl_111_t1 = TR_123 ;
	7'h2d :
		RG_rl_111_t1 = TR_123 ;
	7'h2e :
		RG_rl_111_t1 = TR_123 ;
	7'h2f :
		RG_rl_111_t1 = TR_123 ;
	7'h30 :
		RG_rl_111_t1 = TR_123 ;
	7'h31 :
		RG_rl_111_t1 = TR_123 ;
	7'h32 :
		RG_rl_111_t1 = TR_123 ;
	7'h33 :
		RG_rl_111_t1 = TR_123 ;
	7'h34 :
		RG_rl_111_t1 = TR_123 ;
	7'h35 :
		RG_rl_111_t1 = TR_123 ;
	7'h36 :
		RG_rl_111_t1 = TR_123 ;
	7'h37 :
		RG_rl_111_t1 = TR_123 ;
	7'h38 :
		RG_rl_111_t1 = TR_123 ;
	7'h39 :
		RG_rl_111_t1 = TR_123 ;
	7'h3a :
		RG_rl_111_t1 = TR_123 ;
	7'h3b :
		RG_rl_111_t1 = TR_123 ;
	7'h3c :
		RG_rl_111_t1 = TR_123 ;
	7'h3d :
		RG_rl_111_t1 = TR_123 ;
	7'h3e :
		RG_rl_111_t1 = TR_123 ;
	7'h3f :
		RG_rl_111_t1 = TR_123 ;
	7'h40 :
		RG_rl_111_t1 = TR_123 ;
	7'h41 :
		RG_rl_111_t1 = TR_123 ;
	7'h42 :
		RG_rl_111_t1 = TR_123 ;
	7'h43 :
		RG_rl_111_t1 = TR_123 ;
	7'h44 :
		RG_rl_111_t1 = TR_123 ;
	7'h45 :
		RG_rl_111_t1 = TR_123 ;
	7'h46 :
		RG_rl_111_t1 = TR_123 ;
	7'h47 :
		RG_rl_111_t1 = TR_123 ;
	7'h48 :
		RG_rl_111_t1 = TR_123 ;
	7'h49 :
		RG_rl_111_t1 = TR_123 ;
	7'h4a :
		RG_rl_111_t1 = TR_123 ;
	7'h4b :
		RG_rl_111_t1 = TR_123 ;
	7'h4c :
		RG_rl_111_t1 = TR_123 ;
	7'h4d :
		RG_rl_111_t1 = TR_123 ;
	7'h4e :
		RG_rl_111_t1 = TR_123 ;
	7'h4f :
		RG_rl_111_t1 = TR_123 ;
	7'h50 :
		RG_rl_111_t1 = TR_123 ;
	7'h51 :
		RG_rl_111_t1 = TR_123 ;
	7'h52 :
		RG_rl_111_t1 = TR_123 ;
	7'h53 :
		RG_rl_111_t1 = TR_123 ;
	7'h54 :
		RG_rl_111_t1 = TR_123 ;
	7'h55 :
		RG_rl_111_t1 = TR_123 ;
	7'h56 :
		RG_rl_111_t1 = TR_123 ;
	7'h57 :
		RG_rl_111_t1 = TR_123 ;
	7'h58 :
		RG_rl_111_t1 = TR_123 ;
	7'h59 :
		RG_rl_111_t1 = TR_123 ;
	7'h5a :
		RG_rl_111_t1 = TR_123 ;
	7'h5b :
		RG_rl_111_t1 = TR_123 ;
	7'h5c :
		RG_rl_111_t1 = TR_123 ;
	7'h5d :
		RG_rl_111_t1 = TR_123 ;
	7'h5e :
		RG_rl_111_t1 = TR_123 ;
	7'h5f :
		RG_rl_111_t1 = TR_123 ;
	7'h60 :
		RG_rl_111_t1 = TR_123 ;
	7'h61 :
		RG_rl_111_t1 = TR_123 ;
	7'h62 :
		RG_rl_111_t1 = TR_123 ;
	7'h63 :
		RG_rl_111_t1 = TR_123 ;
	7'h64 :
		RG_rl_111_t1 = TR_123 ;
	7'h65 :
		RG_rl_111_t1 = TR_123 ;
	7'h66 :
		RG_rl_111_t1 = TR_123 ;
	7'h67 :
		RG_rl_111_t1 = TR_123 ;
	7'h68 :
		RG_rl_111_t1 = TR_123 ;
	7'h69 :
		RG_rl_111_t1 = TR_123 ;
	7'h6a :
		RG_rl_111_t1 = TR_123 ;
	7'h6b :
		RG_rl_111_t1 = TR_123 ;
	7'h6c :
		RG_rl_111_t1 = TR_123 ;
	7'h6d :
		RG_rl_111_t1 = TR_123 ;
	7'h6e :
		RG_rl_111_t1 = TR_123 ;
	7'h6f :
		RG_rl_111_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h70 :
		RG_rl_111_t1 = TR_123 ;
	7'h71 :
		RG_rl_111_t1 = TR_123 ;
	7'h72 :
		RG_rl_111_t1 = TR_123 ;
	7'h73 :
		RG_rl_111_t1 = TR_123 ;
	7'h74 :
		RG_rl_111_t1 = TR_123 ;
	7'h75 :
		RG_rl_111_t1 = TR_123 ;
	7'h76 :
		RG_rl_111_t1 = TR_123 ;
	7'h77 :
		RG_rl_111_t1 = TR_123 ;
	7'h78 :
		RG_rl_111_t1 = TR_123 ;
	7'h79 :
		RG_rl_111_t1 = TR_123 ;
	7'h7a :
		RG_rl_111_t1 = TR_123 ;
	7'h7b :
		RG_rl_111_t1 = TR_123 ;
	7'h7c :
		RG_rl_111_t1 = TR_123 ;
	7'h7d :
		RG_rl_111_t1 = TR_123 ;
	7'h7e :
		RG_rl_111_t1 = TR_123 ;
	7'h7f :
		RG_rl_111_t1 = TR_123 ;
	default :
		RG_rl_111_t1 = 9'hx ;
	endcase
always @ ( RG_rl_111_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_52 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_111_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h6f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_111_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_52 )
		| ( { 9{ U_569 } } & RG_rl_111_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_111_en = ( U_570 | RG_rl_111_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_111_en )
		RG_rl_111 <= RG_rl_111_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_124 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_112_t1 = TR_124 ;
	7'h01 :
		RG_rl_112_t1 = TR_124 ;
	7'h02 :
		RG_rl_112_t1 = TR_124 ;
	7'h03 :
		RG_rl_112_t1 = TR_124 ;
	7'h04 :
		RG_rl_112_t1 = TR_124 ;
	7'h05 :
		RG_rl_112_t1 = TR_124 ;
	7'h06 :
		RG_rl_112_t1 = TR_124 ;
	7'h07 :
		RG_rl_112_t1 = TR_124 ;
	7'h08 :
		RG_rl_112_t1 = TR_124 ;
	7'h09 :
		RG_rl_112_t1 = TR_124 ;
	7'h0a :
		RG_rl_112_t1 = TR_124 ;
	7'h0b :
		RG_rl_112_t1 = TR_124 ;
	7'h0c :
		RG_rl_112_t1 = TR_124 ;
	7'h0d :
		RG_rl_112_t1 = TR_124 ;
	7'h0e :
		RG_rl_112_t1 = TR_124 ;
	7'h0f :
		RG_rl_112_t1 = TR_124 ;
	7'h10 :
		RG_rl_112_t1 = TR_124 ;
	7'h11 :
		RG_rl_112_t1 = TR_124 ;
	7'h12 :
		RG_rl_112_t1 = TR_124 ;
	7'h13 :
		RG_rl_112_t1 = TR_124 ;
	7'h14 :
		RG_rl_112_t1 = TR_124 ;
	7'h15 :
		RG_rl_112_t1 = TR_124 ;
	7'h16 :
		RG_rl_112_t1 = TR_124 ;
	7'h17 :
		RG_rl_112_t1 = TR_124 ;
	7'h18 :
		RG_rl_112_t1 = TR_124 ;
	7'h19 :
		RG_rl_112_t1 = TR_124 ;
	7'h1a :
		RG_rl_112_t1 = TR_124 ;
	7'h1b :
		RG_rl_112_t1 = TR_124 ;
	7'h1c :
		RG_rl_112_t1 = TR_124 ;
	7'h1d :
		RG_rl_112_t1 = TR_124 ;
	7'h1e :
		RG_rl_112_t1 = TR_124 ;
	7'h1f :
		RG_rl_112_t1 = TR_124 ;
	7'h20 :
		RG_rl_112_t1 = TR_124 ;
	7'h21 :
		RG_rl_112_t1 = TR_124 ;
	7'h22 :
		RG_rl_112_t1 = TR_124 ;
	7'h23 :
		RG_rl_112_t1 = TR_124 ;
	7'h24 :
		RG_rl_112_t1 = TR_124 ;
	7'h25 :
		RG_rl_112_t1 = TR_124 ;
	7'h26 :
		RG_rl_112_t1 = TR_124 ;
	7'h27 :
		RG_rl_112_t1 = TR_124 ;
	7'h28 :
		RG_rl_112_t1 = TR_124 ;
	7'h29 :
		RG_rl_112_t1 = TR_124 ;
	7'h2a :
		RG_rl_112_t1 = TR_124 ;
	7'h2b :
		RG_rl_112_t1 = TR_124 ;
	7'h2c :
		RG_rl_112_t1 = TR_124 ;
	7'h2d :
		RG_rl_112_t1 = TR_124 ;
	7'h2e :
		RG_rl_112_t1 = TR_124 ;
	7'h2f :
		RG_rl_112_t1 = TR_124 ;
	7'h30 :
		RG_rl_112_t1 = TR_124 ;
	7'h31 :
		RG_rl_112_t1 = TR_124 ;
	7'h32 :
		RG_rl_112_t1 = TR_124 ;
	7'h33 :
		RG_rl_112_t1 = TR_124 ;
	7'h34 :
		RG_rl_112_t1 = TR_124 ;
	7'h35 :
		RG_rl_112_t1 = TR_124 ;
	7'h36 :
		RG_rl_112_t1 = TR_124 ;
	7'h37 :
		RG_rl_112_t1 = TR_124 ;
	7'h38 :
		RG_rl_112_t1 = TR_124 ;
	7'h39 :
		RG_rl_112_t1 = TR_124 ;
	7'h3a :
		RG_rl_112_t1 = TR_124 ;
	7'h3b :
		RG_rl_112_t1 = TR_124 ;
	7'h3c :
		RG_rl_112_t1 = TR_124 ;
	7'h3d :
		RG_rl_112_t1 = TR_124 ;
	7'h3e :
		RG_rl_112_t1 = TR_124 ;
	7'h3f :
		RG_rl_112_t1 = TR_124 ;
	7'h40 :
		RG_rl_112_t1 = TR_124 ;
	7'h41 :
		RG_rl_112_t1 = TR_124 ;
	7'h42 :
		RG_rl_112_t1 = TR_124 ;
	7'h43 :
		RG_rl_112_t1 = TR_124 ;
	7'h44 :
		RG_rl_112_t1 = TR_124 ;
	7'h45 :
		RG_rl_112_t1 = TR_124 ;
	7'h46 :
		RG_rl_112_t1 = TR_124 ;
	7'h47 :
		RG_rl_112_t1 = TR_124 ;
	7'h48 :
		RG_rl_112_t1 = TR_124 ;
	7'h49 :
		RG_rl_112_t1 = TR_124 ;
	7'h4a :
		RG_rl_112_t1 = TR_124 ;
	7'h4b :
		RG_rl_112_t1 = TR_124 ;
	7'h4c :
		RG_rl_112_t1 = TR_124 ;
	7'h4d :
		RG_rl_112_t1 = TR_124 ;
	7'h4e :
		RG_rl_112_t1 = TR_124 ;
	7'h4f :
		RG_rl_112_t1 = TR_124 ;
	7'h50 :
		RG_rl_112_t1 = TR_124 ;
	7'h51 :
		RG_rl_112_t1 = TR_124 ;
	7'h52 :
		RG_rl_112_t1 = TR_124 ;
	7'h53 :
		RG_rl_112_t1 = TR_124 ;
	7'h54 :
		RG_rl_112_t1 = TR_124 ;
	7'h55 :
		RG_rl_112_t1 = TR_124 ;
	7'h56 :
		RG_rl_112_t1 = TR_124 ;
	7'h57 :
		RG_rl_112_t1 = TR_124 ;
	7'h58 :
		RG_rl_112_t1 = TR_124 ;
	7'h59 :
		RG_rl_112_t1 = TR_124 ;
	7'h5a :
		RG_rl_112_t1 = TR_124 ;
	7'h5b :
		RG_rl_112_t1 = TR_124 ;
	7'h5c :
		RG_rl_112_t1 = TR_124 ;
	7'h5d :
		RG_rl_112_t1 = TR_124 ;
	7'h5e :
		RG_rl_112_t1 = TR_124 ;
	7'h5f :
		RG_rl_112_t1 = TR_124 ;
	7'h60 :
		RG_rl_112_t1 = TR_124 ;
	7'h61 :
		RG_rl_112_t1 = TR_124 ;
	7'h62 :
		RG_rl_112_t1 = TR_124 ;
	7'h63 :
		RG_rl_112_t1 = TR_124 ;
	7'h64 :
		RG_rl_112_t1 = TR_124 ;
	7'h65 :
		RG_rl_112_t1 = TR_124 ;
	7'h66 :
		RG_rl_112_t1 = TR_124 ;
	7'h67 :
		RG_rl_112_t1 = TR_124 ;
	7'h68 :
		RG_rl_112_t1 = TR_124 ;
	7'h69 :
		RG_rl_112_t1 = TR_124 ;
	7'h6a :
		RG_rl_112_t1 = TR_124 ;
	7'h6b :
		RG_rl_112_t1 = TR_124 ;
	7'h6c :
		RG_rl_112_t1 = TR_124 ;
	7'h6d :
		RG_rl_112_t1 = TR_124 ;
	7'h6e :
		RG_rl_112_t1 = TR_124 ;
	7'h6f :
		RG_rl_112_t1 = TR_124 ;
	7'h70 :
		RG_rl_112_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h71 :
		RG_rl_112_t1 = TR_124 ;
	7'h72 :
		RG_rl_112_t1 = TR_124 ;
	7'h73 :
		RG_rl_112_t1 = TR_124 ;
	7'h74 :
		RG_rl_112_t1 = TR_124 ;
	7'h75 :
		RG_rl_112_t1 = TR_124 ;
	7'h76 :
		RG_rl_112_t1 = TR_124 ;
	7'h77 :
		RG_rl_112_t1 = TR_124 ;
	7'h78 :
		RG_rl_112_t1 = TR_124 ;
	7'h79 :
		RG_rl_112_t1 = TR_124 ;
	7'h7a :
		RG_rl_112_t1 = TR_124 ;
	7'h7b :
		RG_rl_112_t1 = TR_124 ;
	7'h7c :
		RG_rl_112_t1 = TR_124 ;
	7'h7d :
		RG_rl_112_t1 = TR_124 ;
	7'h7e :
		RG_rl_112_t1 = TR_124 ;
	7'h7f :
		RG_rl_112_t1 = TR_124 ;
	default :
		RG_rl_112_t1 = 9'hx ;
	endcase
always @ ( RG_rl_112_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_53 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_112_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h70 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_112_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_53 )
		| ( { 9{ U_569 } } & RG_rl_112_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_112_en = ( U_570 | RG_rl_112_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_112_en )
		RG_rl_112 <= RG_rl_112_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_125 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_113_t1 = TR_125 ;
	7'h01 :
		RG_rl_113_t1 = TR_125 ;
	7'h02 :
		RG_rl_113_t1 = TR_125 ;
	7'h03 :
		RG_rl_113_t1 = TR_125 ;
	7'h04 :
		RG_rl_113_t1 = TR_125 ;
	7'h05 :
		RG_rl_113_t1 = TR_125 ;
	7'h06 :
		RG_rl_113_t1 = TR_125 ;
	7'h07 :
		RG_rl_113_t1 = TR_125 ;
	7'h08 :
		RG_rl_113_t1 = TR_125 ;
	7'h09 :
		RG_rl_113_t1 = TR_125 ;
	7'h0a :
		RG_rl_113_t1 = TR_125 ;
	7'h0b :
		RG_rl_113_t1 = TR_125 ;
	7'h0c :
		RG_rl_113_t1 = TR_125 ;
	7'h0d :
		RG_rl_113_t1 = TR_125 ;
	7'h0e :
		RG_rl_113_t1 = TR_125 ;
	7'h0f :
		RG_rl_113_t1 = TR_125 ;
	7'h10 :
		RG_rl_113_t1 = TR_125 ;
	7'h11 :
		RG_rl_113_t1 = TR_125 ;
	7'h12 :
		RG_rl_113_t1 = TR_125 ;
	7'h13 :
		RG_rl_113_t1 = TR_125 ;
	7'h14 :
		RG_rl_113_t1 = TR_125 ;
	7'h15 :
		RG_rl_113_t1 = TR_125 ;
	7'h16 :
		RG_rl_113_t1 = TR_125 ;
	7'h17 :
		RG_rl_113_t1 = TR_125 ;
	7'h18 :
		RG_rl_113_t1 = TR_125 ;
	7'h19 :
		RG_rl_113_t1 = TR_125 ;
	7'h1a :
		RG_rl_113_t1 = TR_125 ;
	7'h1b :
		RG_rl_113_t1 = TR_125 ;
	7'h1c :
		RG_rl_113_t1 = TR_125 ;
	7'h1d :
		RG_rl_113_t1 = TR_125 ;
	7'h1e :
		RG_rl_113_t1 = TR_125 ;
	7'h1f :
		RG_rl_113_t1 = TR_125 ;
	7'h20 :
		RG_rl_113_t1 = TR_125 ;
	7'h21 :
		RG_rl_113_t1 = TR_125 ;
	7'h22 :
		RG_rl_113_t1 = TR_125 ;
	7'h23 :
		RG_rl_113_t1 = TR_125 ;
	7'h24 :
		RG_rl_113_t1 = TR_125 ;
	7'h25 :
		RG_rl_113_t1 = TR_125 ;
	7'h26 :
		RG_rl_113_t1 = TR_125 ;
	7'h27 :
		RG_rl_113_t1 = TR_125 ;
	7'h28 :
		RG_rl_113_t1 = TR_125 ;
	7'h29 :
		RG_rl_113_t1 = TR_125 ;
	7'h2a :
		RG_rl_113_t1 = TR_125 ;
	7'h2b :
		RG_rl_113_t1 = TR_125 ;
	7'h2c :
		RG_rl_113_t1 = TR_125 ;
	7'h2d :
		RG_rl_113_t1 = TR_125 ;
	7'h2e :
		RG_rl_113_t1 = TR_125 ;
	7'h2f :
		RG_rl_113_t1 = TR_125 ;
	7'h30 :
		RG_rl_113_t1 = TR_125 ;
	7'h31 :
		RG_rl_113_t1 = TR_125 ;
	7'h32 :
		RG_rl_113_t1 = TR_125 ;
	7'h33 :
		RG_rl_113_t1 = TR_125 ;
	7'h34 :
		RG_rl_113_t1 = TR_125 ;
	7'h35 :
		RG_rl_113_t1 = TR_125 ;
	7'h36 :
		RG_rl_113_t1 = TR_125 ;
	7'h37 :
		RG_rl_113_t1 = TR_125 ;
	7'h38 :
		RG_rl_113_t1 = TR_125 ;
	7'h39 :
		RG_rl_113_t1 = TR_125 ;
	7'h3a :
		RG_rl_113_t1 = TR_125 ;
	7'h3b :
		RG_rl_113_t1 = TR_125 ;
	7'h3c :
		RG_rl_113_t1 = TR_125 ;
	7'h3d :
		RG_rl_113_t1 = TR_125 ;
	7'h3e :
		RG_rl_113_t1 = TR_125 ;
	7'h3f :
		RG_rl_113_t1 = TR_125 ;
	7'h40 :
		RG_rl_113_t1 = TR_125 ;
	7'h41 :
		RG_rl_113_t1 = TR_125 ;
	7'h42 :
		RG_rl_113_t1 = TR_125 ;
	7'h43 :
		RG_rl_113_t1 = TR_125 ;
	7'h44 :
		RG_rl_113_t1 = TR_125 ;
	7'h45 :
		RG_rl_113_t1 = TR_125 ;
	7'h46 :
		RG_rl_113_t1 = TR_125 ;
	7'h47 :
		RG_rl_113_t1 = TR_125 ;
	7'h48 :
		RG_rl_113_t1 = TR_125 ;
	7'h49 :
		RG_rl_113_t1 = TR_125 ;
	7'h4a :
		RG_rl_113_t1 = TR_125 ;
	7'h4b :
		RG_rl_113_t1 = TR_125 ;
	7'h4c :
		RG_rl_113_t1 = TR_125 ;
	7'h4d :
		RG_rl_113_t1 = TR_125 ;
	7'h4e :
		RG_rl_113_t1 = TR_125 ;
	7'h4f :
		RG_rl_113_t1 = TR_125 ;
	7'h50 :
		RG_rl_113_t1 = TR_125 ;
	7'h51 :
		RG_rl_113_t1 = TR_125 ;
	7'h52 :
		RG_rl_113_t1 = TR_125 ;
	7'h53 :
		RG_rl_113_t1 = TR_125 ;
	7'h54 :
		RG_rl_113_t1 = TR_125 ;
	7'h55 :
		RG_rl_113_t1 = TR_125 ;
	7'h56 :
		RG_rl_113_t1 = TR_125 ;
	7'h57 :
		RG_rl_113_t1 = TR_125 ;
	7'h58 :
		RG_rl_113_t1 = TR_125 ;
	7'h59 :
		RG_rl_113_t1 = TR_125 ;
	7'h5a :
		RG_rl_113_t1 = TR_125 ;
	7'h5b :
		RG_rl_113_t1 = TR_125 ;
	7'h5c :
		RG_rl_113_t1 = TR_125 ;
	7'h5d :
		RG_rl_113_t1 = TR_125 ;
	7'h5e :
		RG_rl_113_t1 = TR_125 ;
	7'h5f :
		RG_rl_113_t1 = TR_125 ;
	7'h60 :
		RG_rl_113_t1 = TR_125 ;
	7'h61 :
		RG_rl_113_t1 = TR_125 ;
	7'h62 :
		RG_rl_113_t1 = TR_125 ;
	7'h63 :
		RG_rl_113_t1 = TR_125 ;
	7'h64 :
		RG_rl_113_t1 = TR_125 ;
	7'h65 :
		RG_rl_113_t1 = TR_125 ;
	7'h66 :
		RG_rl_113_t1 = TR_125 ;
	7'h67 :
		RG_rl_113_t1 = TR_125 ;
	7'h68 :
		RG_rl_113_t1 = TR_125 ;
	7'h69 :
		RG_rl_113_t1 = TR_125 ;
	7'h6a :
		RG_rl_113_t1 = TR_125 ;
	7'h6b :
		RG_rl_113_t1 = TR_125 ;
	7'h6c :
		RG_rl_113_t1 = TR_125 ;
	7'h6d :
		RG_rl_113_t1 = TR_125 ;
	7'h6e :
		RG_rl_113_t1 = TR_125 ;
	7'h6f :
		RG_rl_113_t1 = TR_125 ;
	7'h70 :
		RG_rl_113_t1 = TR_125 ;
	7'h71 :
		RG_rl_113_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h72 :
		RG_rl_113_t1 = TR_125 ;
	7'h73 :
		RG_rl_113_t1 = TR_125 ;
	7'h74 :
		RG_rl_113_t1 = TR_125 ;
	7'h75 :
		RG_rl_113_t1 = TR_125 ;
	7'h76 :
		RG_rl_113_t1 = TR_125 ;
	7'h77 :
		RG_rl_113_t1 = TR_125 ;
	7'h78 :
		RG_rl_113_t1 = TR_125 ;
	7'h79 :
		RG_rl_113_t1 = TR_125 ;
	7'h7a :
		RG_rl_113_t1 = TR_125 ;
	7'h7b :
		RG_rl_113_t1 = TR_125 ;
	7'h7c :
		RG_rl_113_t1 = TR_125 ;
	7'h7d :
		RG_rl_113_t1 = TR_125 ;
	7'h7e :
		RG_rl_113_t1 = TR_125 ;
	7'h7f :
		RG_rl_113_t1 = TR_125 ;
	default :
		RG_rl_113_t1 = 9'hx ;
	endcase
always @ ( RG_rl_113_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_54 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_113_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h71 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_113_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_54 )
		| ( { 9{ U_569 } } & RG_rl_113_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_113_en = ( U_570 | RG_rl_113_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_113_en )
		RG_rl_113 <= RG_rl_113_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_126 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_114_t1 = TR_126 ;
	7'h01 :
		RG_rl_114_t1 = TR_126 ;
	7'h02 :
		RG_rl_114_t1 = TR_126 ;
	7'h03 :
		RG_rl_114_t1 = TR_126 ;
	7'h04 :
		RG_rl_114_t1 = TR_126 ;
	7'h05 :
		RG_rl_114_t1 = TR_126 ;
	7'h06 :
		RG_rl_114_t1 = TR_126 ;
	7'h07 :
		RG_rl_114_t1 = TR_126 ;
	7'h08 :
		RG_rl_114_t1 = TR_126 ;
	7'h09 :
		RG_rl_114_t1 = TR_126 ;
	7'h0a :
		RG_rl_114_t1 = TR_126 ;
	7'h0b :
		RG_rl_114_t1 = TR_126 ;
	7'h0c :
		RG_rl_114_t1 = TR_126 ;
	7'h0d :
		RG_rl_114_t1 = TR_126 ;
	7'h0e :
		RG_rl_114_t1 = TR_126 ;
	7'h0f :
		RG_rl_114_t1 = TR_126 ;
	7'h10 :
		RG_rl_114_t1 = TR_126 ;
	7'h11 :
		RG_rl_114_t1 = TR_126 ;
	7'h12 :
		RG_rl_114_t1 = TR_126 ;
	7'h13 :
		RG_rl_114_t1 = TR_126 ;
	7'h14 :
		RG_rl_114_t1 = TR_126 ;
	7'h15 :
		RG_rl_114_t1 = TR_126 ;
	7'h16 :
		RG_rl_114_t1 = TR_126 ;
	7'h17 :
		RG_rl_114_t1 = TR_126 ;
	7'h18 :
		RG_rl_114_t1 = TR_126 ;
	7'h19 :
		RG_rl_114_t1 = TR_126 ;
	7'h1a :
		RG_rl_114_t1 = TR_126 ;
	7'h1b :
		RG_rl_114_t1 = TR_126 ;
	7'h1c :
		RG_rl_114_t1 = TR_126 ;
	7'h1d :
		RG_rl_114_t1 = TR_126 ;
	7'h1e :
		RG_rl_114_t1 = TR_126 ;
	7'h1f :
		RG_rl_114_t1 = TR_126 ;
	7'h20 :
		RG_rl_114_t1 = TR_126 ;
	7'h21 :
		RG_rl_114_t1 = TR_126 ;
	7'h22 :
		RG_rl_114_t1 = TR_126 ;
	7'h23 :
		RG_rl_114_t1 = TR_126 ;
	7'h24 :
		RG_rl_114_t1 = TR_126 ;
	7'h25 :
		RG_rl_114_t1 = TR_126 ;
	7'h26 :
		RG_rl_114_t1 = TR_126 ;
	7'h27 :
		RG_rl_114_t1 = TR_126 ;
	7'h28 :
		RG_rl_114_t1 = TR_126 ;
	7'h29 :
		RG_rl_114_t1 = TR_126 ;
	7'h2a :
		RG_rl_114_t1 = TR_126 ;
	7'h2b :
		RG_rl_114_t1 = TR_126 ;
	7'h2c :
		RG_rl_114_t1 = TR_126 ;
	7'h2d :
		RG_rl_114_t1 = TR_126 ;
	7'h2e :
		RG_rl_114_t1 = TR_126 ;
	7'h2f :
		RG_rl_114_t1 = TR_126 ;
	7'h30 :
		RG_rl_114_t1 = TR_126 ;
	7'h31 :
		RG_rl_114_t1 = TR_126 ;
	7'h32 :
		RG_rl_114_t1 = TR_126 ;
	7'h33 :
		RG_rl_114_t1 = TR_126 ;
	7'h34 :
		RG_rl_114_t1 = TR_126 ;
	7'h35 :
		RG_rl_114_t1 = TR_126 ;
	7'h36 :
		RG_rl_114_t1 = TR_126 ;
	7'h37 :
		RG_rl_114_t1 = TR_126 ;
	7'h38 :
		RG_rl_114_t1 = TR_126 ;
	7'h39 :
		RG_rl_114_t1 = TR_126 ;
	7'h3a :
		RG_rl_114_t1 = TR_126 ;
	7'h3b :
		RG_rl_114_t1 = TR_126 ;
	7'h3c :
		RG_rl_114_t1 = TR_126 ;
	7'h3d :
		RG_rl_114_t1 = TR_126 ;
	7'h3e :
		RG_rl_114_t1 = TR_126 ;
	7'h3f :
		RG_rl_114_t1 = TR_126 ;
	7'h40 :
		RG_rl_114_t1 = TR_126 ;
	7'h41 :
		RG_rl_114_t1 = TR_126 ;
	7'h42 :
		RG_rl_114_t1 = TR_126 ;
	7'h43 :
		RG_rl_114_t1 = TR_126 ;
	7'h44 :
		RG_rl_114_t1 = TR_126 ;
	7'h45 :
		RG_rl_114_t1 = TR_126 ;
	7'h46 :
		RG_rl_114_t1 = TR_126 ;
	7'h47 :
		RG_rl_114_t1 = TR_126 ;
	7'h48 :
		RG_rl_114_t1 = TR_126 ;
	7'h49 :
		RG_rl_114_t1 = TR_126 ;
	7'h4a :
		RG_rl_114_t1 = TR_126 ;
	7'h4b :
		RG_rl_114_t1 = TR_126 ;
	7'h4c :
		RG_rl_114_t1 = TR_126 ;
	7'h4d :
		RG_rl_114_t1 = TR_126 ;
	7'h4e :
		RG_rl_114_t1 = TR_126 ;
	7'h4f :
		RG_rl_114_t1 = TR_126 ;
	7'h50 :
		RG_rl_114_t1 = TR_126 ;
	7'h51 :
		RG_rl_114_t1 = TR_126 ;
	7'h52 :
		RG_rl_114_t1 = TR_126 ;
	7'h53 :
		RG_rl_114_t1 = TR_126 ;
	7'h54 :
		RG_rl_114_t1 = TR_126 ;
	7'h55 :
		RG_rl_114_t1 = TR_126 ;
	7'h56 :
		RG_rl_114_t1 = TR_126 ;
	7'h57 :
		RG_rl_114_t1 = TR_126 ;
	7'h58 :
		RG_rl_114_t1 = TR_126 ;
	7'h59 :
		RG_rl_114_t1 = TR_126 ;
	7'h5a :
		RG_rl_114_t1 = TR_126 ;
	7'h5b :
		RG_rl_114_t1 = TR_126 ;
	7'h5c :
		RG_rl_114_t1 = TR_126 ;
	7'h5d :
		RG_rl_114_t1 = TR_126 ;
	7'h5e :
		RG_rl_114_t1 = TR_126 ;
	7'h5f :
		RG_rl_114_t1 = TR_126 ;
	7'h60 :
		RG_rl_114_t1 = TR_126 ;
	7'h61 :
		RG_rl_114_t1 = TR_126 ;
	7'h62 :
		RG_rl_114_t1 = TR_126 ;
	7'h63 :
		RG_rl_114_t1 = TR_126 ;
	7'h64 :
		RG_rl_114_t1 = TR_126 ;
	7'h65 :
		RG_rl_114_t1 = TR_126 ;
	7'h66 :
		RG_rl_114_t1 = TR_126 ;
	7'h67 :
		RG_rl_114_t1 = TR_126 ;
	7'h68 :
		RG_rl_114_t1 = TR_126 ;
	7'h69 :
		RG_rl_114_t1 = TR_126 ;
	7'h6a :
		RG_rl_114_t1 = TR_126 ;
	7'h6b :
		RG_rl_114_t1 = TR_126 ;
	7'h6c :
		RG_rl_114_t1 = TR_126 ;
	7'h6d :
		RG_rl_114_t1 = TR_126 ;
	7'h6e :
		RG_rl_114_t1 = TR_126 ;
	7'h6f :
		RG_rl_114_t1 = TR_126 ;
	7'h70 :
		RG_rl_114_t1 = TR_126 ;
	7'h71 :
		RG_rl_114_t1 = TR_126 ;
	7'h72 :
		RG_rl_114_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h73 :
		RG_rl_114_t1 = TR_126 ;
	7'h74 :
		RG_rl_114_t1 = TR_126 ;
	7'h75 :
		RG_rl_114_t1 = TR_126 ;
	7'h76 :
		RG_rl_114_t1 = TR_126 ;
	7'h77 :
		RG_rl_114_t1 = TR_126 ;
	7'h78 :
		RG_rl_114_t1 = TR_126 ;
	7'h79 :
		RG_rl_114_t1 = TR_126 ;
	7'h7a :
		RG_rl_114_t1 = TR_126 ;
	7'h7b :
		RG_rl_114_t1 = TR_126 ;
	7'h7c :
		RG_rl_114_t1 = TR_126 ;
	7'h7d :
		RG_rl_114_t1 = TR_126 ;
	7'h7e :
		RG_rl_114_t1 = TR_126 ;
	7'h7f :
		RG_rl_114_t1 = TR_126 ;
	default :
		RG_rl_114_t1 = 9'hx ;
	endcase
always @ ( RG_rl_114_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_55 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_114_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h72 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_114_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_55 )
		| ( { 9{ U_569 } } & RG_rl_114_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_114_en = ( U_570 | RG_rl_114_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_114_en )
		RG_rl_114 <= RG_rl_114_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_127 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_115_t1 = TR_127 ;
	7'h01 :
		RG_rl_115_t1 = TR_127 ;
	7'h02 :
		RG_rl_115_t1 = TR_127 ;
	7'h03 :
		RG_rl_115_t1 = TR_127 ;
	7'h04 :
		RG_rl_115_t1 = TR_127 ;
	7'h05 :
		RG_rl_115_t1 = TR_127 ;
	7'h06 :
		RG_rl_115_t1 = TR_127 ;
	7'h07 :
		RG_rl_115_t1 = TR_127 ;
	7'h08 :
		RG_rl_115_t1 = TR_127 ;
	7'h09 :
		RG_rl_115_t1 = TR_127 ;
	7'h0a :
		RG_rl_115_t1 = TR_127 ;
	7'h0b :
		RG_rl_115_t1 = TR_127 ;
	7'h0c :
		RG_rl_115_t1 = TR_127 ;
	7'h0d :
		RG_rl_115_t1 = TR_127 ;
	7'h0e :
		RG_rl_115_t1 = TR_127 ;
	7'h0f :
		RG_rl_115_t1 = TR_127 ;
	7'h10 :
		RG_rl_115_t1 = TR_127 ;
	7'h11 :
		RG_rl_115_t1 = TR_127 ;
	7'h12 :
		RG_rl_115_t1 = TR_127 ;
	7'h13 :
		RG_rl_115_t1 = TR_127 ;
	7'h14 :
		RG_rl_115_t1 = TR_127 ;
	7'h15 :
		RG_rl_115_t1 = TR_127 ;
	7'h16 :
		RG_rl_115_t1 = TR_127 ;
	7'h17 :
		RG_rl_115_t1 = TR_127 ;
	7'h18 :
		RG_rl_115_t1 = TR_127 ;
	7'h19 :
		RG_rl_115_t1 = TR_127 ;
	7'h1a :
		RG_rl_115_t1 = TR_127 ;
	7'h1b :
		RG_rl_115_t1 = TR_127 ;
	7'h1c :
		RG_rl_115_t1 = TR_127 ;
	7'h1d :
		RG_rl_115_t1 = TR_127 ;
	7'h1e :
		RG_rl_115_t1 = TR_127 ;
	7'h1f :
		RG_rl_115_t1 = TR_127 ;
	7'h20 :
		RG_rl_115_t1 = TR_127 ;
	7'h21 :
		RG_rl_115_t1 = TR_127 ;
	7'h22 :
		RG_rl_115_t1 = TR_127 ;
	7'h23 :
		RG_rl_115_t1 = TR_127 ;
	7'h24 :
		RG_rl_115_t1 = TR_127 ;
	7'h25 :
		RG_rl_115_t1 = TR_127 ;
	7'h26 :
		RG_rl_115_t1 = TR_127 ;
	7'h27 :
		RG_rl_115_t1 = TR_127 ;
	7'h28 :
		RG_rl_115_t1 = TR_127 ;
	7'h29 :
		RG_rl_115_t1 = TR_127 ;
	7'h2a :
		RG_rl_115_t1 = TR_127 ;
	7'h2b :
		RG_rl_115_t1 = TR_127 ;
	7'h2c :
		RG_rl_115_t1 = TR_127 ;
	7'h2d :
		RG_rl_115_t1 = TR_127 ;
	7'h2e :
		RG_rl_115_t1 = TR_127 ;
	7'h2f :
		RG_rl_115_t1 = TR_127 ;
	7'h30 :
		RG_rl_115_t1 = TR_127 ;
	7'h31 :
		RG_rl_115_t1 = TR_127 ;
	7'h32 :
		RG_rl_115_t1 = TR_127 ;
	7'h33 :
		RG_rl_115_t1 = TR_127 ;
	7'h34 :
		RG_rl_115_t1 = TR_127 ;
	7'h35 :
		RG_rl_115_t1 = TR_127 ;
	7'h36 :
		RG_rl_115_t1 = TR_127 ;
	7'h37 :
		RG_rl_115_t1 = TR_127 ;
	7'h38 :
		RG_rl_115_t1 = TR_127 ;
	7'h39 :
		RG_rl_115_t1 = TR_127 ;
	7'h3a :
		RG_rl_115_t1 = TR_127 ;
	7'h3b :
		RG_rl_115_t1 = TR_127 ;
	7'h3c :
		RG_rl_115_t1 = TR_127 ;
	7'h3d :
		RG_rl_115_t1 = TR_127 ;
	7'h3e :
		RG_rl_115_t1 = TR_127 ;
	7'h3f :
		RG_rl_115_t1 = TR_127 ;
	7'h40 :
		RG_rl_115_t1 = TR_127 ;
	7'h41 :
		RG_rl_115_t1 = TR_127 ;
	7'h42 :
		RG_rl_115_t1 = TR_127 ;
	7'h43 :
		RG_rl_115_t1 = TR_127 ;
	7'h44 :
		RG_rl_115_t1 = TR_127 ;
	7'h45 :
		RG_rl_115_t1 = TR_127 ;
	7'h46 :
		RG_rl_115_t1 = TR_127 ;
	7'h47 :
		RG_rl_115_t1 = TR_127 ;
	7'h48 :
		RG_rl_115_t1 = TR_127 ;
	7'h49 :
		RG_rl_115_t1 = TR_127 ;
	7'h4a :
		RG_rl_115_t1 = TR_127 ;
	7'h4b :
		RG_rl_115_t1 = TR_127 ;
	7'h4c :
		RG_rl_115_t1 = TR_127 ;
	7'h4d :
		RG_rl_115_t1 = TR_127 ;
	7'h4e :
		RG_rl_115_t1 = TR_127 ;
	7'h4f :
		RG_rl_115_t1 = TR_127 ;
	7'h50 :
		RG_rl_115_t1 = TR_127 ;
	7'h51 :
		RG_rl_115_t1 = TR_127 ;
	7'h52 :
		RG_rl_115_t1 = TR_127 ;
	7'h53 :
		RG_rl_115_t1 = TR_127 ;
	7'h54 :
		RG_rl_115_t1 = TR_127 ;
	7'h55 :
		RG_rl_115_t1 = TR_127 ;
	7'h56 :
		RG_rl_115_t1 = TR_127 ;
	7'h57 :
		RG_rl_115_t1 = TR_127 ;
	7'h58 :
		RG_rl_115_t1 = TR_127 ;
	7'h59 :
		RG_rl_115_t1 = TR_127 ;
	7'h5a :
		RG_rl_115_t1 = TR_127 ;
	7'h5b :
		RG_rl_115_t1 = TR_127 ;
	7'h5c :
		RG_rl_115_t1 = TR_127 ;
	7'h5d :
		RG_rl_115_t1 = TR_127 ;
	7'h5e :
		RG_rl_115_t1 = TR_127 ;
	7'h5f :
		RG_rl_115_t1 = TR_127 ;
	7'h60 :
		RG_rl_115_t1 = TR_127 ;
	7'h61 :
		RG_rl_115_t1 = TR_127 ;
	7'h62 :
		RG_rl_115_t1 = TR_127 ;
	7'h63 :
		RG_rl_115_t1 = TR_127 ;
	7'h64 :
		RG_rl_115_t1 = TR_127 ;
	7'h65 :
		RG_rl_115_t1 = TR_127 ;
	7'h66 :
		RG_rl_115_t1 = TR_127 ;
	7'h67 :
		RG_rl_115_t1 = TR_127 ;
	7'h68 :
		RG_rl_115_t1 = TR_127 ;
	7'h69 :
		RG_rl_115_t1 = TR_127 ;
	7'h6a :
		RG_rl_115_t1 = TR_127 ;
	7'h6b :
		RG_rl_115_t1 = TR_127 ;
	7'h6c :
		RG_rl_115_t1 = TR_127 ;
	7'h6d :
		RG_rl_115_t1 = TR_127 ;
	7'h6e :
		RG_rl_115_t1 = TR_127 ;
	7'h6f :
		RG_rl_115_t1 = TR_127 ;
	7'h70 :
		RG_rl_115_t1 = TR_127 ;
	7'h71 :
		RG_rl_115_t1 = TR_127 ;
	7'h72 :
		RG_rl_115_t1 = TR_127 ;
	7'h73 :
		RG_rl_115_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h74 :
		RG_rl_115_t1 = TR_127 ;
	7'h75 :
		RG_rl_115_t1 = TR_127 ;
	7'h76 :
		RG_rl_115_t1 = TR_127 ;
	7'h77 :
		RG_rl_115_t1 = TR_127 ;
	7'h78 :
		RG_rl_115_t1 = TR_127 ;
	7'h79 :
		RG_rl_115_t1 = TR_127 ;
	7'h7a :
		RG_rl_115_t1 = TR_127 ;
	7'h7b :
		RG_rl_115_t1 = TR_127 ;
	7'h7c :
		RG_rl_115_t1 = TR_127 ;
	7'h7d :
		RG_rl_115_t1 = TR_127 ;
	7'h7e :
		RG_rl_115_t1 = TR_127 ;
	7'h7f :
		RG_rl_115_t1 = TR_127 ;
	default :
		RG_rl_115_t1 = 9'hx ;
	endcase
always @ ( RG_rl_115_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_56 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_115_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h73 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_115_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_56 )
		| ( { 9{ U_569 } } & RG_rl_115_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_115_en = ( U_570 | RG_rl_115_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_115_en )
		RG_rl_115 <= RG_rl_115_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_128 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_116_t1 = TR_128 ;
	7'h01 :
		RG_rl_116_t1 = TR_128 ;
	7'h02 :
		RG_rl_116_t1 = TR_128 ;
	7'h03 :
		RG_rl_116_t1 = TR_128 ;
	7'h04 :
		RG_rl_116_t1 = TR_128 ;
	7'h05 :
		RG_rl_116_t1 = TR_128 ;
	7'h06 :
		RG_rl_116_t1 = TR_128 ;
	7'h07 :
		RG_rl_116_t1 = TR_128 ;
	7'h08 :
		RG_rl_116_t1 = TR_128 ;
	7'h09 :
		RG_rl_116_t1 = TR_128 ;
	7'h0a :
		RG_rl_116_t1 = TR_128 ;
	7'h0b :
		RG_rl_116_t1 = TR_128 ;
	7'h0c :
		RG_rl_116_t1 = TR_128 ;
	7'h0d :
		RG_rl_116_t1 = TR_128 ;
	7'h0e :
		RG_rl_116_t1 = TR_128 ;
	7'h0f :
		RG_rl_116_t1 = TR_128 ;
	7'h10 :
		RG_rl_116_t1 = TR_128 ;
	7'h11 :
		RG_rl_116_t1 = TR_128 ;
	7'h12 :
		RG_rl_116_t1 = TR_128 ;
	7'h13 :
		RG_rl_116_t1 = TR_128 ;
	7'h14 :
		RG_rl_116_t1 = TR_128 ;
	7'h15 :
		RG_rl_116_t1 = TR_128 ;
	7'h16 :
		RG_rl_116_t1 = TR_128 ;
	7'h17 :
		RG_rl_116_t1 = TR_128 ;
	7'h18 :
		RG_rl_116_t1 = TR_128 ;
	7'h19 :
		RG_rl_116_t1 = TR_128 ;
	7'h1a :
		RG_rl_116_t1 = TR_128 ;
	7'h1b :
		RG_rl_116_t1 = TR_128 ;
	7'h1c :
		RG_rl_116_t1 = TR_128 ;
	7'h1d :
		RG_rl_116_t1 = TR_128 ;
	7'h1e :
		RG_rl_116_t1 = TR_128 ;
	7'h1f :
		RG_rl_116_t1 = TR_128 ;
	7'h20 :
		RG_rl_116_t1 = TR_128 ;
	7'h21 :
		RG_rl_116_t1 = TR_128 ;
	7'h22 :
		RG_rl_116_t1 = TR_128 ;
	7'h23 :
		RG_rl_116_t1 = TR_128 ;
	7'h24 :
		RG_rl_116_t1 = TR_128 ;
	7'h25 :
		RG_rl_116_t1 = TR_128 ;
	7'h26 :
		RG_rl_116_t1 = TR_128 ;
	7'h27 :
		RG_rl_116_t1 = TR_128 ;
	7'h28 :
		RG_rl_116_t1 = TR_128 ;
	7'h29 :
		RG_rl_116_t1 = TR_128 ;
	7'h2a :
		RG_rl_116_t1 = TR_128 ;
	7'h2b :
		RG_rl_116_t1 = TR_128 ;
	7'h2c :
		RG_rl_116_t1 = TR_128 ;
	7'h2d :
		RG_rl_116_t1 = TR_128 ;
	7'h2e :
		RG_rl_116_t1 = TR_128 ;
	7'h2f :
		RG_rl_116_t1 = TR_128 ;
	7'h30 :
		RG_rl_116_t1 = TR_128 ;
	7'h31 :
		RG_rl_116_t1 = TR_128 ;
	7'h32 :
		RG_rl_116_t1 = TR_128 ;
	7'h33 :
		RG_rl_116_t1 = TR_128 ;
	7'h34 :
		RG_rl_116_t1 = TR_128 ;
	7'h35 :
		RG_rl_116_t1 = TR_128 ;
	7'h36 :
		RG_rl_116_t1 = TR_128 ;
	7'h37 :
		RG_rl_116_t1 = TR_128 ;
	7'h38 :
		RG_rl_116_t1 = TR_128 ;
	7'h39 :
		RG_rl_116_t1 = TR_128 ;
	7'h3a :
		RG_rl_116_t1 = TR_128 ;
	7'h3b :
		RG_rl_116_t1 = TR_128 ;
	7'h3c :
		RG_rl_116_t1 = TR_128 ;
	7'h3d :
		RG_rl_116_t1 = TR_128 ;
	7'h3e :
		RG_rl_116_t1 = TR_128 ;
	7'h3f :
		RG_rl_116_t1 = TR_128 ;
	7'h40 :
		RG_rl_116_t1 = TR_128 ;
	7'h41 :
		RG_rl_116_t1 = TR_128 ;
	7'h42 :
		RG_rl_116_t1 = TR_128 ;
	7'h43 :
		RG_rl_116_t1 = TR_128 ;
	7'h44 :
		RG_rl_116_t1 = TR_128 ;
	7'h45 :
		RG_rl_116_t1 = TR_128 ;
	7'h46 :
		RG_rl_116_t1 = TR_128 ;
	7'h47 :
		RG_rl_116_t1 = TR_128 ;
	7'h48 :
		RG_rl_116_t1 = TR_128 ;
	7'h49 :
		RG_rl_116_t1 = TR_128 ;
	7'h4a :
		RG_rl_116_t1 = TR_128 ;
	7'h4b :
		RG_rl_116_t1 = TR_128 ;
	7'h4c :
		RG_rl_116_t1 = TR_128 ;
	7'h4d :
		RG_rl_116_t1 = TR_128 ;
	7'h4e :
		RG_rl_116_t1 = TR_128 ;
	7'h4f :
		RG_rl_116_t1 = TR_128 ;
	7'h50 :
		RG_rl_116_t1 = TR_128 ;
	7'h51 :
		RG_rl_116_t1 = TR_128 ;
	7'h52 :
		RG_rl_116_t1 = TR_128 ;
	7'h53 :
		RG_rl_116_t1 = TR_128 ;
	7'h54 :
		RG_rl_116_t1 = TR_128 ;
	7'h55 :
		RG_rl_116_t1 = TR_128 ;
	7'h56 :
		RG_rl_116_t1 = TR_128 ;
	7'h57 :
		RG_rl_116_t1 = TR_128 ;
	7'h58 :
		RG_rl_116_t1 = TR_128 ;
	7'h59 :
		RG_rl_116_t1 = TR_128 ;
	7'h5a :
		RG_rl_116_t1 = TR_128 ;
	7'h5b :
		RG_rl_116_t1 = TR_128 ;
	7'h5c :
		RG_rl_116_t1 = TR_128 ;
	7'h5d :
		RG_rl_116_t1 = TR_128 ;
	7'h5e :
		RG_rl_116_t1 = TR_128 ;
	7'h5f :
		RG_rl_116_t1 = TR_128 ;
	7'h60 :
		RG_rl_116_t1 = TR_128 ;
	7'h61 :
		RG_rl_116_t1 = TR_128 ;
	7'h62 :
		RG_rl_116_t1 = TR_128 ;
	7'h63 :
		RG_rl_116_t1 = TR_128 ;
	7'h64 :
		RG_rl_116_t1 = TR_128 ;
	7'h65 :
		RG_rl_116_t1 = TR_128 ;
	7'h66 :
		RG_rl_116_t1 = TR_128 ;
	7'h67 :
		RG_rl_116_t1 = TR_128 ;
	7'h68 :
		RG_rl_116_t1 = TR_128 ;
	7'h69 :
		RG_rl_116_t1 = TR_128 ;
	7'h6a :
		RG_rl_116_t1 = TR_128 ;
	7'h6b :
		RG_rl_116_t1 = TR_128 ;
	7'h6c :
		RG_rl_116_t1 = TR_128 ;
	7'h6d :
		RG_rl_116_t1 = TR_128 ;
	7'h6e :
		RG_rl_116_t1 = TR_128 ;
	7'h6f :
		RG_rl_116_t1 = TR_128 ;
	7'h70 :
		RG_rl_116_t1 = TR_128 ;
	7'h71 :
		RG_rl_116_t1 = TR_128 ;
	7'h72 :
		RG_rl_116_t1 = TR_128 ;
	7'h73 :
		RG_rl_116_t1 = TR_128 ;
	7'h74 :
		RG_rl_116_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h75 :
		RG_rl_116_t1 = TR_128 ;
	7'h76 :
		RG_rl_116_t1 = TR_128 ;
	7'h77 :
		RG_rl_116_t1 = TR_128 ;
	7'h78 :
		RG_rl_116_t1 = TR_128 ;
	7'h79 :
		RG_rl_116_t1 = TR_128 ;
	7'h7a :
		RG_rl_116_t1 = TR_128 ;
	7'h7b :
		RG_rl_116_t1 = TR_128 ;
	7'h7c :
		RG_rl_116_t1 = TR_128 ;
	7'h7d :
		RG_rl_116_t1 = TR_128 ;
	7'h7e :
		RG_rl_116_t1 = TR_128 ;
	7'h7f :
		RG_rl_116_t1 = TR_128 ;
	default :
		RG_rl_116_t1 = 9'hx ;
	endcase
always @ ( RG_rl_116_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_242 or M_318 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_116_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h74 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_116_t = ( ( { 9{ M_318 } } & RG_rl_242 )
		| ( { 9{ U_569 } } & RG_rl_116_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_116_en = ( M_318 | RG_rl_116_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_116_en )
		RG_rl_116 <= RG_rl_116_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_129 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_117_t1 = TR_129 ;
	7'h01 :
		RG_rl_117_t1 = TR_129 ;
	7'h02 :
		RG_rl_117_t1 = TR_129 ;
	7'h03 :
		RG_rl_117_t1 = TR_129 ;
	7'h04 :
		RG_rl_117_t1 = TR_129 ;
	7'h05 :
		RG_rl_117_t1 = TR_129 ;
	7'h06 :
		RG_rl_117_t1 = TR_129 ;
	7'h07 :
		RG_rl_117_t1 = TR_129 ;
	7'h08 :
		RG_rl_117_t1 = TR_129 ;
	7'h09 :
		RG_rl_117_t1 = TR_129 ;
	7'h0a :
		RG_rl_117_t1 = TR_129 ;
	7'h0b :
		RG_rl_117_t1 = TR_129 ;
	7'h0c :
		RG_rl_117_t1 = TR_129 ;
	7'h0d :
		RG_rl_117_t1 = TR_129 ;
	7'h0e :
		RG_rl_117_t1 = TR_129 ;
	7'h0f :
		RG_rl_117_t1 = TR_129 ;
	7'h10 :
		RG_rl_117_t1 = TR_129 ;
	7'h11 :
		RG_rl_117_t1 = TR_129 ;
	7'h12 :
		RG_rl_117_t1 = TR_129 ;
	7'h13 :
		RG_rl_117_t1 = TR_129 ;
	7'h14 :
		RG_rl_117_t1 = TR_129 ;
	7'h15 :
		RG_rl_117_t1 = TR_129 ;
	7'h16 :
		RG_rl_117_t1 = TR_129 ;
	7'h17 :
		RG_rl_117_t1 = TR_129 ;
	7'h18 :
		RG_rl_117_t1 = TR_129 ;
	7'h19 :
		RG_rl_117_t1 = TR_129 ;
	7'h1a :
		RG_rl_117_t1 = TR_129 ;
	7'h1b :
		RG_rl_117_t1 = TR_129 ;
	7'h1c :
		RG_rl_117_t1 = TR_129 ;
	7'h1d :
		RG_rl_117_t1 = TR_129 ;
	7'h1e :
		RG_rl_117_t1 = TR_129 ;
	7'h1f :
		RG_rl_117_t1 = TR_129 ;
	7'h20 :
		RG_rl_117_t1 = TR_129 ;
	7'h21 :
		RG_rl_117_t1 = TR_129 ;
	7'h22 :
		RG_rl_117_t1 = TR_129 ;
	7'h23 :
		RG_rl_117_t1 = TR_129 ;
	7'h24 :
		RG_rl_117_t1 = TR_129 ;
	7'h25 :
		RG_rl_117_t1 = TR_129 ;
	7'h26 :
		RG_rl_117_t1 = TR_129 ;
	7'h27 :
		RG_rl_117_t1 = TR_129 ;
	7'h28 :
		RG_rl_117_t1 = TR_129 ;
	7'h29 :
		RG_rl_117_t1 = TR_129 ;
	7'h2a :
		RG_rl_117_t1 = TR_129 ;
	7'h2b :
		RG_rl_117_t1 = TR_129 ;
	7'h2c :
		RG_rl_117_t1 = TR_129 ;
	7'h2d :
		RG_rl_117_t1 = TR_129 ;
	7'h2e :
		RG_rl_117_t1 = TR_129 ;
	7'h2f :
		RG_rl_117_t1 = TR_129 ;
	7'h30 :
		RG_rl_117_t1 = TR_129 ;
	7'h31 :
		RG_rl_117_t1 = TR_129 ;
	7'h32 :
		RG_rl_117_t1 = TR_129 ;
	7'h33 :
		RG_rl_117_t1 = TR_129 ;
	7'h34 :
		RG_rl_117_t1 = TR_129 ;
	7'h35 :
		RG_rl_117_t1 = TR_129 ;
	7'h36 :
		RG_rl_117_t1 = TR_129 ;
	7'h37 :
		RG_rl_117_t1 = TR_129 ;
	7'h38 :
		RG_rl_117_t1 = TR_129 ;
	7'h39 :
		RG_rl_117_t1 = TR_129 ;
	7'h3a :
		RG_rl_117_t1 = TR_129 ;
	7'h3b :
		RG_rl_117_t1 = TR_129 ;
	7'h3c :
		RG_rl_117_t1 = TR_129 ;
	7'h3d :
		RG_rl_117_t1 = TR_129 ;
	7'h3e :
		RG_rl_117_t1 = TR_129 ;
	7'h3f :
		RG_rl_117_t1 = TR_129 ;
	7'h40 :
		RG_rl_117_t1 = TR_129 ;
	7'h41 :
		RG_rl_117_t1 = TR_129 ;
	7'h42 :
		RG_rl_117_t1 = TR_129 ;
	7'h43 :
		RG_rl_117_t1 = TR_129 ;
	7'h44 :
		RG_rl_117_t1 = TR_129 ;
	7'h45 :
		RG_rl_117_t1 = TR_129 ;
	7'h46 :
		RG_rl_117_t1 = TR_129 ;
	7'h47 :
		RG_rl_117_t1 = TR_129 ;
	7'h48 :
		RG_rl_117_t1 = TR_129 ;
	7'h49 :
		RG_rl_117_t1 = TR_129 ;
	7'h4a :
		RG_rl_117_t1 = TR_129 ;
	7'h4b :
		RG_rl_117_t1 = TR_129 ;
	7'h4c :
		RG_rl_117_t1 = TR_129 ;
	7'h4d :
		RG_rl_117_t1 = TR_129 ;
	7'h4e :
		RG_rl_117_t1 = TR_129 ;
	7'h4f :
		RG_rl_117_t1 = TR_129 ;
	7'h50 :
		RG_rl_117_t1 = TR_129 ;
	7'h51 :
		RG_rl_117_t1 = TR_129 ;
	7'h52 :
		RG_rl_117_t1 = TR_129 ;
	7'h53 :
		RG_rl_117_t1 = TR_129 ;
	7'h54 :
		RG_rl_117_t1 = TR_129 ;
	7'h55 :
		RG_rl_117_t1 = TR_129 ;
	7'h56 :
		RG_rl_117_t1 = TR_129 ;
	7'h57 :
		RG_rl_117_t1 = TR_129 ;
	7'h58 :
		RG_rl_117_t1 = TR_129 ;
	7'h59 :
		RG_rl_117_t1 = TR_129 ;
	7'h5a :
		RG_rl_117_t1 = TR_129 ;
	7'h5b :
		RG_rl_117_t1 = TR_129 ;
	7'h5c :
		RG_rl_117_t1 = TR_129 ;
	7'h5d :
		RG_rl_117_t1 = TR_129 ;
	7'h5e :
		RG_rl_117_t1 = TR_129 ;
	7'h5f :
		RG_rl_117_t1 = TR_129 ;
	7'h60 :
		RG_rl_117_t1 = TR_129 ;
	7'h61 :
		RG_rl_117_t1 = TR_129 ;
	7'h62 :
		RG_rl_117_t1 = TR_129 ;
	7'h63 :
		RG_rl_117_t1 = TR_129 ;
	7'h64 :
		RG_rl_117_t1 = TR_129 ;
	7'h65 :
		RG_rl_117_t1 = TR_129 ;
	7'h66 :
		RG_rl_117_t1 = TR_129 ;
	7'h67 :
		RG_rl_117_t1 = TR_129 ;
	7'h68 :
		RG_rl_117_t1 = TR_129 ;
	7'h69 :
		RG_rl_117_t1 = TR_129 ;
	7'h6a :
		RG_rl_117_t1 = TR_129 ;
	7'h6b :
		RG_rl_117_t1 = TR_129 ;
	7'h6c :
		RG_rl_117_t1 = TR_129 ;
	7'h6d :
		RG_rl_117_t1 = TR_129 ;
	7'h6e :
		RG_rl_117_t1 = TR_129 ;
	7'h6f :
		RG_rl_117_t1 = TR_129 ;
	7'h70 :
		RG_rl_117_t1 = TR_129 ;
	7'h71 :
		RG_rl_117_t1 = TR_129 ;
	7'h72 :
		RG_rl_117_t1 = TR_129 ;
	7'h73 :
		RG_rl_117_t1 = TR_129 ;
	7'h74 :
		RG_rl_117_t1 = TR_129 ;
	7'h75 :
		RG_rl_117_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h76 :
		RG_rl_117_t1 = TR_129 ;
	7'h77 :
		RG_rl_117_t1 = TR_129 ;
	7'h78 :
		RG_rl_117_t1 = TR_129 ;
	7'h79 :
		RG_rl_117_t1 = TR_129 ;
	7'h7a :
		RG_rl_117_t1 = TR_129 ;
	7'h7b :
		RG_rl_117_t1 = TR_129 ;
	7'h7c :
		RG_rl_117_t1 = TR_129 ;
	7'h7d :
		RG_rl_117_t1 = TR_129 ;
	7'h7e :
		RG_rl_117_t1 = TR_129 ;
	7'h7f :
		RG_rl_117_t1 = TR_129 ;
	default :
		RG_rl_117_t1 = 9'hx ;
	endcase
always @ ( RG_rl_117_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_57 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_117_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h75 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_117_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_57 )
		| ( { 9{ U_569 } } & RG_rl_117_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_117_en = ( U_570 | RG_rl_117_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_117_en )
		RG_rl_117 <= RG_rl_117_t ;	// line#=../rle.cpp:79,80,83,84,85
assign	M_318 = ( ST1_01d | U_570 ) ;	// line#=../rle.cpp:83,84,85
always @ ( TR_130 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_118_t1 = TR_130 ;
	7'h01 :
		RG_rl_118_t1 = TR_130 ;
	7'h02 :
		RG_rl_118_t1 = TR_130 ;
	7'h03 :
		RG_rl_118_t1 = TR_130 ;
	7'h04 :
		RG_rl_118_t1 = TR_130 ;
	7'h05 :
		RG_rl_118_t1 = TR_130 ;
	7'h06 :
		RG_rl_118_t1 = TR_130 ;
	7'h07 :
		RG_rl_118_t1 = TR_130 ;
	7'h08 :
		RG_rl_118_t1 = TR_130 ;
	7'h09 :
		RG_rl_118_t1 = TR_130 ;
	7'h0a :
		RG_rl_118_t1 = TR_130 ;
	7'h0b :
		RG_rl_118_t1 = TR_130 ;
	7'h0c :
		RG_rl_118_t1 = TR_130 ;
	7'h0d :
		RG_rl_118_t1 = TR_130 ;
	7'h0e :
		RG_rl_118_t1 = TR_130 ;
	7'h0f :
		RG_rl_118_t1 = TR_130 ;
	7'h10 :
		RG_rl_118_t1 = TR_130 ;
	7'h11 :
		RG_rl_118_t1 = TR_130 ;
	7'h12 :
		RG_rl_118_t1 = TR_130 ;
	7'h13 :
		RG_rl_118_t1 = TR_130 ;
	7'h14 :
		RG_rl_118_t1 = TR_130 ;
	7'h15 :
		RG_rl_118_t1 = TR_130 ;
	7'h16 :
		RG_rl_118_t1 = TR_130 ;
	7'h17 :
		RG_rl_118_t1 = TR_130 ;
	7'h18 :
		RG_rl_118_t1 = TR_130 ;
	7'h19 :
		RG_rl_118_t1 = TR_130 ;
	7'h1a :
		RG_rl_118_t1 = TR_130 ;
	7'h1b :
		RG_rl_118_t1 = TR_130 ;
	7'h1c :
		RG_rl_118_t1 = TR_130 ;
	7'h1d :
		RG_rl_118_t1 = TR_130 ;
	7'h1e :
		RG_rl_118_t1 = TR_130 ;
	7'h1f :
		RG_rl_118_t1 = TR_130 ;
	7'h20 :
		RG_rl_118_t1 = TR_130 ;
	7'h21 :
		RG_rl_118_t1 = TR_130 ;
	7'h22 :
		RG_rl_118_t1 = TR_130 ;
	7'h23 :
		RG_rl_118_t1 = TR_130 ;
	7'h24 :
		RG_rl_118_t1 = TR_130 ;
	7'h25 :
		RG_rl_118_t1 = TR_130 ;
	7'h26 :
		RG_rl_118_t1 = TR_130 ;
	7'h27 :
		RG_rl_118_t1 = TR_130 ;
	7'h28 :
		RG_rl_118_t1 = TR_130 ;
	7'h29 :
		RG_rl_118_t1 = TR_130 ;
	7'h2a :
		RG_rl_118_t1 = TR_130 ;
	7'h2b :
		RG_rl_118_t1 = TR_130 ;
	7'h2c :
		RG_rl_118_t1 = TR_130 ;
	7'h2d :
		RG_rl_118_t1 = TR_130 ;
	7'h2e :
		RG_rl_118_t1 = TR_130 ;
	7'h2f :
		RG_rl_118_t1 = TR_130 ;
	7'h30 :
		RG_rl_118_t1 = TR_130 ;
	7'h31 :
		RG_rl_118_t1 = TR_130 ;
	7'h32 :
		RG_rl_118_t1 = TR_130 ;
	7'h33 :
		RG_rl_118_t1 = TR_130 ;
	7'h34 :
		RG_rl_118_t1 = TR_130 ;
	7'h35 :
		RG_rl_118_t1 = TR_130 ;
	7'h36 :
		RG_rl_118_t1 = TR_130 ;
	7'h37 :
		RG_rl_118_t1 = TR_130 ;
	7'h38 :
		RG_rl_118_t1 = TR_130 ;
	7'h39 :
		RG_rl_118_t1 = TR_130 ;
	7'h3a :
		RG_rl_118_t1 = TR_130 ;
	7'h3b :
		RG_rl_118_t1 = TR_130 ;
	7'h3c :
		RG_rl_118_t1 = TR_130 ;
	7'h3d :
		RG_rl_118_t1 = TR_130 ;
	7'h3e :
		RG_rl_118_t1 = TR_130 ;
	7'h3f :
		RG_rl_118_t1 = TR_130 ;
	7'h40 :
		RG_rl_118_t1 = TR_130 ;
	7'h41 :
		RG_rl_118_t1 = TR_130 ;
	7'h42 :
		RG_rl_118_t1 = TR_130 ;
	7'h43 :
		RG_rl_118_t1 = TR_130 ;
	7'h44 :
		RG_rl_118_t1 = TR_130 ;
	7'h45 :
		RG_rl_118_t1 = TR_130 ;
	7'h46 :
		RG_rl_118_t1 = TR_130 ;
	7'h47 :
		RG_rl_118_t1 = TR_130 ;
	7'h48 :
		RG_rl_118_t1 = TR_130 ;
	7'h49 :
		RG_rl_118_t1 = TR_130 ;
	7'h4a :
		RG_rl_118_t1 = TR_130 ;
	7'h4b :
		RG_rl_118_t1 = TR_130 ;
	7'h4c :
		RG_rl_118_t1 = TR_130 ;
	7'h4d :
		RG_rl_118_t1 = TR_130 ;
	7'h4e :
		RG_rl_118_t1 = TR_130 ;
	7'h4f :
		RG_rl_118_t1 = TR_130 ;
	7'h50 :
		RG_rl_118_t1 = TR_130 ;
	7'h51 :
		RG_rl_118_t1 = TR_130 ;
	7'h52 :
		RG_rl_118_t1 = TR_130 ;
	7'h53 :
		RG_rl_118_t1 = TR_130 ;
	7'h54 :
		RG_rl_118_t1 = TR_130 ;
	7'h55 :
		RG_rl_118_t1 = TR_130 ;
	7'h56 :
		RG_rl_118_t1 = TR_130 ;
	7'h57 :
		RG_rl_118_t1 = TR_130 ;
	7'h58 :
		RG_rl_118_t1 = TR_130 ;
	7'h59 :
		RG_rl_118_t1 = TR_130 ;
	7'h5a :
		RG_rl_118_t1 = TR_130 ;
	7'h5b :
		RG_rl_118_t1 = TR_130 ;
	7'h5c :
		RG_rl_118_t1 = TR_130 ;
	7'h5d :
		RG_rl_118_t1 = TR_130 ;
	7'h5e :
		RG_rl_118_t1 = TR_130 ;
	7'h5f :
		RG_rl_118_t1 = TR_130 ;
	7'h60 :
		RG_rl_118_t1 = TR_130 ;
	7'h61 :
		RG_rl_118_t1 = TR_130 ;
	7'h62 :
		RG_rl_118_t1 = TR_130 ;
	7'h63 :
		RG_rl_118_t1 = TR_130 ;
	7'h64 :
		RG_rl_118_t1 = TR_130 ;
	7'h65 :
		RG_rl_118_t1 = TR_130 ;
	7'h66 :
		RG_rl_118_t1 = TR_130 ;
	7'h67 :
		RG_rl_118_t1 = TR_130 ;
	7'h68 :
		RG_rl_118_t1 = TR_130 ;
	7'h69 :
		RG_rl_118_t1 = TR_130 ;
	7'h6a :
		RG_rl_118_t1 = TR_130 ;
	7'h6b :
		RG_rl_118_t1 = TR_130 ;
	7'h6c :
		RG_rl_118_t1 = TR_130 ;
	7'h6d :
		RG_rl_118_t1 = TR_130 ;
	7'h6e :
		RG_rl_118_t1 = TR_130 ;
	7'h6f :
		RG_rl_118_t1 = TR_130 ;
	7'h70 :
		RG_rl_118_t1 = TR_130 ;
	7'h71 :
		RG_rl_118_t1 = TR_130 ;
	7'h72 :
		RG_rl_118_t1 = TR_130 ;
	7'h73 :
		RG_rl_118_t1 = TR_130 ;
	7'h74 :
		RG_rl_118_t1 = TR_130 ;
	7'h75 :
		RG_rl_118_t1 = TR_130 ;
	7'h76 :
		RG_rl_118_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h77 :
		RG_rl_118_t1 = TR_130 ;
	7'h78 :
		RG_rl_118_t1 = TR_130 ;
	7'h79 :
		RG_rl_118_t1 = TR_130 ;
	7'h7a :
		RG_rl_118_t1 = TR_130 ;
	7'h7b :
		RG_rl_118_t1 = TR_130 ;
	7'h7c :
		RG_rl_118_t1 = TR_130 ;
	7'h7d :
		RG_rl_118_t1 = TR_130 ;
	7'h7e :
		RG_rl_118_t1 = TR_130 ;
	7'h7f :
		RG_rl_118_t1 = TR_130 ;
	default :
		RG_rl_118_t1 = 9'hx ;
	endcase
always @ ( RG_rl_118_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_243 or M_318 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_118_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h76 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_118_t = ( ( { 9{ M_318 } } & RG_rl_243 )
		| ( { 9{ U_569 } } & RG_rl_118_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_118_en = ( M_318 | RG_rl_118_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_118_en )
		RG_rl_118 <= RG_rl_118_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_131 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_119_t1 = TR_131 ;
	7'h01 :
		RG_rl_119_t1 = TR_131 ;
	7'h02 :
		RG_rl_119_t1 = TR_131 ;
	7'h03 :
		RG_rl_119_t1 = TR_131 ;
	7'h04 :
		RG_rl_119_t1 = TR_131 ;
	7'h05 :
		RG_rl_119_t1 = TR_131 ;
	7'h06 :
		RG_rl_119_t1 = TR_131 ;
	7'h07 :
		RG_rl_119_t1 = TR_131 ;
	7'h08 :
		RG_rl_119_t1 = TR_131 ;
	7'h09 :
		RG_rl_119_t1 = TR_131 ;
	7'h0a :
		RG_rl_119_t1 = TR_131 ;
	7'h0b :
		RG_rl_119_t1 = TR_131 ;
	7'h0c :
		RG_rl_119_t1 = TR_131 ;
	7'h0d :
		RG_rl_119_t1 = TR_131 ;
	7'h0e :
		RG_rl_119_t1 = TR_131 ;
	7'h0f :
		RG_rl_119_t1 = TR_131 ;
	7'h10 :
		RG_rl_119_t1 = TR_131 ;
	7'h11 :
		RG_rl_119_t1 = TR_131 ;
	7'h12 :
		RG_rl_119_t1 = TR_131 ;
	7'h13 :
		RG_rl_119_t1 = TR_131 ;
	7'h14 :
		RG_rl_119_t1 = TR_131 ;
	7'h15 :
		RG_rl_119_t1 = TR_131 ;
	7'h16 :
		RG_rl_119_t1 = TR_131 ;
	7'h17 :
		RG_rl_119_t1 = TR_131 ;
	7'h18 :
		RG_rl_119_t1 = TR_131 ;
	7'h19 :
		RG_rl_119_t1 = TR_131 ;
	7'h1a :
		RG_rl_119_t1 = TR_131 ;
	7'h1b :
		RG_rl_119_t1 = TR_131 ;
	7'h1c :
		RG_rl_119_t1 = TR_131 ;
	7'h1d :
		RG_rl_119_t1 = TR_131 ;
	7'h1e :
		RG_rl_119_t1 = TR_131 ;
	7'h1f :
		RG_rl_119_t1 = TR_131 ;
	7'h20 :
		RG_rl_119_t1 = TR_131 ;
	7'h21 :
		RG_rl_119_t1 = TR_131 ;
	7'h22 :
		RG_rl_119_t1 = TR_131 ;
	7'h23 :
		RG_rl_119_t1 = TR_131 ;
	7'h24 :
		RG_rl_119_t1 = TR_131 ;
	7'h25 :
		RG_rl_119_t1 = TR_131 ;
	7'h26 :
		RG_rl_119_t1 = TR_131 ;
	7'h27 :
		RG_rl_119_t1 = TR_131 ;
	7'h28 :
		RG_rl_119_t1 = TR_131 ;
	7'h29 :
		RG_rl_119_t1 = TR_131 ;
	7'h2a :
		RG_rl_119_t1 = TR_131 ;
	7'h2b :
		RG_rl_119_t1 = TR_131 ;
	7'h2c :
		RG_rl_119_t1 = TR_131 ;
	7'h2d :
		RG_rl_119_t1 = TR_131 ;
	7'h2e :
		RG_rl_119_t1 = TR_131 ;
	7'h2f :
		RG_rl_119_t1 = TR_131 ;
	7'h30 :
		RG_rl_119_t1 = TR_131 ;
	7'h31 :
		RG_rl_119_t1 = TR_131 ;
	7'h32 :
		RG_rl_119_t1 = TR_131 ;
	7'h33 :
		RG_rl_119_t1 = TR_131 ;
	7'h34 :
		RG_rl_119_t1 = TR_131 ;
	7'h35 :
		RG_rl_119_t1 = TR_131 ;
	7'h36 :
		RG_rl_119_t1 = TR_131 ;
	7'h37 :
		RG_rl_119_t1 = TR_131 ;
	7'h38 :
		RG_rl_119_t1 = TR_131 ;
	7'h39 :
		RG_rl_119_t1 = TR_131 ;
	7'h3a :
		RG_rl_119_t1 = TR_131 ;
	7'h3b :
		RG_rl_119_t1 = TR_131 ;
	7'h3c :
		RG_rl_119_t1 = TR_131 ;
	7'h3d :
		RG_rl_119_t1 = TR_131 ;
	7'h3e :
		RG_rl_119_t1 = TR_131 ;
	7'h3f :
		RG_rl_119_t1 = TR_131 ;
	7'h40 :
		RG_rl_119_t1 = TR_131 ;
	7'h41 :
		RG_rl_119_t1 = TR_131 ;
	7'h42 :
		RG_rl_119_t1 = TR_131 ;
	7'h43 :
		RG_rl_119_t1 = TR_131 ;
	7'h44 :
		RG_rl_119_t1 = TR_131 ;
	7'h45 :
		RG_rl_119_t1 = TR_131 ;
	7'h46 :
		RG_rl_119_t1 = TR_131 ;
	7'h47 :
		RG_rl_119_t1 = TR_131 ;
	7'h48 :
		RG_rl_119_t1 = TR_131 ;
	7'h49 :
		RG_rl_119_t1 = TR_131 ;
	7'h4a :
		RG_rl_119_t1 = TR_131 ;
	7'h4b :
		RG_rl_119_t1 = TR_131 ;
	7'h4c :
		RG_rl_119_t1 = TR_131 ;
	7'h4d :
		RG_rl_119_t1 = TR_131 ;
	7'h4e :
		RG_rl_119_t1 = TR_131 ;
	7'h4f :
		RG_rl_119_t1 = TR_131 ;
	7'h50 :
		RG_rl_119_t1 = TR_131 ;
	7'h51 :
		RG_rl_119_t1 = TR_131 ;
	7'h52 :
		RG_rl_119_t1 = TR_131 ;
	7'h53 :
		RG_rl_119_t1 = TR_131 ;
	7'h54 :
		RG_rl_119_t1 = TR_131 ;
	7'h55 :
		RG_rl_119_t1 = TR_131 ;
	7'h56 :
		RG_rl_119_t1 = TR_131 ;
	7'h57 :
		RG_rl_119_t1 = TR_131 ;
	7'h58 :
		RG_rl_119_t1 = TR_131 ;
	7'h59 :
		RG_rl_119_t1 = TR_131 ;
	7'h5a :
		RG_rl_119_t1 = TR_131 ;
	7'h5b :
		RG_rl_119_t1 = TR_131 ;
	7'h5c :
		RG_rl_119_t1 = TR_131 ;
	7'h5d :
		RG_rl_119_t1 = TR_131 ;
	7'h5e :
		RG_rl_119_t1 = TR_131 ;
	7'h5f :
		RG_rl_119_t1 = TR_131 ;
	7'h60 :
		RG_rl_119_t1 = TR_131 ;
	7'h61 :
		RG_rl_119_t1 = TR_131 ;
	7'h62 :
		RG_rl_119_t1 = TR_131 ;
	7'h63 :
		RG_rl_119_t1 = TR_131 ;
	7'h64 :
		RG_rl_119_t1 = TR_131 ;
	7'h65 :
		RG_rl_119_t1 = TR_131 ;
	7'h66 :
		RG_rl_119_t1 = TR_131 ;
	7'h67 :
		RG_rl_119_t1 = TR_131 ;
	7'h68 :
		RG_rl_119_t1 = TR_131 ;
	7'h69 :
		RG_rl_119_t1 = TR_131 ;
	7'h6a :
		RG_rl_119_t1 = TR_131 ;
	7'h6b :
		RG_rl_119_t1 = TR_131 ;
	7'h6c :
		RG_rl_119_t1 = TR_131 ;
	7'h6d :
		RG_rl_119_t1 = TR_131 ;
	7'h6e :
		RG_rl_119_t1 = TR_131 ;
	7'h6f :
		RG_rl_119_t1 = TR_131 ;
	7'h70 :
		RG_rl_119_t1 = TR_131 ;
	7'h71 :
		RG_rl_119_t1 = TR_131 ;
	7'h72 :
		RG_rl_119_t1 = TR_131 ;
	7'h73 :
		RG_rl_119_t1 = TR_131 ;
	7'h74 :
		RG_rl_119_t1 = TR_131 ;
	7'h75 :
		RG_rl_119_t1 = TR_131 ;
	7'h76 :
		RG_rl_119_t1 = TR_131 ;
	7'h77 :
		RG_rl_119_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h78 :
		RG_rl_119_t1 = TR_131 ;
	7'h79 :
		RG_rl_119_t1 = TR_131 ;
	7'h7a :
		RG_rl_119_t1 = TR_131 ;
	7'h7b :
		RG_rl_119_t1 = TR_131 ;
	7'h7c :
		RG_rl_119_t1 = TR_131 ;
	7'h7d :
		RG_rl_119_t1 = TR_131 ;
	7'h7e :
		RG_rl_119_t1 = TR_131 ;
	7'h7f :
		RG_rl_119_t1 = TR_131 ;
	default :
		RG_rl_119_t1 = 9'hx ;
	endcase
always @ ( RG_rl_119_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_58 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_119_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h77 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_119_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_58 )
		| ( { 9{ U_569 } } & RG_rl_119_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_119_en = ( U_570 | RG_rl_119_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_119_en )
		RG_rl_119 <= RG_rl_119_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_132 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_120_t1 = TR_132 ;
	7'h01 :
		RG_rl_120_t1 = TR_132 ;
	7'h02 :
		RG_rl_120_t1 = TR_132 ;
	7'h03 :
		RG_rl_120_t1 = TR_132 ;
	7'h04 :
		RG_rl_120_t1 = TR_132 ;
	7'h05 :
		RG_rl_120_t1 = TR_132 ;
	7'h06 :
		RG_rl_120_t1 = TR_132 ;
	7'h07 :
		RG_rl_120_t1 = TR_132 ;
	7'h08 :
		RG_rl_120_t1 = TR_132 ;
	7'h09 :
		RG_rl_120_t1 = TR_132 ;
	7'h0a :
		RG_rl_120_t1 = TR_132 ;
	7'h0b :
		RG_rl_120_t1 = TR_132 ;
	7'h0c :
		RG_rl_120_t1 = TR_132 ;
	7'h0d :
		RG_rl_120_t1 = TR_132 ;
	7'h0e :
		RG_rl_120_t1 = TR_132 ;
	7'h0f :
		RG_rl_120_t1 = TR_132 ;
	7'h10 :
		RG_rl_120_t1 = TR_132 ;
	7'h11 :
		RG_rl_120_t1 = TR_132 ;
	7'h12 :
		RG_rl_120_t1 = TR_132 ;
	7'h13 :
		RG_rl_120_t1 = TR_132 ;
	7'h14 :
		RG_rl_120_t1 = TR_132 ;
	7'h15 :
		RG_rl_120_t1 = TR_132 ;
	7'h16 :
		RG_rl_120_t1 = TR_132 ;
	7'h17 :
		RG_rl_120_t1 = TR_132 ;
	7'h18 :
		RG_rl_120_t1 = TR_132 ;
	7'h19 :
		RG_rl_120_t1 = TR_132 ;
	7'h1a :
		RG_rl_120_t1 = TR_132 ;
	7'h1b :
		RG_rl_120_t1 = TR_132 ;
	7'h1c :
		RG_rl_120_t1 = TR_132 ;
	7'h1d :
		RG_rl_120_t1 = TR_132 ;
	7'h1e :
		RG_rl_120_t1 = TR_132 ;
	7'h1f :
		RG_rl_120_t1 = TR_132 ;
	7'h20 :
		RG_rl_120_t1 = TR_132 ;
	7'h21 :
		RG_rl_120_t1 = TR_132 ;
	7'h22 :
		RG_rl_120_t1 = TR_132 ;
	7'h23 :
		RG_rl_120_t1 = TR_132 ;
	7'h24 :
		RG_rl_120_t1 = TR_132 ;
	7'h25 :
		RG_rl_120_t1 = TR_132 ;
	7'h26 :
		RG_rl_120_t1 = TR_132 ;
	7'h27 :
		RG_rl_120_t1 = TR_132 ;
	7'h28 :
		RG_rl_120_t1 = TR_132 ;
	7'h29 :
		RG_rl_120_t1 = TR_132 ;
	7'h2a :
		RG_rl_120_t1 = TR_132 ;
	7'h2b :
		RG_rl_120_t1 = TR_132 ;
	7'h2c :
		RG_rl_120_t1 = TR_132 ;
	7'h2d :
		RG_rl_120_t1 = TR_132 ;
	7'h2e :
		RG_rl_120_t1 = TR_132 ;
	7'h2f :
		RG_rl_120_t1 = TR_132 ;
	7'h30 :
		RG_rl_120_t1 = TR_132 ;
	7'h31 :
		RG_rl_120_t1 = TR_132 ;
	7'h32 :
		RG_rl_120_t1 = TR_132 ;
	7'h33 :
		RG_rl_120_t1 = TR_132 ;
	7'h34 :
		RG_rl_120_t1 = TR_132 ;
	7'h35 :
		RG_rl_120_t1 = TR_132 ;
	7'h36 :
		RG_rl_120_t1 = TR_132 ;
	7'h37 :
		RG_rl_120_t1 = TR_132 ;
	7'h38 :
		RG_rl_120_t1 = TR_132 ;
	7'h39 :
		RG_rl_120_t1 = TR_132 ;
	7'h3a :
		RG_rl_120_t1 = TR_132 ;
	7'h3b :
		RG_rl_120_t1 = TR_132 ;
	7'h3c :
		RG_rl_120_t1 = TR_132 ;
	7'h3d :
		RG_rl_120_t1 = TR_132 ;
	7'h3e :
		RG_rl_120_t1 = TR_132 ;
	7'h3f :
		RG_rl_120_t1 = TR_132 ;
	7'h40 :
		RG_rl_120_t1 = TR_132 ;
	7'h41 :
		RG_rl_120_t1 = TR_132 ;
	7'h42 :
		RG_rl_120_t1 = TR_132 ;
	7'h43 :
		RG_rl_120_t1 = TR_132 ;
	7'h44 :
		RG_rl_120_t1 = TR_132 ;
	7'h45 :
		RG_rl_120_t1 = TR_132 ;
	7'h46 :
		RG_rl_120_t1 = TR_132 ;
	7'h47 :
		RG_rl_120_t1 = TR_132 ;
	7'h48 :
		RG_rl_120_t1 = TR_132 ;
	7'h49 :
		RG_rl_120_t1 = TR_132 ;
	7'h4a :
		RG_rl_120_t1 = TR_132 ;
	7'h4b :
		RG_rl_120_t1 = TR_132 ;
	7'h4c :
		RG_rl_120_t1 = TR_132 ;
	7'h4d :
		RG_rl_120_t1 = TR_132 ;
	7'h4e :
		RG_rl_120_t1 = TR_132 ;
	7'h4f :
		RG_rl_120_t1 = TR_132 ;
	7'h50 :
		RG_rl_120_t1 = TR_132 ;
	7'h51 :
		RG_rl_120_t1 = TR_132 ;
	7'h52 :
		RG_rl_120_t1 = TR_132 ;
	7'h53 :
		RG_rl_120_t1 = TR_132 ;
	7'h54 :
		RG_rl_120_t1 = TR_132 ;
	7'h55 :
		RG_rl_120_t1 = TR_132 ;
	7'h56 :
		RG_rl_120_t1 = TR_132 ;
	7'h57 :
		RG_rl_120_t1 = TR_132 ;
	7'h58 :
		RG_rl_120_t1 = TR_132 ;
	7'h59 :
		RG_rl_120_t1 = TR_132 ;
	7'h5a :
		RG_rl_120_t1 = TR_132 ;
	7'h5b :
		RG_rl_120_t1 = TR_132 ;
	7'h5c :
		RG_rl_120_t1 = TR_132 ;
	7'h5d :
		RG_rl_120_t1 = TR_132 ;
	7'h5e :
		RG_rl_120_t1 = TR_132 ;
	7'h5f :
		RG_rl_120_t1 = TR_132 ;
	7'h60 :
		RG_rl_120_t1 = TR_132 ;
	7'h61 :
		RG_rl_120_t1 = TR_132 ;
	7'h62 :
		RG_rl_120_t1 = TR_132 ;
	7'h63 :
		RG_rl_120_t1 = TR_132 ;
	7'h64 :
		RG_rl_120_t1 = TR_132 ;
	7'h65 :
		RG_rl_120_t1 = TR_132 ;
	7'h66 :
		RG_rl_120_t1 = TR_132 ;
	7'h67 :
		RG_rl_120_t1 = TR_132 ;
	7'h68 :
		RG_rl_120_t1 = TR_132 ;
	7'h69 :
		RG_rl_120_t1 = TR_132 ;
	7'h6a :
		RG_rl_120_t1 = TR_132 ;
	7'h6b :
		RG_rl_120_t1 = TR_132 ;
	7'h6c :
		RG_rl_120_t1 = TR_132 ;
	7'h6d :
		RG_rl_120_t1 = TR_132 ;
	7'h6e :
		RG_rl_120_t1 = TR_132 ;
	7'h6f :
		RG_rl_120_t1 = TR_132 ;
	7'h70 :
		RG_rl_120_t1 = TR_132 ;
	7'h71 :
		RG_rl_120_t1 = TR_132 ;
	7'h72 :
		RG_rl_120_t1 = TR_132 ;
	7'h73 :
		RG_rl_120_t1 = TR_132 ;
	7'h74 :
		RG_rl_120_t1 = TR_132 ;
	7'h75 :
		RG_rl_120_t1 = TR_132 ;
	7'h76 :
		RG_rl_120_t1 = TR_132 ;
	7'h77 :
		RG_rl_120_t1 = TR_132 ;
	7'h78 :
		RG_rl_120_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h79 :
		RG_rl_120_t1 = TR_132 ;
	7'h7a :
		RG_rl_120_t1 = TR_132 ;
	7'h7b :
		RG_rl_120_t1 = TR_132 ;
	7'h7c :
		RG_rl_120_t1 = TR_132 ;
	7'h7d :
		RG_rl_120_t1 = TR_132 ;
	7'h7e :
		RG_rl_120_t1 = TR_132 ;
	7'h7f :
		RG_rl_120_t1 = TR_132 ;
	default :
		RG_rl_120_t1 = 9'hx ;
	endcase
always @ ( RG_rl_120_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_244 or M_318 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_120_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h78 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_120_t = ( ( { 9{ M_318 } } & RG_rl_244 )
		| ( { 9{ U_569 } } & RG_rl_120_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_120_en = ( M_318 | RG_rl_120_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_120_en )
		RG_rl_120 <= RG_rl_120_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_133 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_121_t1 = TR_133 ;
	7'h01 :
		RG_rl_121_t1 = TR_133 ;
	7'h02 :
		RG_rl_121_t1 = TR_133 ;
	7'h03 :
		RG_rl_121_t1 = TR_133 ;
	7'h04 :
		RG_rl_121_t1 = TR_133 ;
	7'h05 :
		RG_rl_121_t1 = TR_133 ;
	7'h06 :
		RG_rl_121_t1 = TR_133 ;
	7'h07 :
		RG_rl_121_t1 = TR_133 ;
	7'h08 :
		RG_rl_121_t1 = TR_133 ;
	7'h09 :
		RG_rl_121_t1 = TR_133 ;
	7'h0a :
		RG_rl_121_t1 = TR_133 ;
	7'h0b :
		RG_rl_121_t1 = TR_133 ;
	7'h0c :
		RG_rl_121_t1 = TR_133 ;
	7'h0d :
		RG_rl_121_t1 = TR_133 ;
	7'h0e :
		RG_rl_121_t1 = TR_133 ;
	7'h0f :
		RG_rl_121_t1 = TR_133 ;
	7'h10 :
		RG_rl_121_t1 = TR_133 ;
	7'h11 :
		RG_rl_121_t1 = TR_133 ;
	7'h12 :
		RG_rl_121_t1 = TR_133 ;
	7'h13 :
		RG_rl_121_t1 = TR_133 ;
	7'h14 :
		RG_rl_121_t1 = TR_133 ;
	7'h15 :
		RG_rl_121_t1 = TR_133 ;
	7'h16 :
		RG_rl_121_t1 = TR_133 ;
	7'h17 :
		RG_rl_121_t1 = TR_133 ;
	7'h18 :
		RG_rl_121_t1 = TR_133 ;
	7'h19 :
		RG_rl_121_t1 = TR_133 ;
	7'h1a :
		RG_rl_121_t1 = TR_133 ;
	7'h1b :
		RG_rl_121_t1 = TR_133 ;
	7'h1c :
		RG_rl_121_t1 = TR_133 ;
	7'h1d :
		RG_rl_121_t1 = TR_133 ;
	7'h1e :
		RG_rl_121_t1 = TR_133 ;
	7'h1f :
		RG_rl_121_t1 = TR_133 ;
	7'h20 :
		RG_rl_121_t1 = TR_133 ;
	7'h21 :
		RG_rl_121_t1 = TR_133 ;
	7'h22 :
		RG_rl_121_t1 = TR_133 ;
	7'h23 :
		RG_rl_121_t1 = TR_133 ;
	7'h24 :
		RG_rl_121_t1 = TR_133 ;
	7'h25 :
		RG_rl_121_t1 = TR_133 ;
	7'h26 :
		RG_rl_121_t1 = TR_133 ;
	7'h27 :
		RG_rl_121_t1 = TR_133 ;
	7'h28 :
		RG_rl_121_t1 = TR_133 ;
	7'h29 :
		RG_rl_121_t1 = TR_133 ;
	7'h2a :
		RG_rl_121_t1 = TR_133 ;
	7'h2b :
		RG_rl_121_t1 = TR_133 ;
	7'h2c :
		RG_rl_121_t1 = TR_133 ;
	7'h2d :
		RG_rl_121_t1 = TR_133 ;
	7'h2e :
		RG_rl_121_t1 = TR_133 ;
	7'h2f :
		RG_rl_121_t1 = TR_133 ;
	7'h30 :
		RG_rl_121_t1 = TR_133 ;
	7'h31 :
		RG_rl_121_t1 = TR_133 ;
	7'h32 :
		RG_rl_121_t1 = TR_133 ;
	7'h33 :
		RG_rl_121_t1 = TR_133 ;
	7'h34 :
		RG_rl_121_t1 = TR_133 ;
	7'h35 :
		RG_rl_121_t1 = TR_133 ;
	7'h36 :
		RG_rl_121_t1 = TR_133 ;
	7'h37 :
		RG_rl_121_t1 = TR_133 ;
	7'h38 :
		RG_rl_121_t1 = TR_133 ;
	7'h39 :
		RG_rl_121_t1 = TR_133 ;
	7'h3a :
		RG_rl_121_t1 = TR_133 ;
	7'h3b :
		RG_rl_121_t1 = TR_133 ;
	7'h3c :
		RG_rl_121_t1 = TR_133 ;
	7'h3d :
		RG_rl_121_t1 = TR_133 ;
	7'h3e :
		RG_rl_121_t1 = TR_133 ;
	7'h3f :
		RG_rl_121_t1 = TR_133 ;
	7'h40 :
		RG_rl_121_t1 = TR_133 ;
	7'h41 :
		RG_rl_121_t1 = TR_133 ;
	7'h42 :
		RG_rl_121_t1 = TR_133 ;
	7'h43 :
		RG_rl_121_t1 = TR_133 ;
	7'h44 :
		RG_rl_121_t1 = TR_133 ;
	7'h45 :
		RG_rl_121_t1 = TR_133 ;
	7'h46 :
		RG_rl_121_t1 = TR_133 ;
	7'h47 :
		RG_rl_121_t1 = TR_133 ;
	7'h48 :
		RG_rl_121_t1 = TR_133 ;
	7'h49 :
		RG_rl_121_t1 = TR_133 ;
	7'h4a :
		RG_rl_121_t1 = TR_133 ;
	7'h4b :
		RG_rl_121_t1 = TR_133 ;
	7'h4c :
		RG_rl_121_t1 = TR_133 ;
	7'h4d :
		RG_rl_121_t1 = TR_133 ;
	7'h4e :
		RG_rl_121_t1 = TR_133 ;
	7'h4f :
		RG_rl_121_t1 = TR_133 ;
	7'h50 :
		RG_rl_121_t1 = TR_133 ;
	7'h51 :
		RG_rl_121_t1 = TR_133 ;
	7'h52 :
		RG_rl_121_t1 = TR_133 ;
	7'h53 :
		RG_rl_121_t1 = TR_133 ;
	7'h54 :
		RG_rl_121_t1 = TR_133 ;
	7'h55 :
		RG_rl_121_t1 = TR_133 ;
	7'h56 :
		RG_rl_121_t1 = TR_133 ;
	7'h57 :
		RG_rl_121_t1 = TR_133 ;
	7'h58 :
		RG_rl_121_t1 = TR_133 ;
	7'h59 :
		RG_rl_121_t1 = TR_133 ;
	7'h5a :
		RG_rl_121_t1 = TR_133 ;
	7'h5b :
		RG_rl_121_t1 = TR_133 ;
	7'h5c :
		RG_rl_121_t1 = TR_133 ;
	7'h5d :
		RG_rl_121_t1 = TR_133 ;
	7'h5e :
		RG_rl_121_t1 = TR_133 ;
	7'h5f :
		RG_rl_121_t1 = TR_133 ;
	7'h60 :
		RG_rl_121_t1 = TR_133 ;
	7'h61 :
		RG_rl_121_t1 = TR_133 ;
	7'h62 :
		RG_rl_121_t1 = TR_133 ;
	7'h63 :
		RG_rl_121_t1 = TR_133 ;
	7'h64 :
		RG_rl_121_t1 = TR_133 ;
	7'h65 :
		RG_rl_121_t1 = TR_133 ;
	7'h66 :
		RG_rl_121_t1 = TR_133 ;
	7'h67 :
		RG_rl_121_t1 = TR_133 ;
	7'h68 :
		RG_rl_121_t1 = TR_133 ;
	7'h69 :
		RG_rl_121_t1 = TR_133 ;
	7'h6a :
		RG_rl_121_t1 = TR_133 ;
	7'h6b :
		RG_rl_121_t1 = TR_133 ;
	7'h6c :
		RG_rl_121_t1 = TR_133 ;
	7'h6d :
		RG_rl_121_t1 = TR_133 ;
	7'h6e :
		RG_rl_121_t1 = TR_133 ;
	7'h6f :
		RG_rl_121_t1 = TR_133 ;
	7'h70 :
		RG_rl_121_t1 = TR_133 ;
	7'h71 :
		RG_rl_121_t1 = TR_133 ;
	7'h72 :
		RG_rl_121_t1 = TR_133 ;
	7'h73 :
		RG_rl_121_t1 = TR_133 ;
	7'h74 :
		RG_rl_121_t1 = TR_133 ;
	7'h75 :
		RG_rl_121_t1 = TR_133 ;
	7'h76 :
		RG_rl_121_t1 = TR_133 ;
	7'h77 :
		RG_rl_121_t1 = TR_133 ;
	7'h78 :
		RG_rl_121_t1 = TR_133 ;
	7'h79 :
		RG_rl_121_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7a :
		RG_rl_121_t1 = TR_133 ;
	7'h7b :
		RG_rl_121_t1 = TR_133 ;
	7'h7c :
		RG_rl_121_t1 = TR_133 ;
	7'h7d :
		RG_rl_121_t1 = TR_133 ;
	7'h7e :
		RG_rl_121_t1 = TR_133 ;
	7'h7f :
		RG_rl_121_t1 = TR_133 ;
	default :
		RG_rl_121_t1 = 9'hx ;
	endcase
always @ ( RG_rl_121_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_59 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_121_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h79 ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_121_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_59 )
		| ( { 9{ U_569 } } & RG_rl_121_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_121_en = ( U_570 | RG_rl_121_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_121_en )
		RG_rl_121 <= RG_rl_121_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_134 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_122_t1 = TR_134 ;
	7'h01 :
		RG_rl_122_t1 = TR_134 ;
	7'h02 :
		RG_rl_122_t1 = TR_134 ;
	7'h03 :
		RG_rl_122_t1 = TR_134 ;
	7'h04 :
		RG_rl_122_t1 = TR_134 ;
	7'h05 :
		RG_rl_122_t1 = TR_134 ;
	7'h06 :
		RG_rl_122_t1 = TR_134 ;
	7'h07 :
		RG_rl_122_t1 = TR_134 ;
	7'h08 :
		RG_rl_122_t1 = TR_134 ;
	7'h09 :
		RG_rl_122_t1 = TR_134 ;
	7'h0a :
		RG_rl_122_t1 = TR_134 ;
	7'h0b :
		RG_rl_122_t1 = TR_134 ;
	7'h0c :
		RG_rl_122_t1 = TR_134 ;
	7'h0d :
		RG_rl_122_t1 = TR_134 ;
	7'h0e :
		RG_rl_122_t1 = TR_134 ;
	7'h0f :
		RG_rl_122_t1 = TR_134 ;
	7'h10 :
		RG_rl_122_t1 = TR_134 ;
	7'h11 :
		RG_rl_122_t1 = TR_134 ;
	7'h12 :
		RG_rl_122_t1 = TR_134 ;
	7'h13 :
		RG_rl_122_t1 = TR_134 ;
	7'h14 :
		RG_rl_122_t1 = TR_134 ;
	7'h15 :
		RG_rl_122_t1 = TR_134 ;
	7'h16 :
		RG_rl_122_t1 = TR_134 ;
	7'h17 :
		RG_rl_122_t1 = TR_134 ;
	7'h18 :
		RG_rl_122_t1 = TR_134 ;
	7'h19 :
		RG_rl_122_t1 = TR_134 ;
	7'h1a :
		RG_rl_122_t1 = TR_134 ;
	7'h1b :
		RG_rl_122_t1 = TR_134 ;
	7'h1c :
		RG_rl_122_t1 = TR_134 ;
	7'h1d :
		RG_rl_122_t1 = TR_134 ;
	7'h1e :
		RG_rl_122_t1 = TR_134 ;
	7'h1f :
		RG_rl_122_t1 = TR_134 ;
	7'h20 :
		RG_rl_122_t1 = TR_134 ;
	7'h21 :
		RG_rl_122_t1 = TR_134 ;
	7'h22 :
		RG_rl_122_t1 = TR_134 ;
	7'h23 :
		RG_rl_122_t1 = TR_134 ;
	7'h24 :
		RG_rl_122_t1 = TR_134 ;
	7'h25 :
		RG_rl_122_t1 = TR_134 ;
	7'h26 :
		RG_rl_122_t1 = TR_134 ;
	7'h27 :
		RG_rl_122_t1 = TR_134 ;
	7'h28 :
		RG_rl_122_t1 = TR_134 ;
	7'h29 :
		RG_rl_122_t1 = TR_134 ;
	7'h2a :
		RG_rl_122_t1 = TR_134 ;
	7'h2b :
		RG_rl_122_t1 = TR_134 ;
	7'h2c :
		RG_rl_122_t1 = TR_134 ;
	7'h2d :
		RG_rl_122_t1 = TR_134 ;
	7'h2e :
		RG_rl_122_t1 = TR_134 ;
	7'h2f :
		RG_rl_122_t1 = TR_134 ;
	7'h30 :
		RG_rl_122_t1 = TR_134 ;
	7'h31 :
		RG_rl_122_t1 = TR_134 ;
	7'h32 :
		RG_rl_122_t1 = TR_134 ;
	7'h33 :
		RG_rl_122_t1 = TR_134 ;
	7'h34 :
		RG_rl_122_t1 = TR_134 ;
	7'h35 :
		RG_rl_122_t1 = TR_134 ;
	7'h36 :
		RG_rl_122_t1 = TR_134 ;
	7'h37 :
		RG_rl_122_t1 = TR_134 ;
	7'h38 :
		RG_rl_122_t1 = TR_134 ;
	7'h39 :
		RG_rl_122_t1 = TR_134 ;
	7'h3a :
		RG_rl_122_t1 = TR_134 ;
	7'h3b :
		RG_rl_122_t1 = TR_134 ;
	7'h3c :
		RG_rl_122_t1 = TR_134 ;
	7'h3d :
		RG_rl_122_t1 = TR_134 ;
	7'h3e :
		RG_rl_122_t1 = TR_134 ;
	7'h3f :
		RG_rl_122_t1 = TR_134 ;
	7'h40 :
		RG_rl_122_t1 = TR_134 ;
	7'h41 :
		RG_rl_122_t1 = TR_134 ;
	7'h42 :
		RG_rl_122_t1 = TR_134 ;
	7'h43 :
		RG_rl_122_t1 = TR_134 ;
	7'h44 :
		RG_rl_122_t1 = TR_134 ;
	7'h45 :
		RG_rl_122_t1 = TR_134 ;
	7'h46 :
		RG_rl_122_t1 = TR_134 ;
	7'h47 :
		RG_rl_122_t1 = TR_134 ;
	7'h48 :
		RG_rl_122_t1 = TR_134 ;
	7'h49 :
		RG_rl_122_t1 = TR_134 ;
	7'h4a :
		RG_rl_122_t1 = TR_134 ;
	7'h4b :
		RG_rl_122_t1 = TR_134 ;
	7'h4c :
		RG_rl_122_t1 = TR_134 ;
	7'h4d :
		RG_rl_122_t1 = TR_134 ;
	7'h4e :
		RG_rl_122_t1 = TR_134 ;
	7'h4f :
		RG_rl_122_t1 = TR_134 ;
	7'h50 :
		RG_rl_122_t1 = TR_134 ;
	7'h51 :
		RG_rl_122_t1 = TR_134 ;
	7'h52 :
		RG_rl_122_t1 = TR_134 ;
	7'h53 :
		RG_rl_122_t1 = TR_134 ;
	7'h54 :
		RG_rl_122_t1 = TR_134 ;
	7'h55 :
		RG_rl_122_t1 = TR_134 ;
	7'h56 :
		RG_rl_122_t1 = TR_134 ;
	7'h57 :
		RG_rl_122_t1 = TR_134 ;
	7'h58 :
		RG_rl_122_t1 = TR_134 ;
	7'h59 :
		RG_rl_122_t1 = TR_134 ;
	7'h5a :
		RG_rl_122_t1 = TR_134 ;
	7'h5b :
		RG_rl_122_t1 = TR_134 ;
	7'h5c :
		RG_rl_122_t1 = TR_134 ;
	7'h5d :
		RG_rl_122_t1 = TR_134 ;
	7'h5e :
		RG_rl_122_t1 = TR_134 ;
	7'h5f :
		RG_rl_122_t1 = TR_134 ;
	7'h60 :
		RG_rl_122_t1 = TR_134 ;
	7'h61 :
		RG_rl_122_t1 = TR_134 ;
	7'h62 :
		RG_rl_122_t1 = TR_134 ;
	7'h63 :
		RG_rl_122_t1 = TR_134 ;
	7'h64 :
		RG_rl_122_t1 = TR_134 ;
	7'h65 :
		RG_rl_122_t1 = TR_134 ;
	7'h66 :
		RG_rl_122_t1 = TR_134 ;
	7'h67 :
		RG_rl_122_t1 = TR_134 ;
	7'h68 :
		RG_rl_122_t1 = TR_134 ;
	7'h69 :
		RG_rl_122_t1 = TR_134 ;
	7'h6a :
		RG_rl_122_t1 = TR_134 ;
	7'h6b :
		RG_rl_122_t1 = TR_134 ;
	7'h6c :
		RG_rl_122_t1 = TR_134 ;
	7'h6d :
		RG_rl_122_t1 = TR_134 ;
	7'h6e :
		RG_rl_122_t1 = TR_134 ;
	7'h6f :
		RG_rl_122_t1 = TR_134 ;
	7'h70 :
		RG_rl_122_t1 = TR_134 ;
	7'h71 :
		RG_rl_122_t1 = TR_134 ;
	7'h72 :
		RG_rl_122_t1 = TR_134 ;
	7'h73 :
		RG_rl_122_t1 = TR_134 ;
	7'h74 :
		RG_rl_122_t1 = TR_134 ;
	7'h75 :
		RG_rl_122_t1 = TR_134 ;
	7'h76 :
		RG_rl_122_t1 = TR_134 ;
	7'h77 :
		RG_rl_122_t1 = TR_134 ;
	7'h78 :
		RG_rl_122_t1 = TR_134 ;
	7'h79 :
		RG_rl_122_t1 = TR_134 ;
	7'h7a :
		RG_rl_122_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7b :
		RG_rl_122_t1 = TR_134 ;
	7'h7c :
		RG_rl_122_t1 = TR_134 ;
	7'h7d :
		RG_rl_122_t1 = TR_134 ;
	7'h7e :
		RG_rl_122_t1 = TR_134 ;
	7'h7f :
		RG_rl_122_t1 = TR_134 ;
	default :
		RG_rl_122_t1 = 9'hx ;
	endcase
always @ ( RG_rl_122_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_245 or M_318 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_122_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h7a ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_122_t = ( ( { 9{ M_318 } } & RG_rl_245 )
		| ( { 9{ U_569 } } & RG_rl_122_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_122_en = ( M_318 | RG_rl_122_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_122_en )
		RG_rl_122 <= RG_rl_122_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_135 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_123_t1 = TR_135 ;
	7'h01 :
		RG_rl_123_t1 = TR_135 ;
	7'h02 :
		RG_rl_123_t1 = TR_135 ;
	7'h03 :
		RG_rl_123_t1 = TR_135 ;
	7'h04 :
		RG_rl_123_t1 = TR_135 ;
	7'h05 :
		RG_rl_123_t1 = TR_135 ;
	7'h06 :
		RG_rl_123_t1 = TR_135 ;
	7'h07 :
		RG_rl_123_t1 = TR_135 ;
	7'h08 :
		RG_rl_123_t1 = TR_135 ;
	7'h09 :
		RG_rl_123_t1 = TR_135 ;
	7'h0a :
		RG_rl_123_t1 = TR_135 ;
	7'h0b :
		RG_rl_123_t1 = TR_135 ;
	7'h0c :
		RG_rl_123_t1 = TR_135 ;
	7'h0d :
		RG_rl_123_t1 = TR_135 ;
	7'h0e :
		RG_rl_123_t1 = TR_135 ;
	7'h0f :
		RG_rl_123_t1 = TR_135 ;
	7'h10 :
		RG_rl_123_t1 = TR_135 ;
	7'h11 :
		RG_rl_123_t1 = TR_135 ;
	7'h12 :
		RG_rl_123_t1 = TR_135 ;
	7'h13 :
		RG_rl_123_t1 = TR_135 ;
	7'h14 :
		RG_rl_123_t1 = TR_135 ;
	7'h15 :
		RG_rl_123_t1 = TR_135 ;
	7'h16 :
		RG_rl_123_t1 = TR_135 ;
	7'h17 :
		RG_rl_123_t1 = TR_135 ;
	7'h18 :
		RG_rl_123_t1 = TR_135 ;
	7'h19 :
		RG_rl_123_t1 = TR_135 ;
	7'h1a :
		RG_rl_123_t1 = TR_135 ;
	7'h1b :
		RG_rl_123_t1 = TR_135 ;
	7'h1c :
		RG_rl_123_t1 = TR_135 ;
	7'h1d :
		RG_rl_123_t1 = TR_135 ;
	7'h1e :
		RG_rl_123_t1 = TR_135 ;
	7'h1f :
		RG_rl_123_t1 = TR_135 ;
	7'h20 :
		RG_rl_123_t1 = TR_135 ;
	7'h21 :
		RG_rl_123_t1 = TR_135 ;
	7'h22 :
		RG_rl_123_t1 = TR_135 ;
	7'h23 :
		RG_rl_123_t1 = TR_135 ;
	7'h24 :
		RG_rl_123_t1 = TR_135 ;
	7'h25 :
		RG_rl_123_t1 = TR_135 ;
	7'h26 :
		RG_rl_123_t1 = TR_135 ;
	7'h27 :
		RG_rl_123_t1 = TR_135 ;
	7'h28 :
		RG_rl_123_t1 = TR_135 ;
	7'h29 :
		RG_rl_123_t1 = TR_135 ;
	7'h2a :
		RG_rl_123_t1 = TR_135 ;
	7'h2b :
		RG_rl_123_t1 = TR_135 ;
	7'h2c :
		RG_rl_123_t1 = TR_135 ;
	7'h2d :
		RG_rl_123_t1 = TR_135 ;
	7'h2e :
		RG_rl_123_t1 = TR_135 ;
	7'h2f :
		RG_rl_123_t1 = TR_135 ;
	7'h30 :
		RG_rl_123_t1 = TR_135 ;
	7'h31 :
		RG_rl_123_t1 = TR_135 ;
	7'h32 :
		RG_rl_123_t1 = TR_135 ;
	7'h33 :
		RG_rl_123_t1 = TR_135 ;
	7'h34 :
		RG_rl_123_t1 = TR_135 ;
	7'h35 :
		RG_rl_123_t1 = TR_135 ;
	7'h36 :
		RG_rl_123_t1 = TR_135 ;
	7'h37 :
		RG_rl_123_t1 = TR_135 ;
	7'h38 :
		RG_rl_123_t1 = TR_135 ;
	7'h39 :
		RG_rl_123_t1 = TR_135 ;
	7'h3a :
		RG_rl_123_t1 = TR_135 ;
	7'h3b :
		RG_rl_123_t1 = TR_135 ;
	7'h3c :
		RG_rl_123_t1 = TR_135 ;
	7'h3d :
		RG_rl_123_t1 = TR_135 ;
	7'h3e :
		RG_rl_123_t1 = TR_135 ;
	7'h3f :
		RG_rl_123_t1 = TR_135 ;
	7'h40 :
		RG_rl_123_t1 = TR_135 ;
	7'h41 :
		RG_rl_123_t1 = TR_135 ;
	7'h42 :
		RG_rl_123_t1 = TR_135 ;
	7'h43 :
		RG_rl_123_t1 = TR_135 ;
	7'h44 :
		RG_rl_123_t1 = TR_135 ;
	7'h45 :
		RG_rl_123_t1 = TR_135 ;
	7'h46 :
		RG_rl_123_t1 = TR_135 ;
	7'h47 :
		RG_rl_123_t1 = TR_135 ;
	7'h48 :
		RG_rl_123_t1 = TR_135 ;
	7'h49 :
		RG_rl_123_t1 = TR_135 ;
	7'h4a :
		RG_rl_123_t1 = TR_135 ;
	7'h4b :
		RG_rl_123_t1 = TR_135 ;
	7'h4c :
		RG_rl_123_t1 = TR_135 ;
	7'h4d :
		RG_rl_123_t1 = TR_135 ;
	7'h4e :
		RG_rl_123_t1 = TR_135 ;
	7'h4f :
		RG_rl_123_t1 = TR_135 ;
	7'h50 :
		RG_rl_123_t1 = TR_135 ;
	7'h51 :
		RG_rl_123_t1 = TR_135 ;
	7'h52 :
		RG_rl_123_t1 = TR_135 ;
	7'h53 :
		RG_rl_123_t1 = TR_135 ;
	7'h54 :
		RG_rl_123_t1 = TR_135 ;
	7'h55 :
		RG_rl_123_t1 = TR_135 ;
	7'h56 :
		RG_rl_123_t1 = TR_135 ;
	7'h57 :
		RG_rl_123_t1 = TR_135 ;
	7'h58 :
		RG_rl_123_t1 = TR_135 ;
	7'h59 :
		RG_rl_123_t1 = TR_135 ;
	7'h5a :
		RG_rl_123_t1 = TR_135 ;
	7'h5b :
		RG_rl_123_t1 = TR_135 ;
	7'h5c :
		RG_rl_123_t1 = TR_135 ;
	7'h5d :
		RG_rl_123_t1 = TR_135 ;
	7'h5e :
		RG_rl_123_t1 = TR_135 ;
	7'h5f :
		RG_rl_123_t1 = TR_135 ;
	7'h60 :
		RG_rl_123_t1 = TR_135 ;
	7'h61 :
		RG_rl_123_t1 = TR_135 ;
	7'h62 :
		RG_rl_123_t1 = TR_135 ;
	7'h63 :
		RG_rl_123_t1 = TR_135 ;
	7'h64 :
		RG_rl_123_t1 = TR_135 ;
	7'h65 :
		RG_rl_123_t1 = TR_135 ;
	7'h66 :
		RG_rl_123_t1 = TR_135 ;
	7'h67 :
		RG_rl_123_t1 = TR_135 ;
	7'h68 :
		RG_rl_123_t1 = TR_135 ;
	7'h69 :
		RG_rl_123_t1 = TR_135 ;
	7'h6a :
		RG_rl_123_t1 = TR_135 ;
	7'h6b :
		RG_rl_123_t1 = TR_135 ;
	7'h6c :
		RG_rl_123_t1 = TR_135 ;
	7'h6d :
		RG_rl_123_t1 = TR_135 ;
	7'h6e :
		RG_rl_123_t1 = TR_135 ;
	7'h6f :
		RG_rl_123_t1 = TR_135 ;
	7'h70 :
		RG_rl_123_t1 = TR_135 ;
	7'h71 :
		RG_rl_123_t1 = TR_135 ;
	7'h72 :
		RG_rl_123_t1 = TR_135 ;
	7'h73 :
		RG_rl_123_t1 = TR_135 ;
	7'h74 :
		RG_rl_123_t1 = TR_135 ;
	7'h75 :
		RG_rl_123_t1 = TR_135 ;
	7'h76 :
		RG_rl_123_t1 = TR_135 ;
	7'h77 :
		RG_rl_123_t1 = TR_135 ;
	7'h78 :
		RG_rl_123_t1 = TR_135 ;
	7'h79 :
		RG_rl_123_t1 = TR_135 ;
	7'h7a :
		RG_rl_123_t1 = TR_135 ;
	7'h7b :
		RG_rl_123_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7c :
		RG_rl_123_t1 = TR_135 ;
	7'h7d :
		RG_rl_123_t1 = TR_135 ;
	7'h7e :
		RG_rl_123_t1 = TR_135 ;
	7'h7f :
		RG_rl_123_t1 = TR_135 ;
	default :
		RG_rl_123_t1 = 9'hx ;
	endcase
always @ ( RG_rl_123_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_60 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_123_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h7b ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_123_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_60 )
		| ( { 9{ U_569 } } & RG_rl_123_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_123_en = ( U_570 | RG_rl_123_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_123_en )
		RG_rl_123 <= RG_rl_123_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_136 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_124_t1 = TR_136 ;
	7'h01 :
		RG_rl_124_t1 = TR_136 ;
	7'h02 :
		RG_rl_124_t1 = TR_136 ;
	7'h03 :
		RG_rl_124_t1 = TR_136 ;
	7'h04 :
		RG_rl_124_t1 = TR_136 ;
	7'h05 :
		RG_rl_124_t1 = TR_136 ;
	7'h06 :
		RG_rl_124_t1 = TR_136 ;
	7'h07 :
		RG_rl_124_t1 = TR_136 ;
	7'h08 :
		RG_rl_124_t1 = TR_136 ;
	7'h09 :
		RG_rl_124_t1 = TR_136 ;
	7'h0a :
		RG_rl_124_t1 = TR_136 ;
	7'h0b :
		RG_rl_124_t1 = TR_136 ;
	7'h0c :
		RG_rl_124_t1 = TR_136 ;
	7'h0d :
		RG_rl_124_t1 = TR_136 ;
	7'h0e :
		RG_rl_124_t1 = TR_136 ;
	7'h0f :
		RG_rl_124_t1 = TR_136 ;
	7'h10 :
		RG_rl_124_t1 = TR_136 ;
	7'h11 :
		RG_rl_124_t1 = TR_136 ;
	7'h12 :
		RG_rl_124_t1 = TR_136 ;
	7'h13 :
		RG_rl_124_t1 = TR_136 ;
	7'h14 :
		RG_rl_124_t1 = TR_136 ;
	7'h15 :
		RG_rl_124_t1 = TR_136 ;
	7'h16 :
		RG_rl_124_t1 = TR_136 ;
	7'h17 :
		RG_rl_124_t1 = TR_136 ;
	7'h18 :
		RG_rl_124_t1 = TR_136 ;
	7'h19 :
		RG_rl_124_t1 = TR_136 ;
	7'h1a :
		RG_rl_124_t1 = TR_136 ;
	7'h1b :
		RG_rl_124_t1 = TR_136 ;
	7'h1c :
		RG_rl_124_t1 = TR_136 ;
	7'h1d :
		RG_rl_124_t1 = TR_136 ;
	7'h1e :
		RG_rl_124_t1 = TR_136 ;
	7'h1f :
		RG_rl_124_t1 = TR_136 ;
	7'h20 :
		RG_rl_124_t1 = TR_136 ;
	7'h21 :
		RG_rl_124_t1 = TR_136 ;
	7'h22 :
		RG_rl_124_t1 = TR_136 ;
	7'h23 :
		RG_rl_124_t1 = TR_136 ;
	7'h24 :
		RG_rl_124_t1 = TR_136 ;
	7'h25 :
		RG_rl_124_t1 = TR_136 ;
	7'h26 :
		RG_rl_124_t1 = TR_136 ;
	7'h27 :
		RG_rl_124_t1 = TR_136 ;
	7'h28 :
		RG_rl_124_t1 = TR_136 ;
	7'h29 :
		RG_rl_124_t1 = TR_136 ;
	7'h2a :
		RG_rl_124_t1 = TR_136 ;
	7'h2b :
		RG_rl_124_t1 = TR_136 ;
	7'h2c :
		RG_rl_124_t1 = TR_136 ;
	7'h2d :
		RG_rl_124_t1 = TR_136 ;
	7'h2e :
		RG_rl_124_t1 = TR_136 ;
	7'h2f :
		RG_rl_124_t1 = TR_136 ;
	7'h30 :
		RG_rl_124_t1 = TR_136 ;
	7'h31 :
		RG_rl_124_t1 = TR_136 ;
	7'h32 :
		RG_rl_124_t1 = TR_136 ;
	7'h33 :
		RG_rl_124_t1 = TR_136 ;
	7'h34 :
		RG_rl_124_t1 = TR_136 ;
	7'h35 :
		RG_rl_124_t1 = TR_136 ;
	7'h36 :
		RG_rl_124_t1 = TR_136 ;
	7'h37 :
		RG_rl_124_t1 = TR_136 ;
	7'h38 :
		RG_rl_124_t1 = TR_136 ;
	7'h39 :
		RG_rl_124_t1 = TR_136 ;
	7'h3a :
		RG_rl_124_t1 = TR_136 ;
	7'h3b :
		RG_rl_124_t1 = TR_136 ;
	7'h3c :
		RG_rl_124_t1 = TR_136 ;
	7'h3d :
		RG_rl_124_t1 = TR_136 ;
	7'h3e :
		RG_rl_124_t1 = TR_136 ;
	7'h3f :
		RG_rl_124_t1 = TR_136 ;
	7'h40 :
		RG_rl_124_t1 = TR_136 ;
	7'h41 :
		RG_rl_124_t1 = TR_136 ;
	7'h42 :
		RG_rl_124_t1 = TR_136 ;
	7'h43 :
		RG_rl_124_t1 = TR_136 ;
	7'h44 :
		RG_rl_124_t1 = TR_136 ;
	7'h45 :
		RG_rl_124_t1 = TR_136 ;
	7'h46 :
		RG_rl_124_t1 = TR_136 ;
	7'h47 :
		RG_rl_124_t1 = TR_136 ;
	7'h48 :
		RG_rl_124_t1 = TR_136 ;
	7'h49 :
		RG_rl_124_t1 = TR_136 ;
	7'h4a :
		RG_rl_124_t1 = TR_136 ;
	7'h4b :
		RG_rl_124_t1 = TR_136 ;
	7'h4c :
		RG_rl_124_t1 = TR_136 ;
	7'h4d :
		RG_rl_124_t1 = TR_136 ;
	7'h4e :
		RG_rl_124_t1 = TR_136 ;
	7'h4f :
		RG_rl_124_t1 = TR_136 ;
	7'h50 :
		RG_rl_124_t1 = TR_136 ;
	7'h51 :
		RG_rl_124_t1 = TR_136 ;
	7'h52 :
		RG_rl_124_t1 = TR_136 ;
	7'h53 :
		RG_rl_124_t1 = TR_136 ;
	7'h54 :
		RG_rl_124_t1 = TR_136 ;
	7'h55 :
		RG_rl_124_t1 = TR_136 ;
	7'h56 :
		RG_rl_124_t1 = TR_136 ;
	7'h57 :
		RG_rl_124_t1 = TR_136 ;
	7'h58 :
		RG_rl_124_t1 = TR_136 ;
	7'h59 :
		RG_rl_124_t1 = TR_136 ;
	7'h5a :
		RG_rl_124_t1 = TR_136 ;
	7'h5b :
		RG_rl_124_t1 = TR_136 ;
	7'h5c :
		RG_rl_124_t1 = TR_136 ;
	7'h5d :
		RG_rl_124_t1 = TR_136 ;
	7'h5e :
		RG_rl_124_t1 = TR_136 ;
	7'h5f :
		RG_rl_124_t1 = TR_136 ;
	7'h60 :
		RG_rl_124_t1 = TR_136 ;
	7'h61 :
		RG_rl_124_t1 = TR_136 ;
	7'h62 :
		RG_rl_124_t1 = TR_136 ;
	7'h63 :
		RG_rl_124_t1 = TR_136 ;
	7'h64 :
		RG_rl_124_t1 = TR_136 ;
	7'h65 :
		RG_rl_124_t1 = TR_136 ;
	7'h66 :
		RG_rl_124_t1 = TR_136 ;
	7'h67 :
		RG_rl_124_t1 = TR_136 ;
	7'h68 :
		RG_rl_124_t1 = TR_136 ;
	7'h69 :
		RG_rl_124_t1 = TR_136 ;
	7'h6a :
		RG_rl_124_t1 = TR_136 ;
	7'h6b :
		RG_rl_124_t1 = TR_136 ;
	7'h6c :
		RG_rl_124_t1 = TR_136 ;
	7'h6d :
		RG_rl_124_t1 = TR_136 ;
	7'h6e :
		RG_rl_124_t1 = TR_136 ;
	7'h6f :
		RG_rl_124_t1 = TR_136 ;
	7'h70 :
		RG_rl_124_t1 = TR_136 ;
	7'h71 :
		RG_rl_124_t1 = TR_136 ;
	7'h72 :
		RG_rl_124_t1 = TR_136 ;
	7'h73 :
		RG_rl_124_t1 = TR_136 ;
	7'h74 :
		RG_rl_124_t1 = TR_136 ;
	7'h75 :
		RG_rl_124_t1 = TR_136 ;
	7'h76 :
		RG_rl_124_t1 = TR_136 ;
	7'h77 :
		RG_rl_124_t1 = TR_136 ;
	7'h78 :
		RG_rl_124_t1 = TR_136 ;
	7'h79 :
		RG_rl_124_t1 = TR_136 ;
	7'h7a :
		RG_rl_124_t1 = TR_136 ;
	7'h7b :
		RG_rl_124_t1 = TR_136 ;
	7'h7c :
		RG_rl_124_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7d :
		RG_rl_124_t1 = TR_136 ;
	7'h7e :
		RG_rl_124_t1 = TR_136 ;
	7'h7f :
		RG_rl_124_t1 = TR_136 ;
	default :
		RG_rl_124_t1 = 9'hx ;
	endcase
always @ ( RG_rl_124_t1 or U_569 or sub8u_71ot or U_571 or RG_rl_246 or M_318 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_124_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h7c ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_124_t = ( ( { 9{ M_318 } } & RG_rl_246 )
		| ( { 9{ U_569 } } & RG_rl_124_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_124_en = ( M_318 | RG_rl_124_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_124_en )
		RG_rl_124 <= RG_rl_124_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_137 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_125_t1 = TR_137 ;
	7'h01 :
		RG_rl_125_t1 = TR_137 ;
	7'h02 :
		RG_rl_125_t1 = TR_137 ;
	7'h03 :
		RG_rl_125_t1 = TR_137 ;
	7'h04 :
		RG_rl_125_t1 = TR_137 ;
	7'h05 :
		RG_rl_125_t1 = TR_137 ;
	7'h06 :
		RG_rl_125_t1 = TR_137 ;
	7'h07 :
		RG_rl_125_t1 = TR_137 ;
	7'h08 :
		RG_rl_125_t1 = TR_137 ;
	7'h09 :
		RG_rl_125_t1 = TR_137 ;
	7'h0a :
		RG_rl_125_t1 = TR_137 ;
	7'h0b :
		RG_rl_125_t1 = TR_137 ;
	7'h0c :
		RG_rl_125_t1 = TR_137 ;
	7'h0d :
		RG_rl_125_t1 = TR_137 ;
	7'h0e :
		RG_rl_125_t1 = TR_137 ;
	7'h0f :
		RG_rl_125_t1 = TR_137 ;
	7'h10 :
		RG_rl_125_t1 = TR_137 ;
	7'h11 :
		RG_rl_125_t1 = TR_137 ;
	7'h12 :
		RG_rl_125_t1 = TR_137 ;
	7'h13 :
		RG_rl_125_t1 = TR_137 ;
	7'h14 :
		RG_rl_125_t1 = TR_137 ;
	7'h15 :
		RG_rl_125_t1 = TR_137 ;
	7'h16 :
		RG_rl_125_t1 = TR_137 ;
	7'h17 :
		RG_rl_125_t1 = TR_137 ;
	7'h18 :
		RG_rl_125_t1 = TR_137 ;
	7'h19 :
		RG_rl_125_t1 = TR_137 ;
	7'h1a :
		RG_rl_125_t1 = TR_137 ;
	7'h1b :
		RG_rl_125_t1 = TR_137 ;
	7'h1c :
		RG_rl_125_t1 = TR_137 ;
	7'h1d :
		RG_rl_125_t1 = TR_137 ;
	7'h1e :
		RG_rl_125_t1 = TR_137 ;
	7'h1f :
		RG_rl_125_t1 = TR_137 ;
	7'h20 :
		RG_rl_125_t1 = TR_137 ;
	7'h21 :
		RG_rl_125_t1 = TR_137 ;
	7'h22 :
		RG_rl_125_t1 = TR_137 ;
	7'h23 :
		RG_rl_125_t1 = TR_137 ;
	7'h24 :
		RG_rl_125_t1 = TR_137 ;
	7'h25 :
		RG_rl_125_t1 = TR_137 ;
	7'h26 :
		RG_rl_125_t1 = TR_137 ;
	7'h27 :
		RG_rl_125_t1 = TR_137 ;
	7'h28 :
		RG_rl_125_t1 = TR_137 ;
	7'h29 :
		RG_rl_125_t1 = TR_137 ;
	7'h2a :
		RG_rl_125_t1 = TR_137 ;
	7'h2b :
		RG_rl_125_t1 = TR_137 ;
	7'h2c :
		RG_rl_125_t1 = TR_137 ;
	7'h2d :
		RG_rl_125_t1 = TR_137 ;
	7'h2e :
		RG_rl_125_t1 = TR_137 ;
	7'h2f :
		RG_rl_125_t1 = TR_137 ;
	7'h30 :
		RG_rl_125_t1 = TR_137 ;
	7'h31 :
		RG_rl_125_t1 = TR_137 ;
	7'h32 :
		RG_rl_125_t1 = TR_137 ;
	7'h33 :
		RG_rl_125_t1 = TR_137 ;
	7'h34 :
		RG_rl_125_t1 = TR_137 ;
	7'h35 :
		RG_rl_125_t1 = TR_137 ;
	7'h36 :
		RG_rl_125_t1 = TR_137 ;
	7'h37 :
		RG_rl_125_t1 = TR_137 ;
	7'h38 :
		RG_rl_125_t1 = TR_137 ;
	7'h39 :
		RG_rl_125_t1 = TR_137 ;
	7'h3a :
		RG_rl_125_t1 = TR_137 ;
	7'h3b :
		RG_rl_125_t1 = TR_137 ;
	7'h3c :
		RG_rl_125_t1 = TR_137 ;
	7'h3d :
		RG_rl_125_t1 = TR_137 ;
	7'h3e :
		RG_rl_125_t1 = TR_137 ;
	7'h3f :
		RG_rl_125_t1 = TR_137 ;
	7'h40 :
		RG_rl_125_t1 = TR_137 ;
	7'h41 :
		RG_rl_125_t1 = TR_137 ;
	7'h42 :
		RG_rl_125_t1 = TR_137 ;
	7'h43 :
		RG_rl_125_t1 = TR_137 ;
	7'h44 :
		RG_rl_125_t1 = TR_137 ;
	7'h45 :
		RG_rl_125_t1 = TR_137 ;
	7'h46 :
		RG_rl_125_t1 = TR_137 ;
	7'h47 :
		RG_rl_125_t1 = TR_137 ;
	7'h48 :
		RG_rl_125_t1 = TR_137 ;
	7'h49 :
		RG_rl_125_t1 = TR_137 ;
	7'h4a :
		RG_rl_125_t1 = TR_137 ;
	7'h4b :
		RG_rl_125_t1 = TR_137 ;
	7'h4c :
		RG_rl_125_t1 = TR_137 ;
	7'h4d :
		RG_rl_125_t1 = TR_137 ;
	7'h4e :
		RG_rl_125_t1 = TR_137 ;
	7'h4f :
		RG_rl_125_t1 = TR_137 ;
	7'h50 :
		RG_rl_125_t1 = TR_137 ;
	7'h51 :
		RG_rl_125_t1 = TR_137 ;
	7'h52 :
		RG_rl_125_t1 = TR_137 ;
	7'h53 :
		RG_rl_125_t1 = TR_137 ;
	7'h54 :
		RG_rl_125_t1 = TR_137 ;
	7'h55 :
		RG_rl_125_t1 = TR_137 ;
	7'h56 :
		RG_rl_125_t1 = TR_137 ;
	7'h57 :
		RG_rl_125_t1 = TR_137 ;
	7'h58 :
		RG_rl_125_t1 = TR_137 ;
	7'h59 :
		RG_rl_125_t1 = TR_137 ;
	7'h5a :
		RG_rl_125_t1 = TR_137 ;
	7'h5b :
		RG_rl_125_t1 = TR_137 ;
	7'h5c :
		RG_rl_125_t1 = TR_137 ;
	7'h5d :
		RG_rl_125_t1 = TR_137 ;
	7'h5e :
		RG_rl_125_t1 = TR_137 ;
	7'h5f :
		RG_rl_125_t1 = TR_137 ;
	7'h60 :
		RG_rl_125_t1 = TR_137 ;
	7'h61 :
		RG_rl_125_t1 = TR_137 ;
	7'h62 :
		RG_rl_125_t1 = TR_137 ;
	7'h63 :
		RG_rl_125_t1 = TR_137 ;
	7'h64 :
		RG_rl_125_t1 = TR_137 ;
	7'h65 :
		RG_rl_125_t1 = TR_137 ;
	7'h66 :
		RG_rl_125_t1 = TR_137 ;
	7'h67 :
		RG_rl_125_t1 = TR_137 ;
	7'h68 :
		RG_rl_125_t1 = TR_137 ;
	7'h69 :
		RG_rl_125_t1 = TR_137 ;
	7'h6a :
		RG_rl_125_t1 = TR_137 ;
	7'h6b :
		RG_rl_125_t1 = TR_137 ;
	7'h6c :
		RG_rl_125_t1 = TR_137 ;
	7'h6d :
		RG_rl_125_t1 = TR_137 ;
	7'h6e :
		RG_rl_125_t1 = TR_137 ;
	7'h6f :
		RG_rl_125_t1 = TR_137 ;
	7'h70 :
		RG_rl_125_t1 = TR_137 ;
	7'h71 :
		RG_rl_125_t1 = TR_137 ;
	7'h72 :
		RG_rl_125_t1 = TR_137 ;
	7'h73 :
		RG_rl_125_t1 = TR_137 ;
	7'h74 :
		RG_rl_125_t1 = TR_137 ;
	7'h75 :
		RG_rl_125_t1 = TR_137 ;
	7'h76 :
		RG_rl_125_t1 = TR_137 ;
	7'h77 :
		RG_rl_125_t1 = TR_137 ;
	7'h78 :
		RG_rl_125_t1 = TR_137 ;
	7'h79 :
		RG_rl_125_t1 = TR_137 ;
	7'h7a :
		RG_rl_125_t1 = TR_137 ;
	7'h7b :
		RG_rl_125_t1 = TR_137 ;
	7'h7c :
		RG_rl_125_t1 = TR_137 ;
	7'h7d :
		RG_rl_125_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7e :
		RG_rl_125_t1 = TR_137 ;
	7'h7f :
		RG_rl_125_t1 = TR_137 ;
	default :
		RG_rl_125_t1 = 9'hx ;
	endcase
always @ ( RG_rl_125_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_61 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_125_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h7d ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_125_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_61 )
		| ( { 9{ U_569 } } & RG_rl_125_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_125_en = ( U_570 | RG_rl_125_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_125_en )
		RG_rl_125 <= RG_rl_125_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_138 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_126_t1 = TR_138 ;
	7'h01 :
		RG_rl_126_t1 = TR_138 ;
	7'h02 :
		RG_rl_126_t1 = TR_138 ;
	7'h03 :
		RG_rl_126_t1 = TR_138 ;
	7'h04 :
		RG_rl_126_t1 = TR_138 ;
	7'h05 :
		RG_rl_126_t1 = TR_138 ;
	7'h06 :
		RG_rl_126_t1 = TR_138 ;
	7'h07 :
		RG_rl_126_t1 = TR_138 ;
	7'h08 :
		RG_rl_126_t1 = TR_138 ;
	7'h09 :
		RG_rl_126_t1 = TR_138 ;
	7'h0a :
		RG_rl_126_t1 = TR_138 ;
	7'h0b :
		RG_rl_126_t1 = TR_138 ;
	7'h0c :
		RG_rl_126_t1 = TR_138 ;
	7'h0d :
		RG_rl_126_t1 = TR_138 ;
	7'h0e :
		RG_rl_126_t1 = TR_138 ;
	7'h0f :
		RG_rl_126_t1 = TR_138 ;
	7'h10 :
		RG_rl_126_t1 = TR_138 ;
	7'h11 :
		RG_rl_126_t1 = TR_138 ;
	7'h12 :
		RG_rl_126_t1 = TR_138 ;
	7'h13 :
		RG_rl_126_t1 = TR_138 ;
	7'h14 :
		RG_rl_126_t1 = TR_138 ;
	7'h15 :
		RG_rl_126_t1 = TR_138 ;
	7'h16 :
		RG_rl_126_t1 = TR_138 ;
	7'h17 :
		RG_rl_126_t1 = TR_138 ;
	7'h18 :
		RG_rl_126_t1 = TR_138 ;
	7'h19 :
		RG_rl_126_t1 = TR_138 ;
	7'h1a :
		RG_rl_126_t1 = TR_138 ;
	7'h1b :
		RG_rl_126_t1 = TR_138 ;
	7'h1c :
		RG_rl_126_t1 = TR_138 ;
	7'h1d :
		RG_rl_126_t1 = TR_138 ;
	7'h1e :
		RG_rl_126_t1 = TR_138 ;
	7'h1f :
		RG_rl_126_t1 = TR_138 ;
	7'h20 :
		RG_rl_126_t1 = TR_138 ;
	7'h21 :
		RG_rl_126_t1 = TR_138 ;
	7'h22 :
		RG_rl_126_t1 = TR_138 ;
	7'h23 :
		RG_rl_126_t1 = TR_138 ;
	7'h24 :
		RG_rl_126_t1 = TR_138 ;
	7'h25 :
		RG_rl_126_t1 = TR_138 ;
	7'h26 :
		RG_rl_126_t1 = TR_138 ;
	7'h27 :
		RG_rl_126_t1 = TR_138 ;
	7'h28 :
		RG_rl_126_t1 = TR_138 ;
	7'h29 :
		RG_rl_126_t1 = TR_138 ;
	7'h2a :
		RG_rl_126_t1 = TR_138 ;
	7'h2b :
		RG_rl_126_t1 = TR_138 ;
	7'h2c :
		RG_rl_126_t1 = TR_138 ;
	7'h2d :
		RG_rl_126_t1 = TR_138 ;
	7'h2e :
		RG_rl_126_t1 = TR_138 ;
	7'h2f :
		RG_rl_126_t1 = TR_138 ;
	7'h30 :
		RG_rl_126_t1 = TR_138 ;
	7'h31 :
		RG_rl_126_t1 = TR_138 ;
	7'h32 :
		RG_rl_126_t1 = TR_138 ;
	7'h33 :
		RG_rl_126_t1 = TR_138 ;
	7'h34 :
		RG_rl_126_t1 = TR_138 ;
	7'h35 :
		RG_rl_126_t1 = TR_138 ;
	7'h36 :
		RG_rl_126_t1 = TR_138 ;
	7'h37 :
		RG_rl_126_t1 = TR_138 ;
	7'h38 :
		RG_rl_126_t1 = TR_138 ;
	7'h39 :
		RG_rl_126_t1 = TR_138 ;
	7'h3a :
		RG_rl_126_t1 = TR_138 ;
	7'h3b :
		RG_rl_126_t1 = TR_138 ;
	7'h3c :
		RG_rl_126_t1 = TR_138 ;
	7'h3d :
		RG_rl_126_t1 = TR_138 ;
	7'h3e :
		RG_rl_126_t1 = TR_138 ;
	7'h3f :
		RG_rl_126_t1 = TR_138 ;
	7'h40 :
		RG_rl_126_t1 = TR_138 ;
	7'h41 :
		RG_rl_126_t1 = TR_138 ;
	7'h42 :
		RG_rl_126_t1 = TR_138 ;
	7'h43 :
		RG_rl_126_t1 = TR_138 ;
	7'h44 :
		RG_rl_126_t1 = TR_138 ;
	7'h45 :
		RG_rl_126_t1 = TR_138 ;
	7'h46 :
		RG_rl_126_t1 = TR_138 ;
	7'h47 :
		RG_rl_126_t1 = TR_138 ;
	7'h48 :
		RG_rl_126_t1 = TR_138 ;
	7'h49 :
		RG_rl_126_t1 = TR_138 ;
	7'h4a :
		RG_rl_126_t1 = TR_138 ;
	7'h4b :
		RG_rl_126_t1 = TR_138 ;
	7'h4c :
		RG_rl_126_t1 = TR_138 ;
	7'h4d :
		RG_rl_126_t1 = TR_138 ;
	7'h4e :
		RG_rl_126_t1 = TR_138 ;
	7'h4f :
		RG_rl_126_t1 = TR_138 ;
	7'h50 :
		RG_rl_126_t1 = TR_138 ;
	7'h51 :
		RG_rl_126_t1 = TR_138 ;
	7'h52 :
		RG_rl_126_t1 = TR_138 ;
	7'h53 :
		RG_rl_126_t1 = TR_138 ;
	7'h54 :
		RG_rl_126_t1 = TR_138 ;
	7'h55 :
		RG_rl_126_t1 = TR_138 ;
	7'h56 :
		RG_rl_126_t1 = TR_138 ;
	7'h57 :
		RG_rl_126_t1 = TR_138 ;
	7'h58 :
		RG_rl_126_t1 = TR_138 ;
	7'h59 :
		RG_rl_126_t1 = TR_138 ;
	7'h5a :
		RG_rl_126_t1 = TR_138 ;
	7'h5b :
		RG_rl_126_t1 = TR_138 ;
	7'h5c :
		RG_rl_126_t1 = TR_138 ;
	7'h5d :
		RG_rl_126_t1 = TR_138 ;
	7'h5e :
		RG_rl_126_t1 = TR_138 ;
	7'h5f :
		RG_rl_126_t1 = TR_138 ;
	7'h60 :
		RG_rl_126_t1 = TR_138 ;
	7'h61 :
		RG_rl_126_t1 = TR_138 ;
	7'h62 :
		RG_rl_126_t1 = TR_138 ;
	7'h63 :
		RG_rl_126_t1 = TR_138 ;
	7'h64 :
		RG_rl_126_t1 = TR_138 ;
	7'h65 :
		RG_rl_126_t1 = TR_138 ;
	7'h66 :
		RG_rl_126_t1 = TR_138 ;
	7'h67 :
		RG_rl_126_t1 = TR_138 ;
	7'h68 :
		RG_rl_126_t1 = TR_138 ;
	7'h69 :
		RG_rl_126_t1 = TR_138 ;
	7'h6a :
		RG_rl_126_t1 = TR_138 ;
	7'h6b :
		RG_rl_126_t1 = TR_138 ;
	7'h6c :
		RG_rl_126_t1 = TR_138 ;
	7'h6d :
		RG_rl_126_t1 = TR_138 ;
	7'h6e :
		RG_rl_126_t1 = TR_138 ;
	7'h6f :
		RG_rl_126_t1 = TR_138 ;
	7'h70 :
		RG_rl_126_t1 = TR_138 ;
	7'h71 :
		RG_rl_126_t1 = TR_138 ;
	7'h72 :
		RG_rl_126_t1 = TR_138 ;
	7'h73 :
		RG_rl_126_t1 = TR_138 ;
	7'h74 :
		RG_rl_126_t1 = TR_138 ;
	7'h75 :
		RG_rl_126_t1 = TR_138 ;
	7'h76 :
		RG_rl_126_t1 = TR_138 ;
	7'h77 :
		RG_rl_126_t1 = TR_138 ;
	7'h78 :
		RG_rl_126_t1 = TR_138 ;
	7'h79 :
		RG_rl_126_t1 = TR_138 ;
	7'h7a :
		RG_rl_126_t1 = TR_138 ;
	7'h7b :
		RG_rl_126_t1 = TR_138 ;
	7'h7c :
		RG_rl_126_t1 = TR_138 ;
	7'h7d :
		RG_rl_126_t1 = TR_138 ;
	7'h7e :
		RG_rl_126_t1 = 9'h000 ;	// line#=../rle.cpp:80
	7'h7f :
		RG_rl_126_t1 = TR_138 ;
	default :
		RG_rl_126_t1 = 9'hx ;
	endcase
always @ ( RG_rl_126_t1 or U_569 or sub8u_71ot or U_571 or RG_previous_dc_rl_1 or 
	M_318 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_126_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h7e ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_126_t = ( ( { 9{ M_318 } } & RG_previous_dc_rl_1 )
		| ( { 9{ U_569 } } & RG_rl_126_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_126_en = ( M_318 | RG_rl_126_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_126_en )
		RG_rl_126 <= RG_rl_126_t ;	// line#=../rle.cpp:79,80,83,84,85
always @ ( TR_11 or incr8u1ot )	// line#=../rle.cpp:79,80
	case ( incr8u1ot [6:0] )
	7'h00 :
		RG_rl_127_t1 = TR_11 ;
	7'h01 :
		RG_rl_127_t1 = TR_11 ;
	7'h02 :
		RG_rl_127_t1 = TR_11 ;
	7'h03 :
		RG_rl_127_t1 = TR_11 ;
	7'h04 :
		RG_rl_127_t1 = TR_11 ;
	7'h05 :
		RG_rl_127_t1 = TR_11 ;
	7'h06 :
		RG_rl_127_t1 = TR_11 ;
	7'h07 :
		RG_rl_127_t1 = TR_11 ;
	7'h08 :
		RG_rl_127_t1 = TR_11 ;
	7'h09 :
		RG_rl_127_t1 = TR_11 ;
	7'h0a :
		RG_rl_127_t1 = TR_11 ;
	7'h0b :
		RG_rl_127_t1 = TR_11 ;
	7'h0c :
		RG_rl_127_t1 = TR_11 ;
	7'h0d :
		RG_rl_127_t1 = TR_11 ;
	7'h0e :
		RG_rl_127_t1 = TR_11 ;
	7'h0f :
		RG_rl_127_t1 = TR_11 ;
	7'h10 :
		RG_rl_127_t1 = TR_11 ;
	7'h11 :
		RG_rl_127_t1 = TR_11 ;
	7'h12 :
		RG_rl_127_t1 = TR_11 ;
	7'h13 :
		RG_rl_127_t1 = TR_11 ;
	7'h14 :
		RG_rl_127_t1 = TR_11 ;
	7'h15 :
		RG_rl_127_t1 = TR_11 ;
	7'h16 :
		RG_rl_127_t1 = TR_11 ;
	7'h17 :
		RG_rl_127_t1 = TR_11 ;
	7'h18 :
		RG_rl_127_t1 = TR_11 ;
	7'h19 :
		RG_rl_127_t1 = TR_11 ;
	7'h1a :
		RG_rl_127_t1 = TR_11 ;
	7'h1b :
		RG_rl_127_t1 = TR_11 ;
	7'h1c :
		RG_rl_127_t1 = TR_11 ;
	7'h1d :
		RG_rl_127_t1 = TR_11 ;
	7'h1e :
		RG_rl_127_t1 = TR_11 ;
	7'h1f :
		RG_rl_127_t1 = TR_11 ;
	7'h20 :
		RG_rl_127_t1 = TR_11 ;
	7'h21 :
		RG_rl_127_t1 = TR_11 ;
	7'h22 :
		RG_rl_127_t1 = TR_11 ;
	7'h23 :
		RG_rl_127_t1 = TR_11 ;
	7'h24 :
		RG_rl_127_t1 = TR_11 ;
	7'h25 :
		RG_rl_127_t1 = TR_11 ;
	7'h26 :
		RG_rl_127_t1 = TR_11 ;
	7'h27 :
		RG_rl_127_t1 = TR_11 ;
	7'h28 :
		RG_rl_127_t1 = TR_11 ;
	7'h29 :
		RG_rl_127_t1 = TR_11 ;
	7'h2a :
		RG_rl_127_t1 = TR_11 ;
	7'h2b :
		RG_rl_127_t1 = TR_11 ;
	7'h2c :
		RG_rl_127_t1 = TR_11 ;
	7'h2d :
		RG_rl_127_t1 = TR_11 ;
	7'h2e :
		RG_rl_127_t1 = TR_11 ;
	7'h2f :
		RG_rl_127_t1 = TR_11 ;
	7'h30 :
		RG_rl_127_t1 = TR_11 ;
	7'h31 :
		RG_rl_127_t1 = TR_11 ;
	7'h32 :
		RG_rl_127_t1 = TR_11 ;
	7'h33 :
		RG_rl_127_t1 = TR_11 ;
	7'h34 :
		RG_rl_127_t1 = TR_11 ;
	7'h35 :
		RG_rl_127_t1 = TR_11 ;
	7'h36 :
		RG_rl_127_t1 = TR_11 ;
	7'h37 :
		RG_rl_127_t1 = TR_11 ;
	7'h38 :
		RG_rl_127_t1 = TR_11 ;
	7'h39 :
		RG_rl_127_t1 = TR_11 ;
	7'h3a :
		RG_rl_127_t1 = TR_11 ;
	7'h3b :
		RG_rl_127_t1 = TR_11 ;
	7'h3c :
		RG_rl_127_t1 = TR_11 ;
	7'h3d :
		RG_rl_127_t1 = TR_11 ;
	7'h3e :
		RG_rl_127_t1 = TR_11 ;
	7'h3f :
		RG_rl_127_t1 = TR_11 ;
	7'h40 :
		RG_rl_127_t1 = TR_11 ;
	7'h41 :
		RG_rl_127_t1 = TR_11 ;
	7'h42 :
		RG_rl_127_t1 = TR_11 ;
	7'h43 :
		RG_rl_127_t1 = TR_11 ;
	7'h44 :
		RG_rl_127_t1 = TR_11 ;
	7'h45 :
		RG_rl_127_t1 = TR_11 ;
	7'h46 :
		RG_rl_127_t1 = TR_11 ;
	7'h47 :
		RG_rl_127_t1 = TR_11 ;
	7'h48 :
		RG_rl_127_t1 = TR_11 ;
	7'h49 :
		RG_rl_127_t1 = TR_11 ;
	7'h4a :
		RG_rl_127_t1 = TR_11 ;
	7'h4b :
		RG_rl_127_t1 = TR_11 ;
	7'h4c :
		RG_rl_127_t1 = TR_11 ;
	7'h4d :
		RG_rl_127_t1 = TR_11 ;
	7'h4e :
		RG_rl_127_t1 = TR_11 ;
	7'h4f :
		RG_rl_127_t1 = TR_11 ;
	7'h50 :
		RG_rl_127_t1 = TR_11 ;
	7'h51 :
		RG_rl_127_t1 = TR_11 ;
	7'h52 :
		RG_rl_127_t1 = TR_11 ;
	7'h53 :
		RG_rl_127_t1 = TR_11 ;
	7'h54 :
		RG_rl_127_t1 = TR_11 ;
	7'h55 :
		RG_rl_127_t1 = TR_11 ;
	7'h56 :
		RG_rl_127_t1 = TR_11 ;
	7'h57 :
		RG_rl_127_t1 = TR_11 ;
	7'h58 :
		RG_rl_127_t1 = TR_11 ;
	7'h59 :
		RG_rl_127_t1 = TR_11 ;
	7'h5a :
		RG_rl_127_t1 = TR_11 ;
	7'h5b :
		RG_rl_127_t1 = TR_11 ;
	7'h5c :
		RG_rl_127_t1 = TR_11 ;
	7'h5d :
		RG_rl_127_t1 = TR_11 ;
	7'h5e :
		RG_rl_127_t1 = TR_11 ;
	7'h5f :
		RG_rl_127_t1 = TR_11 ;
	7'h60 :
		RG_rl_127_t1 = TR_11 ;
	7'h61 :
		RG_rl_127_t1 = TR_11 ;
	7'h62 :
		RG_rl_127_t1 = TR_11 ;
	7'h63 :
		RG_rl_127_t1 = TR_11 ;
	7'h64 :
		RG_rl_127_t1 = TR_11 ;
	7'h65 :
		RG_rl_127_t1 = TR_11 ;
	7'h66 :
		RG_rl_127_t1 = TR_11 ;
	7'h67 :
		RG_rl_127_t1 = TR_11 ;
	7'h68 :
		RG_rl_127_t1 = TR_11 ;
	7'h69 :
		RG_rl_127_t1 = TR_11 ;
	7'h6a :
		RG_rl_127_t1 = TR_11 ;
	7'h6b :
		RG_rl_127_t1 = TR_11 ;
	7'h6c :
		RG_rl_127_t1 = TR_11 ;
	7'h6d :
		RG_rl_127_t1 = TR_11 ;
	7'h6e :
		RG_rl_127_t1 = TR_11 ;
	7'h6f :
		RG_rl_127_t1 = TR_11 ;
	7'h70 :
		RG_rl_127_t1 = TR_11 ;
	7'h71 :
		RG_rl_127_t1 = TR_11 ;
	7'h72 :
		RG_rl_127_t1 = TR_11 ;
	7'h73 :
		RG_rl_127_t1 = TR_11 ;
	7'h74 :
		RG_rl_127_t1 = TR_11 ;
	7'h75 :
		RG_rl_127_t1 = TR_11 ;
	7'h76 :
		RG_rl_127_t1 = TR_11 ;
	7'h77 :
		RG_rl_127_t1 = TR_11 ;
	7'h78 :
		RG_rl_127_t1 = TR_11 ;
	7'h79 :
		RG_rl_127_t1 = TR_11 ;
	7'h7a :
		RG_rl_127_t1 = TR_11 ;
	7'h7b :
		RG_rl_127_t1 = TR_11 ;
	7'h7c :
		RG_rl_127_t1 = TR_11 ;
	7'h7d :
		RG_rl_127_t1 = TR_11 ;
	7'h7e :
		RG_rl_127_t1 = TR_11 ;
	7'h7f :
		RG_rl_127_t1 = 9'h000 ;	// line#=../rle.cpp:80
	default :
		RG_rl_127_t1 = 9'hx ;
	endcase
always @ ( RG_rl_127_t1 or U_569 or sub8u_71ot or U_571 or RG_quantized_block_rl_62 or 
	U_570 )	// line#=../rle.cpp:83,84,85
	begin
	RG_rl_127_t_c1 = ( U_571 & ( ~|( sub8u_71ot ^ 7'h7f ) ) ) ;	// line#=../rle.cpp:85
	RG_rl_127_t = ( ( { 9{ U_570 } } & RG_quantized_block_rl_62 )
		| ( { 9{ U_569 } } & RG_rl_127_t1 )	// line#=../rle.cpp:79,80
		) ;	// line#=../rle.cpp:85
	end
assign	RG_rl_127_en = ( U_570 | RG_rl_127_t_c1 | U_569 ) ;	// line#=../rle.cpp:83,84,85
always @ ( posedge clk )	// line#=../rle.cpp:83,84,85
	if ( RG_rl_127_en )
		RG_rl_127 <= RG_rl_127_t ;	// line#=../rle.cpp:79,80,83,84,85
assign	RG_previous_dc_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_previous_dc_en )
		RG_previous_dc <= RG_previous_dc_rl_1 ;
assign	RG_rl_128_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_128_en )
		RG_rl_128 <= RG_rl_185 ;
assign	RG_rl_129_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_129_en )
		RG_rl_129 <= RG_rl_186 ;
assign	RG_rl_130_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_130_en )
		RG_rl_130 <= RG_rl_187 ;
assign	RG_rl_131_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_131_en )
		RG_rl_131 <= RG_rl_188 ;
assign	RG_rl_132_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_132_en )
		RG_rl_132 <= RG_rl_189 ;
assign	RG_rl_133_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_133_en )
		RG_rl_133 <= RG_rl_190 ;
assign	RG_rl_134_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_134_en )
		RG_rl_134 <= RG_rl_191 ;
assign	RG_rl_135_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_135_en )
		RG_rl_135 <= RG_rl_192 ;
assign	RG_rl_136_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_136_en )
		RG_rl_136 <= RG_rl_193 ;
assign	RG_rl_137_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_137_en )
		RG_rl_137 <= RG_rl_194 ;
assign	RG_rl_138_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_138_en )
		RG_rl_138 <= RG_rl_195 ;
assign	RG_rl_139_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_139_en )
		RG_rl_139 <= RG_rl_196 ;
assign	RG_rl_140_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_140_en )
		RG_rl_140 <= RG_rl_197 ;
assign	RG_rl_141_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_141_en )
		RG_rl_141 <= RG_rl_198 ;
assign	RG_rl_142_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_142_en )
		RG_rl_142 <= RG_rl_199 ;
assign	RG_rl_143_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_143_en )
		RG_rl_143 <= RG_rl_200 ;
assign	RG_rl_144_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_144_en )
		RG_rl_144 <= RG_rl_201 ;
assign	RG_rl_145_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_145_en )
		RG_rl_145 <= RG_rl_202 ;
assign	RG_rl_146_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_146_en )
		RG_rl_146 <= RG_rl_203 ;
assign	RG_rl_147_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_147_en )
		RG_rl_147 <= RG_rl_204 ;
assign	RG_rl_148_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_148_en )
		RG_rl_148 <= RG_rl_205 ;
assign	RG_rl_149_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_149_en )
		RG_rl_149 <= RG_rl_206 ;
assign	RG_rl_150_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_150_en )
		RG_rl_150 <= RG_rl_207 ;
assign	RG_rl_151_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_151_en )
		RG_rl_151 <= RG_rl_208 ;
assign	RG_rl_152_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_152_en )
		RG_rl_152 <= RG_rl_209 ;
assign	RG_rl_153_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_153_en )
		RG_rl_153 <= RG_rl_210 ;
assign	RG_rl_154_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_154_en )
		RG_rl_154 <= RG_rl_211 ;
assign	RG_rl_155_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_155_en )
		RG_rl_155 <= RG_rl_212 ;
assign	RG_rl_156_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_156_en )
		RG_rl_156 <= RG_rl_213 ;
assign	RG_rl_157_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_157_en )
		RG_rl_157 <= RG_rl_214 ;
assign	RG_rl_158_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_158_en )
		RG_rl_158 <= RG_rl_215 ;
assign	RG_rl_159_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_159_en )
		RG_rl_159 <= RG_rl_216 ;
assign	RG_rl_160_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_160_en )
		RG_rl_160 <= RG_rl_217 ;
assign	RG_rl_161_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_161_en )
		RG_rl_161 <= RG_rl_218 ;
assign	RG_rl_162_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_162_en )
		RG_rl_162 <= RG_rl_219 ;
assign	RG_rl_163_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_163_en )
		RG_rl_163 <= RG_rl_220 ;
assign	RG_rl_164_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_164_en )
		RG_rl_164 <= RG_rl_221 ;
assign	RG_rl_165_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_165_en )
		RG_rl_165 <= RG_rl_222 ;
assign	RG_rl_166_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_166_en )
		RG_rl_166 <= RG_rl_223 ;
assign	RG_rl_167_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_167_en )
		RG_rl_167 <= RG_rl_224 ;
assign	RG_rl_168_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_168_en )
		RG_rl_168 <= RG_rl_225 ;
assign	RG_rl_169_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_169_en )
		RG_rl_169 <= RG_rl_226 ;
assign	RG_rl_170_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_170_en )
		RG_rl_170 <= RG_rl_227 ;
assign	RG_rl_171_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_171_en )
		RG_rl_171 <= RG_rl_228 ;
assign	RG_rl_172_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_172_en )
		RG_rl_172 <= RG_rl_229 ;
assign	RG_rl_173_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_173_en )
		RG_rl_173 <= RG_rl_230 ;
assign	RG_rl_174_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_174_en )
		RG_rl_174 <= RG_rl_231 ;
assign	RG_rl_175_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_175_en )
		RG_rl_175 <= RG_rl_232 ;
assign	RG_rl_176_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_176_en )
		RG_rl_176 <= RG_rl_233 ;
assign	RG_rl_177_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_177_en )
		RG_rl_177 <= RG_rl_234 ;
assign	RG_rl_178_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_178_en )
		RG_rl_178 <= RG_rl_235 ;
assign	RG_rl_179_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_179_en )
		RG_rl_179 <= RG_rl_236 ;
assign	RG_rl_180_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_180_en )
		RG_rl_180 <= RG_rl_237 ;
assign	RG_rl_181_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_181_en )
		RG_rl_181 <= RG_rl_238 ;
assign	RG_rl_182_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_182_en )
		RG_rl_182 <= RG_rl_239 ;
assign	RG_rl_183_en = ST1_02d ;
always @ ( posedge clk )
	if ( RG_rl_183_en )
		RG_rl_183 <= RG_rl_240 ;
always @ ( rl_a00_t4 or ST1_09d or RG_i_k_01 or RG_len or U_174 or sub12s_91ot or 
	ST1_06d or RG_rl_241 or ST1_02d )	// line#=../rle.cpp:73
	begin
	RG_rl_184_t_c1 = ( U_174 & ( ~|RG_len [6:0] ) ) ;	// line#=../rle.cpp:73
	RG_rl_184_t = ( ( { 9{ ST1_02d } } & RG_rl_241 )
		| ( { 9{ ST1_06d } } & sub12s_91ot )		// line#=../rle.cpp:52
		| ( { 9{ RG_rl_184_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a00_t4 ) ) ;
	end
assign	RG_rl_184_en = ( ST1_02d | ST1_06d | RG_rl_184_t_c1 | ST1_09d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_184_en )
		RG_rl_184 <= RG_rl_184_t ;	// line#=../rle.cpp:52,73
always @ ( rl_a01_t4 or ST1_09d or RG_i_k_01 or RG_len or U_174 or RG_rl_185 or 
	ST1_06d or RG_previous_dc or ST1_05d or RG_quantized_block_rl or ST1_02d )	// line#=../rle.cpp:73
	begin
	RG_previous_dc_rl_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h01 ) ) ) ;	// line#=../rle.cpp:73
	RG_previous_dc_rl_t = ( ( { 9{ ST1_02d } } & RG_quantized_block_rl )
		| ( { 9{ ST1_05d } } & RG_previous_dc )
		| ( { 9{ ST1_06d } } & RG_rl_185 )
		| ( { 9{ RG_previous_dc_rl_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a01_t4 ) ) ;
	end
assign	RG_previous_dc_rl_en = ( ST1_02d | ST1_05d | ST1_06d | RG_previous_dc_rl_t_c1 | 
	ST1_09d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( !rst )
		RG_previous_dc_rl <= 9'h000 ;
	else if ( RG_previous_dc_rl_en )
		RG_previous_dc_rl <= RG_previous_dc_rl_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_1 or ST1_11d or rl_a02_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_186 or ST1_06d or RG_rl_128 or ST1_05d or RG_quantized_block_rl_1 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_185_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h02 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_185_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_1 )
		| ( { 9{ ST1_05d } } & RG_rl_128 )
		| ( { 9{ ST1_06d } } & RG_rl_186 )
		| ( { 9{ RG_rl_185_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a02_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_1 ) ) ;
	end
assign	RG_rl_185_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_185_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_185_en )
		RG_rl_185 <= RG_rl_185_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_2 or ST1_11d or rl_a03_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_187 or ST1_06d or RG_rl_129 or ST1_05d or RG_quantized_block_rl_2 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_186_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h03 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_186_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_2 )
		| ( { 9{ ST1_05d } } & RG_rl_129 )
		| ( { 9{ ST1_06d } } & RG_rl_187 )
		| ( { 9{ RG_rl_186_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a03_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_2 ) ) ;
	end
assign	RG_rl_186_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_186_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_186_en )
		RG_rl_186 <= RG_rl_186_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_3 or ST1_11d or rl_a04_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_188 or ST1_06d or RG_rl_130 or ST1_05d or RG_quantized_block_rl_3 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_187_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h04 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_187_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_3 )
		| ( { 9{ ST1_05d } } & RG_rl_130 )
		| ( { 9{ ST1_06d } } & RG_rl_188 )
		| ( { 9{ RG_rl_187_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a04_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_3 ) ) ;
	end
assign	RG_rl_187_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_187_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_187_en )
		RG_rl_187 <= RG_rl_187_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_4 or ST1_11d or rl_a05_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_189 or ST1_06d or RG_rl_131 or ST1_05d or RG_quantized_block_rl_4 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_188_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h05 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_188_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_4 )
		| ( { 9{ ST1_05d } } & RG_rl_131 )
		| ( { 9{ ST1_06d } } & RG_rl_189 )
		| ( { 9{ RG_rl_188_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a05_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_4 ) ) ;
	end
assign	RG_rl_188_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_188_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_188_en )
		RG_rl_188 <= RG_rl_188_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_5 or ST1_11d or rl_a06_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_190 or ST1_06d or RG_rl_132 or ST1_05d or RG_quantized_block_rl_5 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_189_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h06 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_189_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_5 )
		| ( { 9{ ST1_05d } } & RG_rl_132 )
		| ( { 9{ ST1_06d } } & RG_rl_190 )
		| ( { 9{ RG_rl_189_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a06_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_5 ) ) ;
	end
assign	RG_rl_189_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_189_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_189_en )
		RG_rl_189 <= RG_rl_189_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_6 or ST1_11d or rl_a07_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_191 or ST1_06d or RG_rl_133 or ST1_05d or RG_quantized_block_rl_6 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_190_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h07 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_190_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_6 )
		| ( { 9{ ST1_05d } } & RG_rl_133 )
		| ( { 9{ ST1_06d } } & RG_rl_191 )
		| ( { 9{ RG_rl_190_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a07_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_6 ) ) ;
	end
assign	RG_rl_190_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_190_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_190_en )
		RG_rl_190 <= RG_rl_190_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_7 or ST1_11d or rl_a08_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_192 or ST1_06d or RG_rl_134 or ST1_05d or RG_quantized_block_rl_7 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_191_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h08 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_191_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_7 )
		| ( { 9{ ST1_05d } } & RG_rl_134 )
		| ( { 9{ ST1_06d } } & RG_rl_192 )
		| ( { 9{ RG_rl_191_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a08_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_7 ) ) ;
	end
assign	RG_rl_191_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_191_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_191_en )
		RG_rl_191 <= RG_rl_191_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_8 or ST1_11d or rl_a09_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_193 or ST1_06d or RG_rl_135 or ST1_05d or RG_quantized_block_rl_8 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_192_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h09 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_192_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_8 )
		| ( { 9{ ST1_05d } } & RG_rl_135 )
		| ( { 9{ ST1_06d } } & RG_rl_193 )
		| ( { 9{ RG_rl_192_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a09_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_8 ) ) ;
	end
assign	RG_rl_192_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_192_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_192_en )
		RG_rl_192 <= RG_rl_192_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_9 or ST1_11d or rl_a10_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_194 or ST1_06d or RG_rl_136 or ST1_05d or RG_quantized_block_rl_9 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_193_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h0a ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_193_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_9 )
		| ( { 9{ ST1_05d } } & RG_rl_136 )
		| ( { 9{ ST1_06d } } & RG_rl_194 )
		| ( { 9{ RG_rl_193_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a10_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_9 ) ) ;
	end
assign	RG_rl_193_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_193_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_193_en )
		RG_rl_193 <= RG_rl_193_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_10 or ST1_11d or rl_a11_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_195 or ST1_06d or RG_rl_137 or ST1_05d or RG_quantized_block_rl_10 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_194_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h0b ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_194_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_10 )
		| ( { 9{ ST1_05d } } & RG_rl_137 )
		| ( { 9{ ST1_06d } } & RG_rl_195 )
		| ( { 9{ RG_rl_194_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a11_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_10 ) ) ;
	end
assign	RG_rl_194_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_194_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_194_en )
		RG_rl_194 <= RG_rl_194_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_11 or ST1_11d or rl_a12_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_196 or ST1_06d or RG_rl_138 or ST1_05d or RG_quantized_block_rl_11 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_195_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h0c ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_195_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_11 )
		| ( { 9{ ST1_05d } } & RG_rl_138 )
		| ( { 9{ ST1_06d } } & RG_rl_196 )
		| ( { 9{ RG_rl_195_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a12_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_11 ) ) ;
	end
assign	RG_rl_195_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_195_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_195_en )
		RG_rl_195 <= RG_rl_195_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_12 or ST1_11d or rl_a13_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_197 or ST1_06d or RG_rl_139 or ST1_05d or RG_quantized_block_rl_12 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_196_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h0d ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_196_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_12 )
		| ( { 9{ ST1_05d } } & RG_rl_139 )
		| ( { 9{ ST1_06d } } & RG_rl_197 )
		| ( { 9{ RG_rl_196_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a13_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_12 ) ) ;
	end
assign	RG_rl_196_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_196_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_196_en )
		RG_rl_196 <= RG_rl_196_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_13 or ST1_11d or rl_a14_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_198 or ST1_06d or RG_rl_140 or ST1_05d or RG_quantized_block_rl_13 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_197_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h0e ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_197_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_13 )
		| ( { 9{ ST1_05d } } & RG_rl_140 )
		| ( { 9{ ST1_06d } } & RG_rl_198 )
		| ( { 9{ RG_rl_197_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a14_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_13 ) ) ;
	end
assign	RG_rl_197_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_197_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_197_en )
		RG_rl_197 <= RG_rl_197_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_14 or ST1_11d or rl_a15_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_199 or ST1_06d or RG_rl_141 or ST1_05d or RG_quantized_block_rl_14 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_198_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h0f ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_198_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_14 )
		| ( { 9{ ST1_05d } } & RG_rl_141 )
		| ( { 9{ ST1_06d } } & RG_rl_199 )
		| ( { 9{ RG_rl_198_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a15_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_14 ) ) ;
	end
assign	RG_rl_198_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_198_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_198_en )
		RG_rl_198 <= RG_rl_198_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_15 or ST1_11d or rl_a16_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_200 or ST1_06d or RG_rl_142 or ST1_05d or RG_quantized_block_rl_15 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_199_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h10 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_199_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_15 )
		| ( { 9{ ST1_05d } } & RG_rl_142 )
		| ( { 9{ ST1_06d } } & RG_rl_200 )
		| ( { 9{ RG_rl_199_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a16_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_15 ) ) ;
	end
assign	RG_rl_199_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_199_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_199_en )
		RG_rl_199 <= RG_rl_199_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_16 or ST1_11d or rl_a17_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_201 or ST1_06d or RG_rl_143 or ST1_05d or RG_quantized_block_rl_16 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_200_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h11 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_200_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_16 )
		| ( { 9{ ST1_05d } } & RG_rl_143 )
		| ( { 9{ ST1_06d } } & RG_rl_201 )
		| ( { 9{ RG_rl_200_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a17_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_16 ) ) ;
	end
assign	RG_rl_200_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_200_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_200_en )
		RG_rl_200 <= RG_rl_200_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_17 or ST1_11d or rl_a18_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_202 or ST1_06d or RG_rl_144 or ST1_05d or RG_quantized_block_rl_17 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_201_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h12 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_201_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_17 )
		| ( { 9{ ST1_05d } } & RG_rl_144 )
		| ( { 9{ ST1_06d } } & RG_rl_202 )
		| ( { 9{ RG_rl_201_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a18_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_17 ) ) ;
	end
assign	RG_rl_201_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_201_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_201_en )
		RG_rl_201 <= RG_rl_201_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_18 or ST1_11d or rl_a19_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_203 or ST1_06d or RG_rl_145 or ST1_05d or RG_quantized_block_rl_18 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_202_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h13 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_202_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_18 )
		| ( { 9{ ST1_05d } } & RG_rl_145 )
		| ( { 9{ ST1_06d } } & RG_rl_203 )
		| ( { 9{ RG_rl_202_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a19_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_18 ) ) ;
	end
assign	RG_rl_202_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_202_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_202_en )
		RG_rl_202 <= RG_rl_202_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_19 or ST1_11d or rl_a20_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_204 or ST1_06d or RG_rl_146 or ST1_05d or RG_quantized_block_rl_19 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_203_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h14 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_203_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_19 )
		| ( { 9{ ST1_05d } } & RG_rl_146 )
		| ( { 9{ ST1_06d } } & RG_rl_204 )
		| ( { 9{ RG_rl_203_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a20_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_19 ) ) ;
	end
assign	RG_rl_203_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_203_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_203_en )
		RG_rl_203 <= RG_rl_203_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_20 or ST1_11d or rl_a21_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_205 or ST1_06d or RG_rl_147 or ST1_05d or RG_quantized_block_rl_20 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_204_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h15 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_204_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_20 )
		| ( { 9{ ST1_05d } } & RG_rl_147 )
		| ( { 9{ ST1_06d } } & RG_rl_205 )
		| ( { 9{ RG_rl_204_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a21_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_20 ) ) ;
	end
assign	RG_rl_204_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_204_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_204_en )
		RG_rl_204 <= RG_rl_204_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_21 or ST1_11d or rl_a22_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_206 or ST1_06d or RG_rl_148 or ST1_05d or RG_quantized_block_rl_21 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_205_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h16 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_205_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_21 )
		| ( { 9{ ST1_05d } } & RG_rl_148 )
		| ( { 9{ ST1_06d } } & RG_rl_206 )
		| ( { 9{ RG_rl_205_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a22_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_21 ) ) ;
	end
assign	RG_rl_205_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_205_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_205_en )
		RG_rl_205 <= RG_rl_205_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_22 or ST1_11d or rl_a23_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_207 or ST1_06d or RG_rl_149 or ST1_05d or RG_quantized_block_rl_22 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_206_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h17 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_206_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_22 )
		| ( { 9{ ST1_05d } } & RG_rl_149 )
		| ( { 9{ ST1_06d } } & RG_rl_207 )
		| ( { 9{ RG_rl_206_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a23_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_22 ) ) ;
	end
assign	RG_rl_206_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_206_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_206_en )
		RG_rl_206 <= RG_rl_206_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_23 or ST1_11d or rl_a24_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_208 or ST1_06d or RG_rl_150 or ST1_05d or RG_quantized_block_rl_23 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_207_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h18 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_207_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_23 )
		| ( { 9{ ST1_05d } } & RG_rl_150 )
		| ( { 9{ ST1_06d } } & RG_rl_208 )
		| ( { 9{ RG_rl_207_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a24_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_23 ) ) ;
	end
assign	RG_rl_207_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_207_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_207_en )
		RG_rl_207 <= RG_rl_207_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_24 or ST1_11d or rl_a25_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_209 or ST1_06d or RG_rl_151 or ST1_05d or RG_quantized_block_rl_24 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_208_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h19 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_208_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_24 )
		| ( { 9{ ST1_05d } } & RG_rl_151 )
		| ( { 9{ ST1_06d } } & RG_rl_209 )
		| ( { 9{ RG_rl_208_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a25_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_24 ) ) ;
	end
assign	RG_rl_208_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_208_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_208_en )
		RG_rl_208 <= RG_rl_208_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_25 or ST1_11d or rl_a26_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_210 or ST1_06d or RG_rl_152 or ST1_05d or RG_quantized_block_rl_25 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_209_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h1a ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_209_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_25 )
		| ( { 9{ ST1_05d } } & RG_rl_152 )
		| ( { 9{ ST1_06d } } & RG_rl_210 )
		| ( { 9{ RG_rl_209_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a26_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_25 ) ) ;
	end
assign	RG_rl_209_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_209_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_209_en )
		RG_rl_209 <= RG_rl_209_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_26 or ST1_11d or rl_a27_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_211 or ST1_06d or RG_rl_153 or ST1_05d or RG_quantized_block_rl_26 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_210_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h1b ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_210_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_26 )
		| ( { 9{ ST1_05d } } & RG_rl_153 )
		| ( { 9{ ST1_06d } } & RG_rl_211 )
		| ( { 9{ RG_rl_210_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a27_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_26 ) ) ;
	end
assign	RG_rl_210_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_210_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_210_en )
		RG_rl_210 <= RG_rl_210_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_27 or ST1_11d or rl_a28_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_212 or ST1_06d or RG_rl_154 or ST1_05d or RG_quantized_block_rl_27 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_211_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h1c ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_211_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_27 )
		| ( { 9{ ST1_05d } } & RG_rl_154 )
		| ( { 9{ ST1_06d } } & RG_rl_212 )
		| ( { 9{ RG_rl_211_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a28_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_27 ) ) ;
	end
assign	RG_rl_211_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_211_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_211_en )
		RG_rl_211 <= RG_rl_211_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_28 or ST1_11d or rl_a29_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_213 or ST1_06d or RG_rl_155 or ST1_05d or RG_quantized_block_rl_28 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_212_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h1d ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_212_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_28 )
		| ( { 9{ ST1_05d } } & RG_rl_155 )
		| ( { 9{ ST1_06d } } & RG_rl_213 )
		| ( { 9{ RG_rl_212_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a29_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_28 ) ) ;
	end
assign	RG_rl_212_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_212_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_212_en )
		RG_rl_212 <= RG_rl_212_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_29 or ST1_11d or rl_a30_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_214 or ST1_06d or RG_rl_156 or ST1_05d or RG_quantized_block_rl_29 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_213_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h1e ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_213_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_29 )
		| ( { 9{ ST1_05d } } & RG_rl_156 )
		| ( { 9{ ST1_06d } } & RG_rl_214 )
		| ( { 9{ RG_rl_213_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a30_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_29 ) ) ;
	end
assign	RG_rl_213_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_213_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_213_en )
		RG_rl_213 <= RG_rl_213_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_30 or ST1_11d or rl_a31_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_215 or ST1_06d or RG_rl_157 or ST1_05d or RG_quantized_block_rl_30 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_214_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h1f ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_214_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_30 )
		| ( { 9{ ST1_05d } } & RG_rl_157 )
		| ( { 9{ ST1_06d } } & RG_rl_215 )
		| ( { 9{ RG_rl_214_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a31_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_30 ) ) ;
	end
assign	RG_rl_214_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_214_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_214_en )
		RG_rl_214 <= RG_rl_214_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_31 or ST1_11d or rl_a32_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_216 or ST1_06d or RG_rl_158 or ST1_05d or RG_quantized_block_rl_31 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_215_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h20 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_215_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_31 )
		| ( { 9{ ST1_05d } } & RG_rl_158 )
		| ( { 9{ ST1_06d } } & RG_rl_216 )
		| ( { 9{ RG_rl_215_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a32_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_31 ) ) ;
	end
assign	RG_rl_215_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_215_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_215_en )
		RG_rl_215 <= RG_rl_215_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_32 or ST1_11d or rl_a33_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_217 or ST1_06d or RG_rl_159 or ST1_05d or RG_quantized_block_rl_32 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_216_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h21 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_216_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_32 )
		| ( { 9{ ST1_05d } } & RG_rl_159 )
		| ( { 9{ ST1_06d } } & RG_rl_217 )
		| ( { 9{ RG_rl_216_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a33_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_32 ) ) ;
	end
assign	RG_rl_216_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_216_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_216_en )
		RG_rl_216 <= RG_rl_216_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_33 or ST1_11d or rl_a34_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_218 or ST1_06d or RG_rl_160 or ST1_05d or RG_quantized_block_rl_33 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_217_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h22 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_217_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_33 )
		| ( { 9{ ST1_05d } } & RG_rl_160 )
		| ( { 9{ ST1_06d } } & RG_rl_218 )
		| ( { 9{ RG_rl_217_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a34_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_33 ) ) ;
	end
assign	RG_rl_217_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_217_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_217_en )
		RG_rl_217 <= RG_rl_217_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_34 or ST1_11d or rl_a35_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_219 or ST1_06d or RG_rl_161 or ST1_05d or RG_quantized_block_rl_34 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_218_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h23 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_218_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_34 )
		| ( { 9{ ST1_05d } } & RG_rl_161 )
		| ( { 9{ ST1_06d } } & RG_rl_219 )
		| ( { 9{ RG_rl_218_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a35_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_34 ) ) ;
	end
assign	RG_rl_218_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_218_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_218_en )
		RG_rl_218 <= RG_rl_218_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_35 or ST1_11d or rl_a36_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_220 or ST1_06d or RG_rl_162 or ST1_05d or RG_quantized_block_rl_35 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_219_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h24 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_219_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_35 )
		| ( { 9{ ST1_05d } } & RG_rl_162 )
		| ( { 9{ ST1_06d } } & RG_rl_220 )
		| ( { 9{ RG_rl_219_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a36_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_35 ) ) ;
	end
assign	RG_rl_219_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_219_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_219_en )
		RG_rl_219 <= RG_rl_219_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_36 or ST1_11d or rl_a37_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_221 or ST1_06d or RG_rl_163 or ST1_05d or RG_quantized_block_rl_36 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_220_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h25 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_220_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_36 )
		| ( { 9{ ST1_05d } } & RG_rl_163 )
		| ( { 9{ ST1_06d } } & RG_rl_221 )
		| ( { 9{ RG_rl_220_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a37_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_36 ) ) ;
	end
assign	RG_rl_220_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_220_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_220_en )
		RG_rl_220 <= RG_rl_220_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_37 or ST1_11d or rl_a38_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_222 or ST1_06d or RG_rl_164 or ST1_05d or RG_quantized_block_rl_37 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_221_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h26 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_221_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_37 )
		| ( { 9{ ST1_05d } } & RG_rl_164 )
		| ( { 9{ ST1_06d } } & RG_rl_222 )
		| ( { 9{ RG_rl_221_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a38_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_37 ) ) ;
	end
assign	RG_rl_221_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_221_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_221_en )
		RG_rl_221 <= RG_rl_221_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_38 or ST1_11d or rl_a39_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_223 or ST1_06d or RG_rl_165 or ST1_05d or RG_quantized_block_rl_38 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_222_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h27 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_222_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_38 )
		| ( { 9{ ST1_05d } } & RG_rl_165 )
		| ( { 9{ ST1_06d } } & RG_rl_223 )
		| ( { 9{ RG_rl_222_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a39_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_38 ) ) ;
	end
assign	RG_rl_222_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_222_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_222_en )
		RG_rl_222 <= RG_rl_222_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_39 or ST1_11d or rl_a40_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_224 or ST1_06d or RG_rl_166 or ST1_05d or RG_quantized_block_rl_39 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_223_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h28 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_223_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_39 )
		| ( { 9{ ST1_05d } } & RG_rl_166 )
		| ( { 9{ ST1_06d } } & RG_rl_224 )
		| ( { 9{ RG_rl_223_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a40_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_39 ) ) ;
	end
assign	RG_rl_223_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_223_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_223_en )
		RG_rl_223 <= RG_rl_223_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_40 or ST1_11d or rl_a41_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_225 or ST1_06d or RG_rl_167 or ST1_05d or RG_quantized_block_rl_40 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_224_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h29 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_224_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_40 )
		| ( { 9{ ST1_05d } } & RG_rl_167 )
		| ( { 9{ ST1_06d } } & RG_rl_225 )
		| ( { 9{ RG_rl_224_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a41_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_40 ) ) ;
	end
assign	RG_rl_224_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_224_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_224_en )
		RG_rl_224 <= RG_rl_224_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_41 or ST1_11d or rl_a42_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_226 or ST1_06d or RG_rl_168 or ST1_05d or RG_quantized_block_rl_41 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_225_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h2a ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_225_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_41 )
		| ( { 9{ ST1_05d } } & RG_rl_168 )
		| ( { 9{ ST1_06d } } & RG_rl_226 )
		| ( { 9{ RG_rl_225_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a42_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_41 ) ) ;
	end
assign	RG_rl_225_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_225_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_225_en )
		RG_rl_225 <= RG_rl_225_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_42 or ST1_11d or rl_a43_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_227 or ST1_06d or RG_rl_169 or ST1_05d or RG_quantized_block_rl_42 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_226_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h2b ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_226_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_42 )
		| ( { 9{ ST1_05d } } & RG_rl_169 )
		| ( { 9{ ST1_06d } } & RG_rl_227 )
		| ( { 9{ RG_rl_226_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a43_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_42 ) ) ;
	end
assign	RG_rl_226_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_226_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_226_en )
		RG_rl_226 <= RG_rl_226_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_43 or ST1_11d or rl_a44_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_228 or ST1_06d or RG_rl_170 or ST1_05d or RG_quantized_block_rl_43 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_227_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h2c ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_227_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_43 )
		| ( { 9{ ST1_05d } } & RG_rl_170 )
		| ( { 9{ ST1_06d } } & RG_rl_228 )
		| ( { 9{ RG_rl_227_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a44_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_43 ) ) ;
	end
assign	RG_rl_227_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_227_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_227_en )
		RG_rl_227 <= RG_rl_227_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_44 or ST1_11d or rl_a45_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_229 or ST1_06d or RG_rl_171 or ST1_05d or RG_quantized_block_rl_44 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_228_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h2d ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_228_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_44 )
		| ( { 9{ ST1_05d } } & RG_rl_171 )
		| ( { 9{ ST1_06d } } & RG_rl_229 )
		| ( { 9{ RG_rl_228_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a45_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_44 ) ) ;
	end
assign	RG_rl_228_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_228_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_228_en )
		RG_rl_228 <= RG_rl_228_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_45 or ST1_11d or rl_a46_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_230 or ST1_06d or RG_rl_172 or ST1_05d or RG_quantized_block_rl_45 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_229_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h2e ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_229_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_45 )
		| ( { 9{ ST1_05d } } & RG_rl_172 )
		| ( { 9{ ST1_06d } } & RG_rl_230 )
		| ( { 9{ RG_rl_229_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a46_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_45 ) ) ;
	end
assign	RG_rl_229_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_229_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_229_en )
		RG_rl_229 <= RG_rl_229_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_46 or ST1_11d or rl_a47_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_231 or ST1_06d or RG_rl_173 or ST1_05d or RG_quantized_block_rl_46 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_230_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h2f ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_230_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_46 )
		| ( { 9{ ST1_05d } } & RG_rl_173 )
		| ( { 9{ ST1_06d } } & RG_rl_231 )
		| ( { 9{ RG_rl_230_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a47_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_46 ) ) ;
	end
assign	RG_rl_230_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_230_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_230_en )
		RG_rl_230 <= RG_rl_230_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_47 or ST1_11d or rl_a48_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_232 or ST1_06d or RG_rl_174 or ST1_05d or RG_quantized_block_rl_47 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_231_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h30 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_231_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_47 )
		| ( { 9{ ST1_05d } } & RG_rl_174 )
		| ( { 9{ ST1_06d } } & RG_rl_232 )
		| ( { 9{ RG_rl_231_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a48_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_47 ) ) ;
	end
assign	RG_rl_231_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_231_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_231_en )
		RG_rl_231 <= RG_rl_231_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_48 or ST1_11d or rl_a49_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_233 or ST1_06d or RG_rl_175 or ST1_05d or RG_quantized_block_rl_48 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_232_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h31 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_232_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_48 )
		| ( { 9{ ST1_05d } } & RG_rl_175 )
		| ( { 9{ ST1_06d } } & RG_rl_233 )
		| ( { 9{ RG_rl_232_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a49_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_48 ) ) ;
	end
assign	RG_rl_232_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_232_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_232_en )
		RG_rl_232 <= RG_rl_232_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_49 or ST1_11d or rl_a50_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_234 or ST1_06d or RG_rl_176 or ST1_05d or RG_quantized_block_rl_49 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_233_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h32 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_233_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_49 )
		| ( { 9{ ST1_05d } } & RG_rl_176 )
		| ( { 9{ ST1_06d } } & RG_rl_234 )
		| ( { 9{ RG_rl_233_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a50_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_49 ) ) ;
	end
assign	RG_rl_233_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_233_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_233_en )
		RG_rl_233 <= RG_rl_233_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_50 or ST1_11d or rl_a51_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_235 or ST1_06d or RG_rl_177 or ST1_05d or RG_quantized_block_rl_50 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_234_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h33 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_234_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_50 )
		| ( { 9{ ST1_05d } } & RG_rl_177 )
		| ( { 9{ ST1_06d } } & RG_rl_235 )
		| ( { 9{ RG_rl_234_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a51_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_50 ) ) ;
	end
assign	RG_rl_234_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_234_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_234_en )
		RG_rl_234 <= RG_rl_234_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_51 or ST1_11d or rl_a52_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_236 or ST1_06d or RG_rl_178 or ST1_05d or RG_quantized_block_rl_51 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_235_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h34 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_235_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_51 )
		| ( { 9{ ST1_05d } } & RG_rl_178 )
		| ( { 9{ ST1_06d } } & RG_rl_236 )
		| ( { 9{ RG_rl_235_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a52_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_51 ) ) ;
	end
assign	RG_rl_235_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_235_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_235_en )
		RG_rl_235 <= RG_rl_235_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_52 or ST1_11d or rl_a53_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_237 or ST1_06d or RG_rl_179 or ST1_05d or RG_quantized_block_rl_52 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_236_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h35 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_236_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_52 )
		| ( { 9{ ST1_05d } } & RG_rl_179 )
		| ( { 9{ ST1_06d } } & RG_rl_237 )
		| ( { 9{ RG_rl_236_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a53_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_52 ) ) ;
	end
assign	RG_rl_236_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_236_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_236_en )
		RG_rl_236 <= RG_rl_236_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_53 or ST1_11d or rl_a54_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_238 or ST1_06d or RG_rl_180 or ST1_05d or RG_quantized_block_rl_53 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_237_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h36 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_237_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_53 )
		| ( { 9{ ST1_05d } } & RG_rl_180 )
		| ( { 9{ ST1_06d } } & RG_rl_238 )
		| ( { 9{ RG_rl_237_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a54_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_53 ) ) ;
	end
assign	RG_rl_237_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_237_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_237_en )
		RG_rl_237 <= RG_rl_237_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_54 or ST1_11d or rl_a55_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_239 or ST1_06d or RG_rl_181 or ST1_05d or RG_quantized_block_rl_54 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_238_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h37 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_238_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_54 )
		| ( { 9{ ST1_05d } } & RG_rl_181 )
		| ( { 9{ ST1_06d } } & RG_rl_239 )
		| ( { 9{ RG_rl_238_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a55_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_54 ) ) ;
	end
assign	RG_rl_238_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_238_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_238_en )
		RG_rl_238 <= RG_rl_238_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_55 or ST1_11d or rl_a56_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_240 or ST1_06d or RG_rl_182 or ST1_05d or RG_quantized_block_rl_55 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_239_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h38 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_239_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_55 )
		| ( { 9{ ST1_05d } } & RG_rl_182 )
		| ( { 9{ ST1_06d } } & RG_rl_240 )
		| ( { 9{ RG_rl_239_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a56_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_55 ) ) ;
	end
assign	RG_rl_239_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_239_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_239_en )
		RG_rl_239 <= RG_rl_239_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_56 or ST1_11d or rl_a57_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_241 or ST1_06d or RG_rl_183 or ST1_05d or RG_quantized_block_rl_56 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_240_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h39 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_240_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_56 )
		| ( { 9{ ST1_05d } } & RG_rl_183 )
		| ( { 9{ ST1_06d } } & RG_rl_241 )
		| ( { 9{ RG_rl_240_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a57_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_56 ) ) ;
	end
assign	RG_rl_240_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_240_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_240_en )
		RG_rl_240 <= RG_rl_240_t ;	// line#=../rle.cpp:73
always @ ( RG_rl_57 or ST1_11d or rl_a58_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl or ST1_06d or RG_rl_184 or ST1_05d or RG_quantized_block_rl_57 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_rl_241_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h3a ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_241_t = ( ( { 9{ U_01 } } & RG_quantized_block_rl_57 )
		| ( { 9{ ST1_05d } } & RG_rl_184 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl )
		| ( { 9{ RG_rl_241_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a58_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_57 ) ) ;
	end
assign	RG_rl_241_en = ( U_01 | ST1_05d | ST1_06d | RG_rl_241_t_c1 | ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_241_en )
		RG_rl_241 <= RG_rl_241_t ;	// line#=../rle.cpp:73
always @ ( FF_j or ST1_11d or incr4s1ot or ST1_02d or ST1_01d )
	RG_j_t = ( ( { 4{ ST1_01d } } & 4'hf /*-4'h1*/ )	// line#=../rle.cpp:34
		| ( { 4{ ST1_02d } } & incr4s1ot )		// line#=../rle.cpp:34
		| ( { 4{ ST1_11d } } & { 3'h0 , FF_j } ) ) ;
always @ ( posedge clk )
	RG_j <= RG_j_t ;	// line#=../rle.cpp:34
assign	M_321 = ( M_320 | U_172 ) ;
always @ ( U_06 )
	TR_01 = ( { 3{ U_06 } } & 3'h7 )	// line#=../rle.cpp:134
		 ;	// line#=../rle.cpp:59,105
always @ ( decr32s1ot or U_165 or U_83 or incr32s1ot or U_166 or U_163 or ST1_04d or 
	U_171 or U_84 or U_81 or TR_01 or U_06 or M_321 )
	begin
	RG_i_k_01_t_c1 = ( M_321 | U_06 ) ;	// line#=../rle.cpp:59,105,134
	RG_i_k_01_t_c2 = ( ( ( U_81 | U_84 ) | U_171 ) | ( ST1_04d & ( U_163 | U_166 ) ) ) ;	// line#=../rle.cpp:64,119,129,150,160
	RG_i_k_01_t_c3 = ( U_83 | ( ST1_04d & U_165 ) ) ;	// line#=../rle.cpp:124,155
	RG_i_k_01_t = ( ( { 32{ RG_i_k_01_t_c1 } } & { 29'h00000000 , TR_01 } )	// line#=../rle.cpp:59,105,134
		| ( { 32{ RG_i_k_01_t_c2 } } & incr32s1ot )			// line#=../rle.cpp:64,119,129,150,160
		| ( { 32{ RG_i_k_01_t_c3 } } & decr32s1ot )			// line#=../rle.cpp:124,155
		) ;
	end
assign	RG_i_k_01_en = ( RG_i_k_01_t_c1 | RG_i_k_01_t_c2 | RG_i_k_01_t_c3 ) ;
always @ ( posedge clk )
	if ( RG_i_k_01_en )
		RG_i_k_01 <= RG_i_k_01_t ;	// line#=../rle.cpp:59,64,105,119,124,129
						// ,134,150,155,160
always @ ( FF_i or U_88 or U_06 )
	TR_02 = ( ( { 1{ U_06 } } & 1'h1 )	// line#=../rle.cpp:135
		| ( { 1{ U_88 } } & FF_i )	// line#=../rle.cpp:140,141
		) ;	// line#=../rle.cpp:105
always @ ( i2_t1 or U_172 or decr32s2ot or U_166 or U_84 or incr32s2ot or U_165 or 
	U_161 or U_87 or U_171 or U_83 or U_79 or TR_02 or U_88 or M_319 )
	begin
	RG_i_j_01_t_c1 = ( M_319 | U_88 ) ;	// line#=../rle.cpp:105,135,140,141
	RG_i_j_01_t_c2 = ( ( ( U_79 | U_83 ) | U_171 ) | ( U_87 & ( U_161 | U_165 ) ) ) ;	// line#=../rle.cpp:63,114,125,145,156
	RG_i_j_01_t_c3 = ( U_84 | ( U_87 & U_166 ) ) ;	// line#=../rle.cpp:130,161
	RG_i_j_01_t = ( ( { 32{ RG_i_j_01_t_c1 } } & { 31'h00000000 , TR_02 } )	// line#=../rle.cpp:105,135,140,141
		| ( { 32{ RG_i_j_01_t_c2 } } & incr32s2ot )			// line#=../rle.cpp:63,114,125,145,156
		| ( { 32{ RG_i_j_01_t_c3 } } & decr32s2ot )			// line#=../rle.cpp:130,161
		| ( { 32{ U_172 } } & i2_t1 ) ) ;
	end
assign	RG_i_j_01_en = ( RG_i_j_01_t_c1 | RG_i_j_01_t_c2 | RG_i_j_01_t_c3 | U_172 ) ;
always @ ( posedge clk )
	if ( RG_i_j_01_en )
		RG_i_j_01 <= RG_i_j_01_t ;	// line#=../rle.cpp:63,105,114,125,130
						// ,135,140,141,145,156,161
always @ ( RG_rl_58 or ST1_11d or rl_a59_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_1 or ST1_06d or RG_previous_dc_rl or ST1_05d or 
	jpeg_in_a00 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h3b ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_t = ( ( { 9{ U_01 } } & jpeg_in_a00 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_previous_dc_rl )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_1 )
		| ( { 9{ RG_quantized_block_rl_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a59_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_58 ) ) ;
	end
assign	RG_quantized_block_rl_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_en )
		RG_quantized_block_rl <= RG_quantized_block_rl_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_59 or ST1_11d or rl_a60_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_2 or ST1_06d or RG_rl_185 or ST1_05d or jpeg_in_a01 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_1_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h3c ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_1_t = ( ( { 9{ U_01 } } & jpeg_in_a01 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_185 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_2 )
		| ( { 9{ RG_quantized_block_rl_1_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a60_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_59 ) ) ;
	end
assign	RG_quantized_block_rl_1_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_1_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_1_en )
		RG_quantized_block_rl_1 <= RG_quantized_block_rl_1_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_60 or ST1_11d or rl_a61_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_3 or ST1_06d or RG_rl_186 or ST1_05d or jpeg_in_a02 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_2_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h3d ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_2_t = ( ( { 9{ U_01 } } & jpeg_in_a02 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_186 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_3 )
		| ( { 9{ RG_quantized_block_rl_2_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a61_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_60 ) ) ;
	end
assign	RG_quantized_block_rl_2_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_2_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_2_en )
		RG_quantized_block_rl_2 <= RG_quantized_block_rl_2_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_61 or ST1_11d or rl_a62_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_4 or ST1_06d or RG_rl_187 or ST1_05d or jpeg_in_a03 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_3_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h3e ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_3_t = ( ( { 9{ U_01 } } & jpeg_in_a03 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_187 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_4 )
		| ( { 9{ RG_quantized_block_rl_3_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a62_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_61 ) ) ;
	end
assign	RG_quantized_block_rl_3_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_3_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_3_en )
		RG_quantized_block_rl_3 <= RG_quantized_block_rl_3_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_62 or ST1_11d or rl_a63_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_5 or ST1_06d or RG_rl_188 or ST1_05d or jpeg_in_a04 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_4_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h3f ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_4_t = ( ( { 9{ U_01 } } & jpeg_in_a04 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_188 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_5 )
		| ( { 9{ RG_quantized_block_rl_4_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a63_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_62 ) ) ;
	end
assign	RG_quantized_block_rl_4_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_4_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_4_en )
		RG_quantized_block_rl_4 <= RG_quantized_block_rl_4_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_63 or ST1_11d or rl_a64_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_6 or ST1_06d or RG_rl_189 or ST1_05d or jpeg_in_a05 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_5_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h40 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_5_t = ( ( { 9{ U_01 } } & jpeg_in_a05 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_189 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_6 )
		| ( { 9{ RG_quantized_block_rl_5_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a64_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_63 ) ) ;
	end
assign	RG_quantized_block_rl_5_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_5_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_5_en )
		RG_quantized_block_rl_5 <= RG_quantized_block_rl_5_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_64 or ST1_11d or rl_a65_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_7 or ST1_06d or RG_rl_190 or ST1_05d or jpeg_in_a06 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_6_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h41 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_6_t = ( ( { 9{ U_01 } } & jpeg_in_a06 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_190 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_7 )
		| ( { 9{ RG_quantized_block_rl_6_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a65_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_64 ) ) ;
	end
assign	RG_quantized_block_rl_6_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_6_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_6_en )
		RG_quantized_block_rl_6 <= RG_quantized_block_rl_6_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_65 or ST1_11d or rl_a66_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_8 or ST1_06d or RG_rl_191 or ST1_05d or jpeg_in_a07 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_7_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h42 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_7_t = ( ( { 9{ U_01 } } & jpeg_in_a07 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_191 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_8 )
		| ( { 9{ RG_quantized_block_rl_7_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a66_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_65 ) ) ;
	end
assign	RG_quantized_block_rl_7_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_7_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_7_en )
		RG_quantized_block_rl_7 <= RG_quantized_block_rl_7_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_66 or ST1_11d or rl_a67_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_9 or ST1_06d or RG_rl_192 or ST1_05d or jpeg_in_a08 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_8_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h43 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_8_t = ( ( { 9{ U_01 } } & jpeg_in_a08 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_192 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_9 )
		| ( { 9{ RG_quantized_block_rl_8_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a67_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_66 ) ) ;
	end
assign	RG_quantized_block_rl_8_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_8_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_8_en )
		RG_quantized_block_rl_8 <= RG_quantized_block_rl_8_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_67 or ST1_11d or rl_a68_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_10 or ST1_06d or RG_rl_193 or ST1_05d or 
	jpeg_in_a09 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_9_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h44 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_9_t = ( ( { 9{ U_01 } } & jpeg_in_a09 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_193 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_10 )
		| ( { 9{ RG_quantized_block_rl_9_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a68_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_67 ) ) ;
	end
assign	RG_quantized_block_rl_9_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_9_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_9_en )
		RG_quantized_block_rl_9 <= RG_quantized_block_rl_9_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_68 or ST1_11d or rl_a69_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_11 or ST1_06d or RG_rl_194 or ST1_05d or 
	jpeg_in_a10 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_10_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h45 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_10_t = ( ( { 9{ U_01 } } & jpeg_in_a10 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_194 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_11 )
		| ( { 9{ RG_quantized_block_rl_10_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a69_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_68 ) ) ;
	end
assign	RG_quantized_block_rl_10_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_10_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_10_en )
		RG_quantized_block_rl_10 <= RG_quantized_block_rl_10_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_69 or ST1_11d or rl_a70_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_12 or ST1_06d or RG_rl_195 or ST1_05d or 
	jpeg_in_a11 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_11_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h46 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_11_t = ( ( { 9{ U_01 } } & jpeg_in_a11 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_195 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_12 )
		| ( { 9{ RG_quantized_block_rl_11_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a70_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_69 ) ) ;
	end
assign	RG_quantized_block_rl_11_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_11_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_11_en )
		RG_quantized_block_rl_11 <= RG_quantized_block_rl_11_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_70 or ST1_11d or rl_a71_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_13 or ST1_06d or RG_rl_196 or ST1_05d or 
	jpeg_in_a12 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_12_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h47 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_12_t = ( ( { 9{ U_01 } } & jpeg_in_a12 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_196 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_13 )
		| ( { 9{ RG_quantized_block_rl_12_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a71_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_70 ) ) ;
	end
assign	RG_quantized_block_rl_12_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_12_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_12_en )
		RG_quantized_block_rl_12 <= RG_quantized_block_rl_12_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_71 or ST1_11d or rl_a72_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_14 or ST1_06d or RG_rl_197 or ST1_05d or 
	jpeg_in_a13 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_13_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h48 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_13_t = ( ( { 9{ U_01 } } & jpeg_in_a13 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_197 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_14 )
		| ( { 9{ RG_quantized_block_rl_13_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a72_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_71 ) ) ;
	end
assign	RG_quantized_block_rl_13_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_13_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_13_en )
		RG_quantized_block_rl_13 <= RG_quantized_block_rl_13_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_72 or ST1_11d or rl_a73_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_15 or ST1_06d or RG_rl_198 or ST1_05d or 
	jpeg_in_a14 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_14_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h49 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_14_t = ( ( { 9{ U_01 } } & jpeg_in_a14 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_198 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_15 )
		| ( { 9{ RG_quantized_block_rl_14_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a73_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_72 ) ) ;
	end
assign	RG_quantized_block_rl_14_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_14_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_14_en )
		RG_quantized_block_rl_14 <= RG_quantized_block_rl_14_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_73 or ST1_11d or rl_a74_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_16 or ST1_06d or RG_rl_199 or ST1_05d or 
	jpeg_in_a15 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_15_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h4a ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_15_t = ( ( { 9{ U_01 } } & jpeg_in_a15 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_199 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_16 )
		| ( { 9{ RG_quantized_block_rl_15_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a74_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_73 ) ) ;
	end
assign	RG_quantized_block_rl_15_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_15_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_15_en )
		RG_quantized_block_rl_15 <= RG_quantized_block_rl_15_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_74 or ST1_11d or rl_a75_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_17 or ST1_06d or RG_rl_200 or ST1_05d or 
	jpeg_in_a16 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_16_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h4b ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_16_t = ( ( { 9{ U_01 } } & jpeg_in_a16 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_200 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_17 )
		| ( { 9{ RG_quantized_block_rl_16_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a75_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_74 ) ) ;
	end
assign	RG_quantized_block_rl_16_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_16_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_16_en )
		RG_quantized_block_rl_16 <= RG_quantized_block_rl_16_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_75 or ST1_11d or rl_a76_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_18 or ST1_06d or RG_rl_201 or ST1_05d or 
	jpeg_in_a17 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_17_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h4c ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_17_t = ( ( { 9{ U_01 } } & jpeg_in_a17 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_201 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_18 )
		| ( { 9{ RG_quantized_block_rl_17_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a76_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_75 ) ) ;
	end
assign	RG_quantized_block_rl_17_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_17_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_17_en )
		RG_quantized_block_rl_17 <= RG_quantized_block_rl_17_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_76 or ST1_11d or rl_a77_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_19 or ST1_06d or RG_rl_202 or ST1_05d or 
	jpeg_in_a18 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_18_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h4d ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_18_t = ( ( { 9{ U_01 } } & jpeg_in_a18 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_202 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_19 )
		| ( { 9{ RG_quantized_block_rl_18_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a77_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_76 ) ) ;
	end
assign	RG_quantized_block_rl_18_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_18_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_18_en )
		RG_quantized_block_rl_18 <= RG_quantized_block_rl_18_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_77 or ST1_11d or rl_a78_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_20 or ST1_06d or RG_rl_203 or ST1_05d or 
	jpeg_in_a19 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_19_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h4e ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_19_t = ( ( { 9{ U_01 } } & jpeg_in_a19 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_203 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_20 )
		| ( { 9{ RG_quantized_block_rl_19_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a78_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_77 ) ) ;
	end
assign	RG_quantized_block_rl_19_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_19_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_19_en )
		RG_quantized_block_rl_19 <= RG_quantized_block_rl_19_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_78 or ST1_11d or rl_a79_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_21 or ST1_06d or RG_rl_204 or ST1_05d or 
	jpeg_in_a20 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_20_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h4f ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_20_t = ( ( { 9{ U_01 } } & jpeg_in_a20 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_204 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_21 )
		| ( { 9{ RG_quantized_block_rl_20_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a79_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_78 ) ) ;
	end
assign	RG_quantized_block_rl_20_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_20_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_20_en )
		RG_quantized_block_rl_20 <= RG_quantized_block_rl_20_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_79 or ST1_11d or rl_a80_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_22 or ST1_06d or RG_rl_205 or ST1_05d or 
	jpeg_in_a21 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_21_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h50 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_21_t = ( ( { 9{ U_01 } } & jpeg_in_a21 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_205 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_22 )
		| ( { 9{ RG_quantized_block_rl_21_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a80_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_79 ) ) ;
	end
assign	RG_quantized_block_rl_21_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_21_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_21_en )
		RG_quantized_block_rl_21 <= RG_quantized_block_rl_21_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_80 or ST1_11d or rl_a81_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_23 or ST1_06d or RG_rl_206 or ST1_05d or 
	jpeg_in_a22 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_22_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h51 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_22_t = ( ( { 9{ U_01 } } & jpeg_in_a22 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_206 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_23 )
		| ( { 9{ RG_quantized_block_rl_22_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a81_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_80 ) ) ;
	end
assign	RG_quantized_block_rl_22_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_22_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_22_en )
		RG_quantized_block_rl_22 <= RG_quantized_block_rl_22_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_81 or ST1_11d or rl_a82_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_24 or ST1_06d or RG_rl_207 or ST1_05d or 
	jpeg_in_a23 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_23_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h52 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_23_t = ( ( { 9{ U_01 } } & jpeg_in_a23 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_207 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_24 )
		| ( { 9{ RG_quantized_block_rl_23_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a82_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_81 ) ) ;
	end
assign	RG_quantized_block_rl_23_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_23_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_23_en )
		RG_quantized_block_rl_23 <= RG_quantized_block_rl_23_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_82 or ST1_11d or rl_a83_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_25 or ST1_06d or RG_rl_208 or ST1_05d or 
	jpeg_in_a24 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_24_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h53 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_24_t = ( ( { 9{ U_01 } } & jpeg_in_a24 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_208 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_25 )
		| ( { 9{ RG_quantized_block_rl_24_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a83_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_82 ) ) ;
	end
assign	RG_quantized_block_rl_24_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_24_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_24_en )
		RG_quantized_block_rl_24 <= RG_quantized_block_rl_24_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_83 or ST1_11d or rl_a84_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_26 or ST1_06d or RG_rl_209 or ST1_05d or 
	jpeg_in_a25 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_25_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h54 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_25_t = ( ( { 9{ U_01 } } & jpeg_in_a25 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_209 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_26 )
		| ( { 9{ RG_quantized_block_rl_25_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a84_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_83 ) ) ;
	end
assign	RG_quantized_block_rl_25_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_25_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_25_en )
		RG_quantized_block_rl_25 <= RG_quantized_block_rl_25_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_84 or ST1_11d or rl_a85_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_27 or ST1_06d or RG_rl_210 or ST1_05d or 
	jpeg_in_a26 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_26_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h55 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_26_t = ( ( { 9{ U_01 } } & jpeg_in_a26 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_210 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_27 )
		| ( { 9{ RG_quantized_block_rl_26_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a85_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_84 ) ) ;
	end
assign	RG_quantized_block_rl_26_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_26_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_26_en )
		RG_quantized_block_rl_26 <= RG_quantized_block_rl_26_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_85 or ST1_11d or rl_a86_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_28 or ST1_06d or RG_rl_211 or ST1_05d or 
	jpeg_in_a27 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_27_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h56 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_27_t = ( ( { 9{ U_01 } } & jpeg_in_a27 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_211 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_28 )
		| ( { 9{ RG_quantized_block_rl_27_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a86_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_85 ) ) ;
	end
assign	RG_quantized_block_rl_27_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_27_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_27_en )
		RG_quantized_block_rl_27 <= RG_quantized_block_rl_27_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_86 or ST1_11d or rl_a87_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_29 or ST1_06d or RG_rl_212 or ST1_05d or 
	jpeg_in_a28 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_28_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h57 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_28_t = ( ( { 9{ U_01 } } & jpeg_in_a28 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_212 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_29 )
		| ( { 9{ RG_quantized_block_rl_28_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a87_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_86 ) ) ;
	end
assign	RG_quantized_block_rl_28_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_28_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_28_en )
		RG_quantized_block_rl_28 <= RG_quantized_block_rl_28_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_87 or ST1_11d or rl_a88_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_30 or ST1_06d or RG_rl_213 or ST1_05d or 
	jpeg_in_a29 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_29_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h58 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_29_t = ( ( { 9{ U_01 } } & jpeg_in_a29 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_213 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_30 )
		| ( { 9{ RG_quantized_block_rl_29_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a88_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_87 ) ) ;
	end
assign	RG_quantized_block_rl_29_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_29_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_29_en )
		RG_quantized_block_rl_29 <= RG_quantized_block_rl_29_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_88 or ST1_11d or rl_a89_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_31 or ST1_06d or RG_rl_214 or ST1_05d or 
	jpeg_in_a30 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_30_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h59 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_30_t = ( ( { 9{ U_01 } } & jpeg_in_a30 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_214 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_31 )
		| ( { 9{ RG_quantized_block_rl_30_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a89_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_88 ) ) ;
	end
assign	RG_quantized_block_rl_30_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_30_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_30_en )
		RG_quantized_block_rl_30 <= RG_quantized_block_rl_30_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_89 or ST1_11d or rl_a90_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_32 or ST1_06d or RG_rl_215 or ST1_05d or 
	jpeg_in_a31 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_31_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h5a ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_31_t = ( ( { 9{ U_01 } } & jpeg_in_a31 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_215 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_32 )
		| ( { 9{ RG_quantized_block_rl_31_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a90_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_89 ) ) ;
	end
assign	RG_quantized_block_rl_31_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_31_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_31_en )
		RG_quantized_block_rl_31 <= RG_quantized_block_rl_31_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_90 or ST1_11d or rl_a91_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_33 or ST1_06d or RG_rl_216 or ST1_05d or 
	jpeg_in_a32 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_32_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h5b ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_32_t = ( ( { 9{ U_01 } } & jpeg_in_a32 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_216 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_33 )
		| ( { 9{ RG_quantized_block_rl_32_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a91_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_90 ) ) ;
	end
assign	RG_quantized_block_rl_32_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_32_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_32_en )
		RG_quantized_block_rl_32 <= RG_quantized_block_rl_32_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_91 or ST1_11d or rl_a92_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_34 or ST1_06d or RG_rl_217 or ST1_05d or 
	jpeg_in_a33 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_33_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h5c ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_33_t = ( ( { 9{ U_01 } } & jpeg_in_a33 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_217 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_34 )
		| ( { 9{ RG_quantized_block_rl_33_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a92_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_91 ) ) ;
	end
assign	RG_quantized_block_rl_33_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_33_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_33_en )
		RG_quantized_block_rl_33 <= RG_quantized_block_rl_33_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_92 or ST1_11d or rl_a93_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_35 or ST1_06d or RG_rl_218 or ST1_05d or 
	jpeg_in_a34 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_34_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h5d ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_34_t = ( ( { 9{ U_01 } } & jpeg_in_a34 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_218 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_35 )
		| ( { 9{ RG_quantized_block_rl_34_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a93_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_92 ) ) ;
	end
assign	RG_quantized_block_rl_34_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_34_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_34_en )
		RG_quantized_block_rl_34 <= RG_quantized_block_rl_34_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_93 or ST1_11d or rl_a94_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_36 or ST1_06d or RG_rl_219 or ST1_05d or 
	jpeg_in_a35 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_35_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h5e ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_35_t = ( ( { 9{ U_01 } } & jpeg_in_a35 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_219 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_36 )
		| ( { 9{ RG_quantized_block_rl_35_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a94_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_93 ) ) ;
	end
assign	RG_quantized_block_rl_35_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_35_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_35_en )
		RG_quantized_block_rl_35 <= RG_quantized_block_rl_35_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_94 or ST1_11d or rl_a95_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_37 or ST1_06d or RG_rl_220 or ST1_05d or 
	jpeg_in_a36 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_36_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h5f ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_36_t = ( ( { 9{ U_01 } } & jpeg_in_a36 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_220 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_37 )
		| ( { 9{ RG_quantized_block_rl_36_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a95_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_94 ) ) ;
	end
assign	RG_quantized_block_rl_36_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_36_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_36_en )
		RG_quantized_block_rl_36 <= RG_quantized_block_rl_36_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_95 or ST1_11d or rl_a96_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_38 or ST1_06d or RG_rl_221 or ST1_05d or 
	jpeg_in_a37 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_37_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h60 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_37_t = ( ( { 9{ U_01 } } & jpeg_in_a37 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_221 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_38 )
		| ( { 9{ RG_quantized_block_rl_37_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a96_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_95 ) ) ;
	end
assign	RG_quantized_block_rl_37_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_37_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_37_en )
		RG_quantized_block_rl_37 <= RG_quantized_block_rl_37_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_96 or ST1_11d or rl_a97_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_39 or ST1_06d or RG_rl_222 or ST1_05d or 
	jpeg_in_a38 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_38_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h61 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_38_t = ( ( { 9{ U_01 } } & jpeg_in_a38 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_222 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_39 )
		| ( { 9{ RG_quantized_block_rl_38_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a97_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_96 ) ) ;
	end
assign	RG_quantized_block_rl_38_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_38_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_38_en )
		RG_quantized_block_rl_38 <= RG_quantized_block_rl_38_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_97 or ST1_11d or rl_a98_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_40 or ST1_06d or RG_rl_223 or ST1_05d or 
	jpeg_in_a39 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_39_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h62 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_39_t = ( ( { 9{ U_01 } } & jpeg_in_a39 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_223 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_40 )
		| ( { 9{ RG_quantized_block_rl_39_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a98_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_97 ) ) ;
	end
assign	RG_quantized_block_rl_39_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_39_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_39_en )
		RG_quantized_block_rl_39 <= RG_quantized_block_rl_39_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_98 or ST1_11d or rl_a99_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_41 or ST1_06d or RG_rl_224 or ST1_05d or 
	jpeg_in_a40 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_40_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h63 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_40_t = ( ( { 9{ U_01 } } & jpeg_in_a40 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_224 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_41 )
		| ( { 9{ RG_quantized_block_rl_40_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a99_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_98 ) ) ;
	end
assign	RG_quantized_block_rl_40_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_40_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_40_en )
		RG_quantized_block_rl_40 <= RG_quantized_block_rl_40_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_99 or ST1_11d or rl_a100_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_42 or ST1_06d or RG_rl_225 or ST1_05d or 
	jpeg_in_a41 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_41_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h64 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_41_t = ( ( { 9{ U_01 } } & jpeg_in_a41 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_225 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_42 )
		| ( { 9{ RG_quantized_block_rl_41_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a100_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_99 ) ) ;
	end
assign	RG_quantized_block_rl_41_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_41_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_41_en )
		RG_quantized_block_rl_41 <= RG_quantized_block_rl_41_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_100 or ST1_11d or rl_a101_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_43 or ST1_06d or RG_rl_226 or ST1_05d or 
	jpeg_in_a42 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_42_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h65 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_42_t = ( ( { 9{ U_01 } } & jpeg_in_a42 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_226 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_43 )
		| ( { 9{ RG_quantized_block_rl_42_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a101_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_100 ) ) ;
	end
assign	RG_quantized_block_rl_42_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_42_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_42_en )
		RG_quantized_block_rl_42 <= RG_quantized_block_rl_42_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_101 or ST1_11d or rl_a102_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_44 or ST1_06d or RG_rl_227 or ST1_05d or 
	jpeg_in_a43 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_43_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h66 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_43_t = ( ( { 9{ U_01 } } & jpeg_in_a43 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_227 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_44 )
		| ( { 9{ RG_quantized_block_rl_43_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a102_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_101 ) ) ;
	end
assign	RG_quantized_block_rl_43_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_43_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_43_en )
		RG_quantized_block_rl_43 <= RG_quantized_block_rl_43_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_102 or ST1_11d or rl_a103_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_45 or ST1_06d or RG_rl_228 or ST1_05d or 
	jpeg_in_a44 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_44_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h67 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_44_t = ( ( { 9{ U_01 } } & jpeg_in_a44 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_228 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_45 )
		| ( { 9{ RG_quantized_block_rl_44_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a103_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_102 ) ) ;
	end
assign	RG_quantized_block_rl_44_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_44_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_44_en )
		RG_quantized_block_rl_44 <= RG_quantized_block_rl_44_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_103 or ST1_11d or rl_a104_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_46 or ST1_06d or RG_rl_229 or ST1_05d or 
	jpeg_in_a45 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_45_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h68 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_45_t = ( ( { 9{ U_01 } } & jpeg_in_a45 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_229 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_46 )
		| ( { 9{ RG_quantized_block_rl_45_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a104_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_103 ) ) ;
	end
assign	RG_quantized_block_rl_45_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_45_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_45_en )
		RG_quantized_block_rl_45 <= RG_quantized_block_rl_45_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_104 or ST1_11d or rl_a105_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_47 or ST1_06d or RG_rl_230 or ST1_05d or 
	jpeg_in_a46 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_46_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h69 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_46_t = ( ( { 9{ U_01 } } & jpeg_in_a46 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_230 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_47 )
		| ( { 9{ RG_quantized_block_rl_46_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a105_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_104 ) ) ;
	end
assign	RG_quantized_block_rl_46_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_46_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_46_en )
		RG_quantized_block_rl_46 <= RG_quantized_block_rl_46_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_105 or ST1_11d or rl_a106_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_48 or ST1_06d or RG_rl_231 or ST1_05d or 
	jpeg_in_a47 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_47_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h6a ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_47_t = ( ( { 9{ U_01 } } & jpeg_in_a47 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_231 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_48 )
		| ( { 9{ RG_quantized_block_rl_47_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a106_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_105 ) ) ;
	end
assign	RG_quantized_block_rl_47_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_47_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_47_en )
		RG_quantized_block_rl_47 <= RG_quantized_block_rl_47_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_106 or ST1_11d or rl_a107_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_49 or ST1_06d or RG_rl_232 or ST1_05d or 
	jpeg_in_a48 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_48_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h6b ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_48_t = ( ( { 9{ U_01 } } & jpeg_in_a48 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_232 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_49 )
		| ( { 9{ RG_quantized_block_rl_48_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a107_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_106 ) ) ;
	end
assign	RG_quantized_block_rl_48_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_48_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_48_en )
		RG_quantized_block_rl_48 <= RG_quantized_block_rl_48_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_107 or ST1_11d or rl_a108_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_50 or ST1_06d or RG_rl_233 or ST1_05d or 
	jpeg_in_a49 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_49_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h6c ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_49_t = ( ( { 9{ U_01 } } & jpeg_in_a49 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_233 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_50 )
		| ( { 9{ RG_quantized_block_rl_49_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a108_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_107 ) ) ;
	end
assign	RG_quantized_block_rl_49_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_49_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_49_en )
		RG_quantized_block_rl_49 <= RG_quantized_block_rl_49_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_108 or ST1_11d or rl_a109_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_51 or ST1_06d or RG_rl_234 or ST1_05d or 
	jpeg_in_a50 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_50_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h6d ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_50_t = ( ( { 9{ U_01 } } & jpeg_in_a50 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_234 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_51 )
		| ( { 9{ RG_quantized_block_rl_50_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a109_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_108 ) ) ;
	end
assign	RG_quantized_block_rl_50_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_50_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_50_en )
		RG_quantized_block_rl_50 <= RG_quantized_block_rl_50_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_109 or ST1_11d or rl_a110_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_52 or ST1_06d or RG_rl_235 or ST1_05d or 
	jpeg_in_a51 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_51_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h6e ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_51_t = ( ( { 9{ U_01 } } & jpeg_in_a51 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_235 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_52 )
		| ( { 9{ RG_quantized_block_rl_51_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a110_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_109 ) ) ;
	end
assign	RG_quantized_block_rl_51_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_51_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_51_en )
		RG_quantized_block_rl_51 <= RG_quantized_block_rl_51_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_110 or ST1_11d or rl_a111_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_53 or ST1_06d or RG_rl_236 or ST1_05d or 
	jpeg_in_a52 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_52_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h6f ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_52_t = ( ( { 9{ U_01 } } & jpeg_in_a52 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_236 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_53 )
		| ( { 9{ RG_quantized_block_rl_52_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a111_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_110 ) ) ;
	end
assign	RG_quantized_block_rl_52_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_52_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_52_en )
		RG_quantized_block_rl_52 <= RG_quantized_block_rl_52_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_111 or ST1_11d or rl_a112_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_54 or ST1_06d or RG_rl_237 or ST1_05d or 
	jpeg_in_a53 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_53_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h70 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_53_t = ( ( { 9{ U_01 } } & jpeg_in_a53 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_237 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_54 )
		| ( { 9{ RG_quantized_block_rl_53_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a112_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_111 ) ) ;
	end
assign	RG_quantized_block_rl_53_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_53_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_53_en )
		RG_quantized_block_rl_53 <= RG_quantized_block_rl_53_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_112 or ST1_11d or rl_a113_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_55 or ST1_06d or RG_rl_238 or ST1_05d or 
	jpeg_in_a54 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_54_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h71 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_54_t = ( ( { 9{ U_01 } } & jpeg_in_a54 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_238 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_55 )
		| ( { 9{ RG_quantized_block_rl_54_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a113_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_112 ) ) ;
	end
assign	RG_quantized_block_rl_54_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_54_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_54_en )
		RG_quantized_block_rl_54 <= RG_quantized_block_rl_54_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_113 or ST1_11d or rl_a114_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_56 or ST1_06d or RG_rl_239 or ST1_05d or 
	jpeg_in_a55 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_55_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h72 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_55_t = ( ( { 9{ U_01 } } & jpeg_in_a55 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_239 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_56 )
		| ( { 9{ RG_quantized_block_rl_55_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a114_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_113 ) ) ;
	end
assign	RG_quantized_block_rl_55_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_55_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_55_en )
		RG_quantized_block_rl_55 <= RG_quantized_block_rl_55_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_114 or ST1_11d or rl_a115_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_quantized_block_rl_57 or ST1_06d or RG_rl_240 or ST1_05d or 
	jpeg_in_a56 or U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_56_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h73 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_56_t = ( ( { 9{ U_01 } } & jpeg_in_a56 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_240 )
		| ( { 9{ ST1_06d } } & RG_quantized_block_rl_57 )
		| ( { 9{ RG_quantized_block_rl_56_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a115_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_114 ) ) ;
	end
assign	RG_quantized_block_rl_56_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_56_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_56_en )
		RG_quantized_block_rl_56 <= RG_quantized_block_rl_56_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_115 or ST1_11d or rl_a117_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_242 or ST1_06d or RG_rl_241 or ST1_05d or jpeg_in_a57 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_57_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h75 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_57_t = ( ( { 9{ U_01 } } & jpeg_in_a57 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_241 )
		| ( { 9{ ST1_06d } } & RG_rl_242 )
		| ( { 9{ RG_quantized_block_rl_57_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a117_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_115 ) ) ;
	end
assign	RG_quantized_block_rl_57_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_57_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_57_en )
		RG_quantized_block_rl_57 <= RG_quantized_block_rl_57_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_117 or ST1_11d or rl_a119_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_243 or ST1_06d or RG_rl_116 or ST1_05d or jpeg_in_a58 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_58_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h77 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_58_t = ( ( { 9{ U_01 } } & jpeg_in_a58 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_116 )
		| ( { 9{ ST1_06d } } & RG_rl_243 )
		| ( { 9{ RG_quantized_block_rl_58_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a119_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_117 ) ) ;
	end
assign	RG_quantized_block_rl_58_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_58_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_58_en )
		RG_quantized_block_rl_58 <= RG_quantized_block_rl_58_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_119 or ST1_11d or rl_a121_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_244 or ST1_06d or RG_rl_118 or ST1_05d or jpeg_in_a59 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_59_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h79 ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_59_t = ( ( { 9{ U_01 } } & jpeg_in_a59 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_118 )
		| ( { 9{ ST1_06d } } & RG_rl_244 )
		| ( { 9{ RG_quantized_block_rl_59_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a121_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_119 ) ) ;
	end
assign	RG_quantized_block_rl_59_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_59_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_59_en )
		RG_quantized_block_rl_59 <= RG_quantized_block_rl_59_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_121 or ST1_11d or rl_a123_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_245 or ST1_06d or RG_rl_120 or ST1_05d or jpeg_in_a60 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_60_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h7b ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_60_t = ( ( { 9{ U_01 } } & jpeg_in_a60 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_120 )
		| ( { 9{ ST1_06d } } & RG_rl_245 )
		| ( { 9{ RG_quantized_block_rl_60_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a123_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_121 ) ) ;
	end
assign	RG_quantized_block_rl_60_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_60_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_60_en )
		RG_quantized_block_rl_60 <= RG_quantized_block_rl_60_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_123 or ST1_11d or rl_a125_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_rl_246 or ST1_06d or RG_rl_122 or ST1_05d or jpeg_in_a61 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_61_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h7d ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_61_t = ( ( { 9{ U_01 } } & jpeg_in_a61 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_122 )
		| ( { 9{ ST1_06d } } & RG_rl_246 )
		| ( { 9{ RG_quantized_block_rl_61_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a125_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_123 ) ) ;
	end
assign	RG_quantized_block_rl_61_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_61_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_61_en )
		RG_quantized_block_rl_61 <= RG_quantized_block_rl_61_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_125 or ST1_11d or rl_a127_t4 or ST1_09d or RG_i_k_01 or RG_len or 
	U_174 or RG_previous_dc_rl_1 or ST1_06d or RG_rl_124 or ST1_05d or jpeg_in_a62 or 
	U_01 )	// line#=../rle.cpp:73
	begin
	RG_quantized_block_rl_62_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h7f ) ) ) ;	// line#=../rle.cpp:73
	RG_quantized_block_rl_62_t = ( ( { 9{ U_01 } } & jpeg_in_a62 )		// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_124 )
		| ( { 9{ ST1_06d } } & RG_previous_dc_rl_1 )
		| ( { 9{ RG_quantized_block_rl_62_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a127_t4 )
		| ( { 9{ ST1_11d } } & RG_rl_125 ) ) ;
	end
assign	RG_quantized_block_rl_62_en = ( U_01 | ST1_05d | ST1_06d | RG_quantized_block_rl_62_t_c1 | 
	ST1_09d | ST1_11d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_quantized_block_rl_62_en )
		RG_quantized_block_rl_62 <= RG_quantized_block_rl_62_t ;	// line#=../rle.cpp:45,73
always @ ( RG_rl_127 or U_572 or zz_RD1 or ST1_06d or RG_rl_126 or ST1_05d or jpeg_in_a63 or 
	U_01 )
	RL_previous_dc_quantized_block_t = ( ( { 9{ U_01 } } & jpeg_in_a63 )	// line#=../rle.cpp:45
		| ( { 9{ ST1_05d } } & RG_rl_126 )
		| ( { 9{ ST1_06d } } & zz_RD1 )					// line#=../rle.cpp:52,53
		| ( { 9{ U_572 } } & RG_rl_127 ) ) ;
assign	RL_previous_dc_quantized_block_en = ( U_01 | ST1_05d | ST1_06d | U_572 ) ;
always @ ( posedge clk )
	if ( RL_previous_dc_quantized_block_en )
		RL_previous_dc_quantized_block <= RL_previous_dc_quantized_block_t ;	// line#=../rle.cpp:45,52,53
always @ ( sub8u1ot or ST1_09d or incr8u1ot or U_172 or incr8u3ot or ST1_04d or 
	U_05 )
	begin
	RG_k_01_t_c1 = ( U_05 | ST1_04d ) ;	// line#=../rle.cpp:111,142
	RG_k_01_t = ( ( { 7{ RG_k_01_t_c1 } } & incr8u3ot [6:0] )	// line#=../rle.cpp:111,142
		| ( { 7{ U_172 } } & incr8u1ot [6:0] )			// line#=../rle.cpp:68,69,73,74
		| ( { 7{ ST1_09d } } & sub8u1ot [6:0] )			// line#=../rle.cpp:77,78
		) ;	// line#=../rle.cpp:105
	end
assign	RG_k_01_en = ( ST1_02d | RG_k_01_t_c1 | U_172 | ST1_09d ) ;
always @ ( posedge clk )
	if ( RG_k_01_en )
		RG_k_01 <= RG_k_01_t ;	// line#=../rle.cpp:68,69,73,74,77,78,105
					// ,111,142
assign	M_319 = ( ST1_02d | U_06 ) ;
always @ ( CT_33 or ST1_08d or U_163 or U_79 or U_161 or ST1_04d or U_81 or M_319 )
	begin
	FF_d_01_t_c1 = ( ( M_319 | U_81 ) | ( ST1_04d & U_161 ) ) ;	// line#=../rle.cpp:105,120,136,146
	FF_d_01_t_c2 = ( U_79 | ( ST1_04d & U_163 ) ) ;	// line#=../rle.cpp:115,151
	FF_d_01_t = ( ( { 1{ FF_d_01_t_c2 } } & 1'h1 )	// line#=../rle.cpp:115,151
		| ( { 1{ ST1_08d } } & CT_33 )		// line#=../rle.cpp:61,62
		) ;	// line#=../rle.cpp:105,120,136,146
	end
assign	FF_d_01_en = ( FF_d_01_t_c1 | FF_d_01_t_c2 | ST1_08d ) ;
always @ ( posedge clk )
	if ( FF_d_01_en )
		FF_d_01 <= FF_d_01_t ;	// line#=../rle.cpp:61,62,105,115,120,136
					// ,146,151
assign	FF_j_en = ST1_02d ;
always @ ( posedge clk )	// line#=../rle.cpp:36
	if ( FF_j_en )
		FF_j <= 1'h0 ;
always @ ( M_317 or ST1_09d or CT_32 or ST1_08d or CT_28 or ST1_07d or ST1_02d )
	FF_i_t = ( ( { 1{ ST1_02d } } & 1'h1 )	// line#=../rle.cpp:37
		| ( { 1{ ST1_07d } } & CT_28 )	// line#=../rle.cpp:61,62
		| ( { 1{ ST1_08d } } & CT_32 )	// line#=../rle.cpp:66,67
		| ( { 1{ ST1_09d } } & M_317 )	// line#=../rle.cpp:77,78
		) ;
assign	FF_i_en = ( ST1_02d | ST1_07d | ST1_08d | ST1_09d ) ;
always @ ( posedge clk )
	if ( FF_i_en )
		FF_i <= FF_i_t ;	// line#=../rle.cpp:37,61,62,66,67,77,78
assign	RG_315_en = ST1_08d ;
always @ ( posedge clk )	// line#=../rle.cpp:57,58
	if ( RG_315_en )
		RG_315 <= ( i2_t1 [31] | ( ~|i2_t1 [30:6] ) ) ;
assign	RG_315_port = RG_315 ;
assign	M_320 = ( ST1_02d | ST1_06d ) ;	// line#=../rle.cpp:73
always @ ( rl_a116_t4 or ST1_09d or RG_i_k_01 or RG_len or U_174 or RG_quantized_block_rl_58 or 
	M_320 )	// line#=../rle.cpp:73
	begin
	RG_rl_242_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h74 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_242_t = ( ( { 9{ M_320 } } & RG_quantized_block_rl_58 )
		| ( { 9{ RG_rl_242_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a116_t4 ) ) ;
	end
assign	RG_rl_242_en = ( M_320 | RG_rl_242_t_c1 | ST1_09d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_242_en )
		RG_rl_242 <= RG_rl_242_t ;	// line#=../rle.cpp:73
always @ ( rl_a118_t4 or ST1_09d or RG_i_k_01 or RG_len or U_174 or RG_quantized_block_rl_59 or 
	M_320 )	// line#=../rle.cpp:73
	begin
	RG_rl_243_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h76 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_243_t = ( ( { 9{ M_320 } } & RG_quantized_block_rl_59 )
		| ( { 9{ RG_rl_243_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a118_t4 ) ) ;
	end
assign	RG_rl_243_en = ( M_320 | RG_rl_243_t_c1 | ST1_09d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_243_en )
		RG_rl_243 <= RG_rl_243_t ;	// line#=../rle.cpp:73
always @ ( rl_a120_t4 or ST1_09d or RG_i_k_01 or RG_len or U_174 or RG_quantized_block_rl_60 or 
	M_320 )	// line#=../rle.cpp:73
	begin
	RG_rl_244_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h78 ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_244_t = ( ( { 9{ M_320 } } & RG_quantized_block_rl_60 )
		| ( { 9{ RG_rl_244_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a120_t4 ) ) ;
	end
assign	RG_rl_244_en = ( M_320 | RG_rl_244_t_c1 | ST1_09d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_244_en )
		RG_rl_244 <= RG_rl_244_t ;	// line#=../rle.cpp:73
always @ ( rl_a122_t4 or ST1_09d or RG_i_k_01 or RG_len or U_174 or RG_quantized_block_rl_61 or 
	M_320 )	// line#=../rle.cpp:73
	begin
	RG_rl_245_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h7a ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_245_t = ( ( { 9{ M_320 } } & RG_quantized_block_rl_61 )
		| ( { 9{ RG_rl_245_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a122_t4 ) ) ;
	end
assign	RG_rl_245_en = ( M_320 | RG_rl_245_t_c1 | ST1_09d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_245_en )
		RG_rl_245 <= RG_rl_245_t ;	// line#=../rle.cpp:73
always @ ( rl_a124_t4 or ST1_09d or RG_i_k_01 or RG_len or U_174 or RG_quantized_block_rl_62 or 
	M_320 )	// line#=../rle.cpp:73
	begin
	RG_rl_246_t_c1 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h7c ) ) ) ;	// line#=../rle.cpp:73
	RG_rl_246_t = ( ( { 9{ M_320 } } & RG_quantized_block_rl_62 )
		| ( { 9{ RG_rl_246_t_c1 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a124_t4 ) ) ;
	end
assign	RG_rl_246_en = ( M_320 | RG_rl_246_t_c1 | ST1_09d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_rl_246_en )
		RG_rl_246 <= RG_rl_246_t ;	// line#=../rle.cpp:73
always @ ( rl_a126_t4 or ST1_09d or RG_i_k_01 or RG_len or U_174 or RL_previous_dc_quantized_block or 
	ST1_11d or ST1_06d or U_01 or RG_previous_dc_rl or ST1_01d )	// line#=../rle.cpp:73
	begin
	RG_previous_dc_rl_1_t_c1 = ( ( U_01 | ST1_06d ) | ST1_11d ) ;
	RG_previous_dc_rl_1_t_c2 = ( U_174 & ( ~|( RG_len [6:0] ^ 7'h7e ) ) ) ;	// line#=../rle.cpp:73
	RG_previous_dc_rl_1_t = ( ( { 9{ ST1_01d } } & RG_previous_dc_rl )
		| ( { 9{ RG_previous_dc_rl_1_t_c1 } } & RL_previous_dc_quantized_block )
		| ( { 9{ RG_previous_dc_rl_1_t_c2 } } & RG_i_k_01 [8:0] )	// line#=../rle.cpp:73
		| ( { 9{ ST1_09d } } & rl_a126_t4 ) ) ;
	end
assign	RG_previous_dc_rl_1_en = ( ST1_01d | RG_previous_dc_rl_1_t_c1 | RG_previous_dc_rl_1_t_c2 | 
	ST1_09d ) ;	// line#=../rle.cpp:73
always @ ( posedge clk )	// line#=../rle.cpp:73
	if ( RG_previous_dc_rl_1_en )
		RG_previous_dc_rl_1 <= RG_previous_dc_rl_1_t ;	// line#=../rle.cpp:73
assign	RG_len_01_en = ST1_04d ;
always @ ( posedge clk )	// line#=../rle.cpp:140,141
	if ( RG_len_01_en )
		RG_len_01 <= { 7'h00 , FF_len } ;
always @ ( sub8u1ot or ST1_11d or incr8u4ot or U_569 or len1_t3 or ST1_09d or incr8u1ot or 
	U_174 or incr8u2ot or U_173 or RG_len_01 or ST1_06d )
	RG_len_t = ( ( { 8{ ST1_06d } } & RG_len_01 )
		| ( { 8{ U_173 } } & incr8u2ot )	// line#=../rle.cpp:69
		| ( { 8{ U_174 } } & incr8u1ot )	// line#=../rle.cpp:73
		| ( { 8{ ST1_09d } } & len1_t3 )
		| ( { 8{ U_569 } } & incr8u4ot )	// line#=../rle.cpp:80
		| ( { 8{ ST1_11d } } & sub8u1ot )	// line#=../rle.cpp:86
		) ;
assign	RG_len_en = ( ST1_06d | U_173 | U_174 | ST1_09d | U_569 | ST1_11d ) ;
always @ ( posedge clk )
	if ( RG_len_en )
		RG_len <= RG_len_t ;	// line#=../rle.cpp:69,73,80,86
always @ ( M_316 or ST1_09d or RG_i_k_01 or ST1_07d or ST1_02d )
	FF_len_t = ( ( { 1{ ST1_02d } } & 1'h1 )		// line#=../rle.cpp:39
		| ( { 1{ ST1_07d } } & ( ~|RG_i_k_01 [30:4] ) )	// line#=../rle.cpp:61,62
		| ( { 1{ ST1_09d } } & M_316 )			// line#=../rle.cpp:77,78
		) ;
assign	FF_len_en = ( ST1_02d | ST1_07d | ST1_09d ) ;
always @ ( posedge clk )
	if ( FF_len_en )
		FF_len <= FF_len_t ;	// line#=../rle.cpp:39,61,62,77,78
assign	JF_01 = ~C_01 ;	// line#=../rle.cpp:35
assign	JF_03 = ~RG_k_01 [6] ;
always @ ( incr32s3ot or RG_i_j_01 or CT_32 )
	begin
	i2_t1_c1 = ~CT_32 ;	// line#=../rle.cpp:74
	i2_t1 = ( ( { 32{ CT_32 } } & RG_i_j_01 )
		| ( { 32{ i2_t1_c1 } } & incr32s3ot )	// line#=../rle.cpp:74
		) ;
	end
always @ ( incr8u3ot or RG_len or FF_i )
	begin
	len1_t3_c1 = ~FF_i ;	// line#=../rle.cpp:74
	len1_t3 = ( ( { 8{ FF_i } } & RG_len )		// line#=../rle.cpp:69
		| ( { 8{ len1_t3_c1 } } & incr8u3ot )	// line#=../rle.cpp:74
		) ;
	end
always @ ( RG_rl_184 or zz_RD1 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a00_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h01 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h02 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h03 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h04 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h05 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h06 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h07 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h08 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h09 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h0a :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h0b :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h0c :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h0d :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h0e :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h0f :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h10 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h11 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h12 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h13 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h14 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h15 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h16 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h17 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h18 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h19 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h1a :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h1b :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h1c :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h1d :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h1e :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h1f :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h20 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h21 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h22 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h23 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h24 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h25 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h26 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h27 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h28 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h29 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h2a :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h2b :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h2c :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h2d :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h2e :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h2f :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h30 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h31 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h32 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h33 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h34 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h35 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h36 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h37 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h38 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h39 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h3a :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h3b :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h3c :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h3d :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h3e :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h3f :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h40 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h41 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h42 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h43 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h44 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h45 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h46 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h47 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h48 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h49 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h4a :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h4b :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h4c :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h4d :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h4e :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h4f :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h50 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h51 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h52 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h53 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h54 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h55 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h56 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h57 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h58 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h59 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h5a :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h5b :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h5c :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h5d :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h5e :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h5f :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h60 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h61 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h62 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h63 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h64 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h65 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h66 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h67 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h68 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h69 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h6a :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h6b :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h6c :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h6d :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h6e :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h6f :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h70 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h71 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h72 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h73 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h74 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h75 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h76 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h77 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h78 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h79 :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h7a :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h7b :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h7c :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h7d :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h7e :
		rl_a00_t4_t1 = RG_rl_184 ;
	7'h7f :
		rl_a00_t4_t1 = RG_rl_184 ;
	default :
		rl_a00_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a00_t4_t1 or rl_a00_t5 or FF_i )
	begin
	rl_a00_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a00_t4 = ( ( { 9{ FF_i } } & rl_a00_t5 )
		| ( { 9{ rl_a00_t4_c1 } } & rl_a00_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_previous_dc_rl or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h01 :
		rl_a01_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h02 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h03 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h04 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h05 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h06 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h07 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h08 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h09 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h0a :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h0b :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h0c :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h0d :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h0e :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h0f :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h10 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h11 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h12 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h13 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h14 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h15 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h16 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h17 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h18 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h19 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h1a :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h1b :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h1c :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h1d :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h1e :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h1f :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h20 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h21 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h22 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h23 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h24 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h25 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h26 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h27 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h28 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h29 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h2a :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h2b :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h2c :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h2d :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h2e :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h2f :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h30 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h31 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h32 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h33 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h34 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h35 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h36 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h37 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h38 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h39 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h3a :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h3b :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h3c :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h3d :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h3e :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h3f :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h40 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h41 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h42 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h43 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h44 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h45 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h46 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h47 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h48 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h49 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h4a :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h4b :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h4c :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h4d :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h4e :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h4f :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h50 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h51 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h52 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h53 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h54 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h55 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h56 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h57 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h58 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h59 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h5a :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h5b :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h5c :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h5d :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h5e :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h5f :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h60 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h61 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h62 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h63 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h64 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h65 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h66 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h67 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h68 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h69 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h6a :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h6b :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h6c :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h6d :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h6e :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h6f :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h70 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h71 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h72 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h73 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h74 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h75 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h76 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h77 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h78 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h79 :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h7a :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h7b :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h7c :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h7d :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h7e :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	7'h7f :
		rl_a01_t4_t1 = RG_previous_dc_rl ;
	default :
		rl_a01_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a01_t4_t1 or rl_a01_t5 or FF_i )
	begin
	rl_a01_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a01_t4 = ( ( { 9{ FF_i } } & rl_a01_t5 )
		| ( { 9{ rl_a01_t4_c1 } } & rl_a01_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_185 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h01 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h02 :
		rl_a02_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h03 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h04 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h05 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h06 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h07 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h08 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h09 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h0a :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h0b :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h0c :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h0d :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h0e :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h0f :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h10 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h11 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h12 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h13 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h14 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h15 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h16 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h17 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h18 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h19 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h1a :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h1b :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h1c :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h1d :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h1e :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h1f :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h20 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h21 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h22 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h23 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h24 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h25 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h26 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h27 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h28 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h29 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h2a :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h2b :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h2c :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h2d :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h2e :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h2f :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h30 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h31 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h32 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h33 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h34 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h35 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h36 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h37 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h38 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h39 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h3a :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h3b :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h3c :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h3d :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h3e :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h3f :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h40 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h41 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h42 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h43 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h44 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h45 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h46 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h47 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h48 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h49 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h4a :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h4b :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h4c :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h4d :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h4e :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h4f :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h50 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h51 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h52 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h53 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h54 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h55 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h56 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h57 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h58 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h59 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h5a :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h5b :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h5c :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h5d :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h5e :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h5f :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h60 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h61 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h62 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h63 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h64 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h65 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h66 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h67 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h68 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h69 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h6a :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h6b :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h6c :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h6d :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h6e :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h6f :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h70 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h71 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h72 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h73 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h74 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h75 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h76 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h77 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h78 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h79 :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h7a :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h7b :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h7c :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h7d :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h7e :
		rl_a02_t4_t1 = RG_rl_185 ;
	7'h7f :
		rl_a02_t4_t1 = RG_rl_185 ;
	default :
		rl_a02_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a02_t4_t1 or rl_a02_t5 or FF_i )
	begin
	rl_a02_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a02_t4 = ( ( { 9{ FF_i } } & rl_a02_t5 )
		| ( { 9{ rl_a02_t4_c1 } } & rl_a02_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_186 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h01 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h02 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h03 :
		rl_a03_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h04 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h05 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h06 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h07 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h08 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h09 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h0a :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h0b :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h0c :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h0d :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h0e :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h0f :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h10 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h11 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h12 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h13 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h14 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h15 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h16 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h17 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h18 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h19 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h1a :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h1b :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h1c :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h1d :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h1e :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h1f :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h20 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h21 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h22 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h23 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h24 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h25 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h26 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h27 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h28 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h29 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h2a :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h2b :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h2c :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h2d :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h2e :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h2f :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h30 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h31 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h32 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h33 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h34 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h35 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h36 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h37 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h38 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h39 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h3a :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h3b :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h3c :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h3d :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h3e :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h3f :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h40 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h41 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h42 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h43 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h44 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h45 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h46 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h47 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h48 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h49 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h4a :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h4b :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h4c :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h4d :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h4e :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h4f :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h50 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h51 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h52 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h53 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h54 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h55 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h56 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h57 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h58 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h59 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h5a :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h5b :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h5c :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h5d :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h5e :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h5f :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h60 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h61 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h62 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h63 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h64 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h65 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h66 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h67 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h68 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h69 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h6a :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h6b :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h6c :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h6d :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h6e :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h6f :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h70 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h71 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h72 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h73 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h74 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h75 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h76 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h77 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h78 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h79 :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h7a :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h7b :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h7c :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h7d :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h7e :
		rl_a03_t4_t1 = RG_rl_186 ;
	7'h7f :
		rl_a03_t4_t1 = RG_rl_186 ;
	default :
		rl_a03_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a03_t4_t1 or rl_a03_t5 or FF_i )
	begin
	rl_a03_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a03_t4 = ( ( { 9{ FF_i } } & rl_a03_t5 )
		| ( { 9{ rl_a03_t4_c1 } } & rl_a03_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_187 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h01 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h02 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h03 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h04 :
		rl_a04_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h05 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h06 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h07 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h08 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h09 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h0a :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h0b :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h0c :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h0d :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h0e :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h0f :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h10 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h11 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h12 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h13 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h14 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h15 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h16 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h17 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h18 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h19 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h1a :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h1b :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h1c :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h1d :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h1e :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h1f :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h20 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h21 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h22 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h23 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h24 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h25 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h26 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h27 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h28 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h29 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h2a :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h2b :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h2c :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h2d :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h2e :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h2f :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h30 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h31 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h32 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h33 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h34 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h35 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h36 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h37 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h38 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h39 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h3a :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h3b :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h3c :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h3d :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h3e :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h3f :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h40 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h41 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h42 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h43 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h44 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h45 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h46 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h47 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h48 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h49 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h4a :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h4b :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h4c :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h4d :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h4e :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h4f :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h50 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h51 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h52 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h53 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h54 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h55 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h56 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h57 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h58 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h59 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h5a :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h5b :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h5c :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h5d :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h5e :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h5f :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h60 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h61 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h62 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h63 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h64 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h65 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h66 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h67 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h68 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h69 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h6a :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h6b :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h6c :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h6d :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h6e :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h6f :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h70 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h71 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h72 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h73 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h74 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h75 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h76 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h77 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h78 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h79 :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h7a :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h7b :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h7c :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h7d :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h7e :
		rl_a04_t4_t1 = RG_rl_187 ;
	7'h7f :
		rl_a04_t4_t1 = RG_rl_187 ;
	default :
		rl_a04_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a04_t4_t1 or rl_a04_t5 or FF_i )
	begin
	rl_a04_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a04_t4 = ( ( { 9{ FF_i } } & rl_a04_t5 )
		| ( { 9{ rl_a04_t4_c1 } } & rl_a04_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_188 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h01 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h02 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h03 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h04 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h05 :
		rl_a05_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h06 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h07 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h08 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h09 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h0a :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h0b :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h0c :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h0d :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h0e :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h0f :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h10 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h11 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h12 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h13 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h14 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h15 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h16 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h17 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h18 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h19 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h1a :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h1b :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h1c :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h1d :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h1e :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h1f :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h20 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h21 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h22 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h23 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h24 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h25 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h26 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h27 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h28 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h29 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h2a :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h2b :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h2c :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h2d :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h2e :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h2f :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h30 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h31 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h32 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h33 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h34 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h35 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h36 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h37 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h38 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h39 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h3a :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h3b :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h3c :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h3d :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h3e :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h3f :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h40 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h41 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h42 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h43 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h44 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h45 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h46 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h47 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h48 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h49 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h4a :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h4b :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h4c :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h4d :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h4e :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h4f :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h50 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h51 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h52 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h53 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h54 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h55 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h56 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h57 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h58 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h59 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h5a :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h5b :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h5c :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h5d :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h5e :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h5f :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h60 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h61 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h62 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h63 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h64 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h65 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h66 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h67 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h68 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h69 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h6a :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h6b :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h6c :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h6d :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h6e :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h6f :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h70 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h71 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h72 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h73 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h74 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h75 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h76 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h77 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h78 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h79 :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h7a :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h7b :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h7c :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h7d :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h7e :
		rl_a05_t4_t1 = RG_rl_188 ;
	7'h7f :
		rl_a05_t4_t1 = RG_rl_188 ;
	default :
		rl_a05_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a05_t4_t1 or rl_a05_t5 or FF_i )
	begin
	rl_a05_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a05_t4 = ( ( { 9{ FF_i } } & rl_a05_t5 )
		| ( { 9{ rl_a05_t4_c1 } } & rl_a05_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_189 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h01 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h02 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h03 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h04 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h05 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h06 :
		rl_a06_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h07 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h08 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h09 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h0a :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h0b :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h0c :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h0d :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h0e :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h0f :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h10 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h11 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h12 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h13 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h14 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h15 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h16 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h17 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h18 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h19 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h1a :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h1b :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h1c :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h1d :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h1e :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h1f :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h20 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h21 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h22 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h23 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h24 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h25 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h26 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h27 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h28 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h29 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h2a :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h2b :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h2c :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h2d :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h2e :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h2f :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h30 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h31 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h32 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h33 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h34 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h35 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h36 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h37 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h38 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h39 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h3a :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h3b :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h3c :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h3d :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h3e :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h3f :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h40 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h41 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h42 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h43 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h44 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h45 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h46 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h47 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h48 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h49 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h4a :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h4b :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h4c :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h4d :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h4e :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h4f :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h50 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h51 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h52 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h53 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h54 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h55 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h56 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h57 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h58 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h59 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h5a :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h5b :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h5c :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h5d :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h5e :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h5f :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h60 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h61 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h62 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h63 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h64 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h65 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h66 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h67 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h68 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h69 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h6a :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h6b :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h6c :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h6d :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h6e :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h6f :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h70 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h71 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h72 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h73 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h74 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h75 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h76 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h77 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h78 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h79 :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h7a :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h7b :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h7c :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h7d :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h7e :
		rl_a06_t4_t1 = RG_rl_189 ;
	7'h7f :
		rl_a06_t4_t1 = RG_rl_189 ;
	default :
		rl_a06_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a06_t4_t1 or rl_a06_t5 or FF_i )
	begin
	rl_a06_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a06_t4 = ( ( { 9{ FF_i } } & rl_a06_t5 )
		| ( { 9{ rl_a06_t4_c1 } } & rl_a06_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_190 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h01 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h02 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h03 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h04 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h05 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h06 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h07 :
		rl_a07_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h08 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h09 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h0a :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h0b :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h0c :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h0d :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h0e :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h0f :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h10 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h11 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h12 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h13 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h14 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h15 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h16 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h17 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h18 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h19 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h1a :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h1b :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h1c :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h1d :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h1e :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h1f :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h20 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h21 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h22 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h23 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h24 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h25 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h26 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h27 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h28 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h29 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h2a :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h2b :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h2c :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h2d :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h2e :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h2f :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h30 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h31 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h32 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h33 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h34 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h35 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h36 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h37 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h38 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h39 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h3a :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h3b :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h3c :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h3d :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h3e :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h3f :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h40 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h41 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h42 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h43 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h44 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h45 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h46 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h47 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h48 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h49 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h4a :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h4b :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h4c :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h4d :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h4e :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h4f :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h50 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h51 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h52 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h53 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h54 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h55 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h56 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h57 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h58 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h59 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h5a :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h5b :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h5c :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h5d :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h5e :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h5f :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h60 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h61 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h62 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h63 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h64 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h65 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h66 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h67 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h68 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h69 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h6a :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h6b :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h6c :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h6d :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h6e :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h6f :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h70 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h71 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h72 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h73 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h74 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h75 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h76 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h77 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h78 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h79 :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h7a :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h7b :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h7c :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h7d :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h7e :
		rl_a07_t4_t1 = RG_rl_190 ;
	7'h7f :
		rl_a07_t4_t1 = RG_rl_190 ;
	default :
		rl_a07_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a07_t4_t1 or rl_a07_t5 or FF_i )
	begin
	rl_a07_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a07_t4 = ( ( { 9{ FF_i } } & rl_a07_t5 )
		| ( { 9{ rl_a07_t4_c1 } } & rl_a07_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_191 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h01 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h02 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h03 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h04 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h05 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h06 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h07 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h08 :
		rl_a08_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h09 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h0a :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h0b :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h0c :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h0d :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h0e :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h0f :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h10 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h11 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h12 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h13 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h14 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h15 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h16 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h17 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h18 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h19 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h1a :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h1b :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h1c :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h1d :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h1e :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h1f :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h20 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h21 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h22 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h23 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h24 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h25 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h26 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h27 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h28 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h29 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h2a :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h2b :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h2c :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h2d :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h2e :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h2f :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h30 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h31 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h32 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h33 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h34 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h35 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h36 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h37 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h38 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h39 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h3a :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h3b :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h3c :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h3d :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h3e :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h3f :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h40 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h41 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h42 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h43 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h44 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h45 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h46 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h47 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h48 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h49 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h4a :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h4b :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h4c :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h4d :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h4e :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h4f :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h50 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h51 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h52 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h53 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h54 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h55 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h56 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h57 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h58 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h59 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h5a :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h5b :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h5c :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h5d :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h5e :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h5f :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h60 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h61 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h62 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h63 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h64 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h65 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h66 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h67 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h68 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h69 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h6a :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h6b :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h6c :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h6d :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h6e :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h6f :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h70 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h71 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h72 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h73 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h74 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h75 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h76 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h77 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h78 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h79 :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h7a :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h7b :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h7c :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h7d :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h7e :
		rl_a08_t4_t1 = RG_rl_191 ;
	7'h7f :
		rl_a08_t4_t1 = RG_rl_191 ;
	default :
		rl_a08_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a08_t4_t1 or rl_a08_t5 or FF_i )
	begin
	rl_a08_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a08_t4 = ( ( { 9{ FF_i } } & rl_a08_t5 )
		| ( { 9{ rl_a08_t4_c1 } } & rl_a08_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_192 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h01 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h02 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h03 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h04 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h05 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h06 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h07 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h08 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h09 :
		rl_a09_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h0a :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h0b :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h0c :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h0d :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h0e :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h0f :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h10 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h11 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h12 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h13 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h14 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h15 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h16 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h17 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h18 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h19 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h1a :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h1b :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h1c :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h1d :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h1e :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h1f :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h20 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h21 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h22 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h23 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h24 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h25 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h26 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h27 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h28 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h29 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h2a :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h2b :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h2c :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h2d :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h2e :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h2f :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h30 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h31 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h32 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h33 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h34 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h35 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h36 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h37 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h38 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h39 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h3a :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h3b :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h3c :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h3d :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h3e :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h3f :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h40 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h41 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h42 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h43 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h44 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h45 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h46 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h47 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h48 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h49 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h4a :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h4b :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h4c :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h4d :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h4e :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h4f :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h50 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h51 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h52 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h53 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h54 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h55 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h56 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h57 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h58 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h59 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h5a :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h5b :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h5c :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h5d :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h5e :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h5f :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h60 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h61 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h62 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h63 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h64 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h65 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h66 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h67 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h68 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h69 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h6a :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h6b :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h6c :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h6d :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h6e :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h6f :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h70 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h71 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h72 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h73 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h74 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h75 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h76 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h77 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h78 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h79 :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h7a :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h7b :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h7c :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h7d :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h7e :
		rl_a09_t4_t1 = RG_rl_192 ;
	7'h7f :
		rl_a09_t4_t1 = RG_rl_192 ;
	default :
		rl_a09_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a09_t4_t1 or rl_a09_t5 or FF_i )
	begin
	rl_a09_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a09_t4 = ( ( { 9{ FF_i } } & rl_a09_t5 )
		| ( { 9{ rl_a09_t4_c1 } } & rl_a09_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_193 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h01 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h02 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h03 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h04 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h05 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h06 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h07 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h08 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h09 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h0a :
		rl_a10_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h0b :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h0c :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h0d :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h0e :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h0f :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h10 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h11 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h12 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h13 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h14 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h15 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h16 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h17 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h18 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h19 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h1a :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h1b :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h1c :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h1d :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h1e :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h1f :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h20 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h21 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h22 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h23 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h24 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h25 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h26 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h27 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h28 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h29 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h2a :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h2b :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h2c :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h2d :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h2e :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h2f :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h30 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h31 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h32 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h33 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h34 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h35 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h36 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h37 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h38 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h39 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h3a :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h3b :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h3c :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h3d :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h3e :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h3f :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h40 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h41 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h42 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h43 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h44 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h45 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h46 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h47 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h48 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h49 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h4a :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h4b :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h4c :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h4d :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h4e :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h4f :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h50 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h51 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h52 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h53 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h54 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h55 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h56 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h57 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h58 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h59 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h5a :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h5b :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h5c :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h5d :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h5e :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h5f :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h60 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h61 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h62 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h63 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h64 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h65 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h66 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h67 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h68 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h69 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h6a :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h6b :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h6c :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h6d :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h6e :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h6f :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h70 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h71 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h72 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h73 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h74 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h75 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h76 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h77 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h78 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h79 :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h7a :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h7b :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h7c :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h7d :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h7e :
		rl_a10_t4_t1 = RG_rl_193 ;
	7'h7f :
		rl_a10_t4_t1 = RG_rl_193 ;
	default :
		rl_a10_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a10_t4_t1 or rl_a10_t5 or FF_i )
	begin
	rl_a10_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a10_t4 = ( ( { 9{ FF_i } } & rl_a10_t5 )
		| ( { 9{ rl_a10_t4_c1 } } & rl_a10_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_194 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h01 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h02 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h03 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h04 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h05 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h06 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h07 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h08 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h09 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h0a :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h0b :
		rl_a11_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h0c :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h0d :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h0e :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h0f :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h10 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h11 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h12 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h13 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h14 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h15 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h16 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h17 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h18 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h19 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h1a :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h1b :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h1c :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h1d :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h1e :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h1f :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h20 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h21 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h22 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h23 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h24 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h25 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h26 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h27 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h28 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h29 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h2a :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h2b :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h2c :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h2d :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h2e :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h2f :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h30 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h31 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h32 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h33 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h34 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h35 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h36 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h37 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h38 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h39 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h3a :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h3b :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h3c :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h3d :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h3e :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h3f :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h40 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h41 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h42 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h43 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h44 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h45 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h46 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h47 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h48 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h49 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h4a :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h4b :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h4c :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h4d :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h4e :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h4f :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h50 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h51 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h52 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h53 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h54 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h55 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h56 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h57 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h58 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h59 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h5a :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h5b :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h5c :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h5d :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h5e :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h5f :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h60 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h61 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h62 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h63 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h64 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h65 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h66 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h67 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h68 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h69 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h6a :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h6b :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h6c :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h6d :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h6e :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h6f :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h70 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h71 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h72 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h73 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h74 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h75 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h76 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h77 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h78 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h79 :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h7a :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h7b :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h7c :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h7d :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h7e :
		rl_a11_t4_t1 = RG_rl_194 ;
	7'h7f :
		rl_a11_t4_t1 = RG_rl_194 ;
	default :
		rl_a11_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a11_t4_t1 or rl_a11_t5 or FF_i )
	begin
	rl_a11_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a11_t4 = ( ( { 9{ FF_i } } & rl_a11_t5 )
		| ( { 9{ rl_a11_t4_c1 } } & rl_a11_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_195 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h01 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h02 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h03 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h04 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h05 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h06 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h07 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h08 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h09 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h0a :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h0b :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h0c :
		rl_a12_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h0d :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h0e :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h0f :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h10 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h11 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h12 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h13 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h14 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h15 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h16 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h17 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h18 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h19 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h1a :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h1b :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h1c :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h1d :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h1e :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h1f :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h20 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h21 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h22 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h23 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h24 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h25 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h26 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h27 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h28 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h29 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h2a :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h2b :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h2c :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h2d :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h2e :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h2f :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h30 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h31 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h32 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h33 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h34 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h35 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h36 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h37 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h38 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h39 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h3a :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h3b :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h3c :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h3d :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h3e :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h3f :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h40 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h41 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h42 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h43 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h44 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h45 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h46 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h47 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h48 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h49 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h4a :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h4b :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h4c :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h4d :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h4e :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h4f :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h50 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h51 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h52 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h53 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h54 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h55 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h56 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h57 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h58 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h59 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h5a :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h5b :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h5c :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h5d :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h5e :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h5f :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h60 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h61 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h62 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h63 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h64 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h65 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h66 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h67 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h68 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h69 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h6a :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h6b :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h6c :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h6d :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h6e :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h6f :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h70 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h71 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h72 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h73 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h74 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h75 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h76 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h77 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h78 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h79 :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h7a :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h7b :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h7c :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h7d :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h7e :
		rl_a12_t4_t1 = RG_rl_195 ;
	7'h7f :
		rl_a12_t4_t1 = RG_rl_195 ;
	default :
		rl_a12_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a12_t4_t1 or rl_a12_t5 or FF_i )
	begin
	rl_a12_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a12_t4 = ( ( { 9{ FF_i } } & rl_a12_t5 )
		| ( { 9{ rl_a12_t4_c1 } } & rl_a12_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_196 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h01 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h02 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h03 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h04 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h05 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h06 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h07 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h08 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h09 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h0a :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h0b :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h0c :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h0d :
		rl_a13_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h0e :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h0f :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h10 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h11 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h12 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h13 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h14 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h15 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h16 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h17 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h18 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h19 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h1a :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h1b :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h1c :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h1d :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h1e :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h1f :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h20 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h21 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h22 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h23 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h24 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h25 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h26 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h27 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h28 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h29 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h2a :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h2b :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h2c :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h2d :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h2e :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h2f :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h30 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h31 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h32 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h33 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h34 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h35 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h36 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h37 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h38 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h39 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h3a :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h3b :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h3c :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h3d :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h3e :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h3f :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h40 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h41 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h42 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h43 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h44 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h45 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h46 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h47 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h48 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h49 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h4a :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h4b :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h4c :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h4d :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h4e :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h4f :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h50 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h51 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h52 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h53 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h54 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h55 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h56 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h57 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h58 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h59 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h5a :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h5b :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h5c :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h5d :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h5e :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h5f :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h60 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h61 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h62 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h63 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h64 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h65 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h66 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h67 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h68 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h69 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h6a :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h6b :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h6c :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h6d :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h6e :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h6f :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h70 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h71 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h72 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h73 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h74 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h75 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h76 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h77 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h78 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h79 :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h7a :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h7b :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h7c :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h7d :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h7e :
		rl_a13_t4_t1 = RG_rl_196 ;
	7'h7f :
		rl_a13_t4_t1 = RG_rl_196 ;
	default :
		rl_a13_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a13_t4_t1 or rl_a13_t5 or FF_i )
	begin
	rl_a13_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a13_t4 = ( ( { 9{ FF_i } } & rl_a13_t5 )
		| ( { 9{ rl_a13_t4_c1 } } & rl_a13_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_197 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h01 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h02 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h03 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h04 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h05 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h06 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h07 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h08 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h09 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h0a :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h0b :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h0c :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h0d :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h0e :
		rl_a14_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h0f :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h10 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h11 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h12 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h13 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h14 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h15 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h16 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h17 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h18 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h19 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h1a :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h1b :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h1c :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h1d :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h1e :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h1f :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h20 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h21 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h22 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h23 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h24 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h25 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h26 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h27 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h28 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h29 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h2a :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h2b :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h2c :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h2d :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h2e :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h2f :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h30 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h31 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h32 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h33 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h34 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h35 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h36 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h37 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h38 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h39 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h3a :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h3b :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h3c :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h3d :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h3e :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h3f :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h40 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h41 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h42 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h43 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h44 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h45 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h46 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h47 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h48 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h49 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h4a :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h4b :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h4c :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h4d :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h4e :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h4f :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h50 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h51 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h52 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h53 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h54 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h55 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h56 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h57 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h58 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h59 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h5a :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h5b :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h5c :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h5d :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h5e :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h5f :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h60 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h61 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h62 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h63 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h64 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h65 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h66 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h67 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h68 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h69 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h6a :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h6b :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h6c :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h6d :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h6e :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h6f :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h70 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h71 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h72 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h73 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h74 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h75 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h76 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h77 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h78 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h79 :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h7a :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h7b :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h7c :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h7d :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h7e :
		rl_a14_t4_t1 = RG_rl_197 ;
	7'h7f :
		rl_a14_t4_t1 = RG_rl_197 ;
	default :
		rl_a14_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a14_t4_t1 or rl_a14_t5 or FF_i )
	begin
	rl_a14_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a14_t4 = ( ( { 9{ FF_i } } & rl_a14_t5 )
		| ( { 9{ rl_a14_t4_c1 } } & rl_a14_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_198 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h01 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h02 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h03 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h04 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h05 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h06 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h07 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h08 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h09 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h0a :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h0b :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h0c :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h0d :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h0e :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h0f :
		rl_a15_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h10 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h11 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h12 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h13 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h14 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h15 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h16 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h17 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h18 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h19 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h1a :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h1b :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h1c :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h1d :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h1e :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h1f :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h20 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h21 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h22 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h23 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h24 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h25 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h26 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h27 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h28 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h29 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h2a :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h2b :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h2c :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h2d :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h2e :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h2f :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h30 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h31 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h32 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h33 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h34 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h35 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h36 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h37 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h38 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h39 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h3a :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h3b :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h3c :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h3d :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h3e :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h3f :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h40 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h41 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h42 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h43 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h44 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h45 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h46 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h47 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h48 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h49 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h4a :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h4b :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h4c :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h4d :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h4e :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h4f :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h50 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h51 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h52 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h53 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h54 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h55 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h56 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h57 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h58 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h59 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h5a :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h5b :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h5c :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h5d :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h5e :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h5f :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h60 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h61 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h62 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h63 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h64 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h65 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h66 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h67 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h68 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h69 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h6a :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h6b :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h6c :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h6d :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h6e :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h6f :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h70 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h71 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h72 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h73 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h74 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h75 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h76 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h77 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h78 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h79 :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h7a :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h7b :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h7c :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h7d :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h7e :
		rl_a15_t4_t1 = RG_rl_198 ;
	7'h7f :
		rl_a15_t4_t1 = RG_rl_198 ;
	default :
		rl_a15_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a15_t4_t1 or rl_a15_t5 or FF_i )
	begin
	rl_a15_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a15_t4 = ( ( { 9{ FF_i } } & rl_a15_t5 )
		| ( { 9{ rl_a15_t4_c1 } } & rl_a15_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_199 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h01 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h02 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h03 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h04 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h05 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h06 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h07 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h08 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h09 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h0a :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h0b :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h0c :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h0d :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h0e :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h0f :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h10 :
		rl_a16_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h11 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h12 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h13 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h14 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h15 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h16 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h17 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h18 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h19 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h1a :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h1b :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h1c :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h1d :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h1e :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h1f :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h20 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h21 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h22 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h23 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h24 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h25 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h26 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h27 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h28 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h29 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h2a :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h2b :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h2c :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h2d :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h2e :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h2f :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h30 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h31 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h32 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h33 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h34 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h35 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h36 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h37 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h38 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h39 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h3a :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h3b :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h3c :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h3d :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h3e :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h3f :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h40 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h41 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h42 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h43 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h44 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h45 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h46 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h47 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h48 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h49 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h4a :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h4b :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h4c :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h4d :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h4e :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h4f :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h50 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h51 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h52 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h53 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h54 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h55 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h56 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h57 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h58 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h59 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h5a :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h5b :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h5c :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h5d :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h5e :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h5f :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h60 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h61 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h62 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h63 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h64 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h65 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h66 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h67 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h68 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h69 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h6a :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h6b :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h6c :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h6d :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h6e :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h6f :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h70 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h71 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h72 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h73 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h74 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h75 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h76 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h77 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h78 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h79 :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h7a :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h7b :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h7c :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h7d :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h7e :
		rl_a16_t4_t1 = RG_rl_199 ;
	7'h7f :
		rl_a16_t4_t1 = RG_rl_199 ;
	default :
		rl_a16_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a16_t4_t1 or rl_a16_t5 or FF_i )
	begin
	rl_a16_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a16_t4 = ( ( { 9{ FF_i } } & rl_a16_t5 )
		| ( { 9{ rl_a16_t4_c1 } } & rl_a16_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_200 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h01 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h02 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h03 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h04 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h05 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h06 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h07 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h08 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h09 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h0a :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h0b :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h0c :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h0d :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h0e :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h0f :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h10 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h11 :
		rl_a17_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h12 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h13 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h14 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h15 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h16 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h17 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h18 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h19 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h1a :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h1b :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h1c :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h1d :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h1e :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h1f :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h20 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h21 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h22 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h23 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h24 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h25 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h26 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h27 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h28 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h29 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h2a :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h2b :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h2c :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h2d :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h2e :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h2f :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h30 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h31 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h32 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h33 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h34 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h35 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h36 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h37 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h38 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h39 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h3a :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h3b :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h3c :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h3d :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h3e :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h3f :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h40 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h41 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h42 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h43 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h44 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h45 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h46 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h47 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h48 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h49 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h4a :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h4b :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h4c :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h4d :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h4e :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h4f :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h50 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h51 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h52 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h53 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h54 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h55 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h56 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h57 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h58 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h59 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h5a :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h5b :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h5c :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h5d :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h5e :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h5f :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h60 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h61 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h62 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h63 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h64 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h65 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h66 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h67 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h68 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h69 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h6a :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h6b :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h6c :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h6d :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h6e :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h6f :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h70 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h71 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h72 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h73 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h74 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h75 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h76 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h77 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h78 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h79 :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h7a :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h7b :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h7c :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h7d :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h7e :
		rl_a17_t4_t1 = RG_rl_200 ;
	7'h7f :
		rl_a17_t4_t1 = RG_rl_200 ;
	default :
		rl_a17_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a17_t4_t1 or rl_a17_t5 or FF_i )
	begin
	rl_a17_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a17_t4 = ( ( { 9{ FF_i } } & rl_a17_t5 )
		| ( { 9{ rl_a17_t4_c1 } } & rl_a17_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_201 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h01 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h02 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h03 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h04 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h05 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h06 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h07 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h08 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h09 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h0a :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h0b :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h0c :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h0d :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h0e :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h0f :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h10 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h11 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h12 :
		rl_a18_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h13 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h14 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h15 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h16 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h17 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h18 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h19 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h1a :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h1b :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h1c :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h1d :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h1e :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h1f :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h20 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h21 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h22 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h23 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h24 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h25 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h26 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h27 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h28 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h29 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h2a :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h2b :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h2c :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h2d :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h2e :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h2f :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h30 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h31 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h32 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h33 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h34 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h35 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h36 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h37 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h38 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h39 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h3a :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h3b :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h3c :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h3d :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h3e :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h3f :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h40 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h41 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h42 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h43 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h44 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h45 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h46 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h47 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h48 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h49 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h4a :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h4b :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h4c :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h4d :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h4e :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h4f :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h50 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h51 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h52 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h53 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h54 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h55 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h56 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h57 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h58 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h59 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h5a :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h5b :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h5c :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h5d :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h5e :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h5f :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h60 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h61 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h62 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h63 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h64 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h65 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h66 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h67 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h68 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h69 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h6a :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h6b :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h6c :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h6d :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h6e :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h6f :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h70 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h71 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h72 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h73 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h74 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h75 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h76 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h77 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h78 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h79 :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h7a :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h7b :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h7c :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h7d :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h7e :
		rl_a18_t4_t1 = RG_rl_201 ;
	7'h7f :
		rl_a18_t4_t1 = RG_rl_201 ;
	default :
		rl_a18_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a18_t4_t1 or rl_a18_t5 or FF_i )
	begin
	rl_a18_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a18_t4 = ( ( { 9{ FF_i } } & rl_a18_t5 )
		| ( { 9{ rl_a18_t4_c1 } } & rl_a18_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_202 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h01 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h02 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h03 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h04 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h05 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h06 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h07 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h08 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h09 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h0a :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h0b :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h0c :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h0d :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h0e :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h0f :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h10 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h11 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h12 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h13 :
		rl_a19_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h14 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h15 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h16 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h17 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h18 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h19 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h1a :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h1b :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h1c :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h1d :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h1e :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h1f :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h20 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h21 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h22 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h23 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h24 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h25 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h26 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h27 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h28 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h29 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h2a :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h2b :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h2c :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h2d :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h2e :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h2f :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h30 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h31 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h32 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h33 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h34 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h35 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h36 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h37 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h38 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h39 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h3a :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h3b :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h3c :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h3d :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h3e :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h3f :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h40 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h41 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h42 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h43 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h44 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h45 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h46 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h47 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h48 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h49 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h4a :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h4b :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h4c :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h4d :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h4e :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h4f :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h50 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h51 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h52 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h53 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h54 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h55 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h56 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h57 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h58 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h59 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h5a :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h5b :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h5c :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h5d :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h5e :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h5f :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h60 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h61 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h62 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h63 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h64 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h65 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h66 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h67 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h68 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h69 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h6a :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h6b :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h6c :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h6d :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h6e :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h6f :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h70 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h71 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h72 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h73 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h74 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h75 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h76 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h77 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h78 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h79 :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h7a :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h7b :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h7c :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h7d :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h7e :
		rl_a19_t4_t1 = RG_rl_202 ;
	7'h7f :
		rl_a19_t4_t1 = RG_rl_202 ;
	default :
		rl_a19_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a19_t4_t1 or rl_a19_t5 or FF_i )
	begin
	rl_a19_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a19_t4 = ( ( { 9{ FF_i } } & rl_a19_t5 )
		| ( { 9{ rl_a19_t4_c1 } } & rl_a19_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_203 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h01 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h02 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h03 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h04 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h05 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h06 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h07 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h08 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h09 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h0a :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h0b :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h0c :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h0d :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h0e :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h0f :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h10 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h11 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h12 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h13 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h14 :
		rl_a20_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h15 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h16 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h17 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h18 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h19 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h1a :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h1b :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h1c :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h1d :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h1e :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h1f :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h20 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h21 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h22 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h23 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h24 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h25 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h26 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h27 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h28 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h29 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h2a :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h2b :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h2c :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h2d :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h2e :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h2f :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h30 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h31 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h32 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h33 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h34 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h35 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h36 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h37 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h38 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h39 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h3a :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h3b :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h3c :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h3d :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h3e :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h3f :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h40 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h41 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h42 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h43 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h44 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h45 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h46 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h47 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h48 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h49 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h4a :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h4b :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h4c :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h4d :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h4e :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h4f :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h50 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h51 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h52 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h53 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h54 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h55 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h56 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h57 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h58 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h59 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h5a :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h5b :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h5c :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h5d :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h5e :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h5f :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h60 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h61 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h62 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h63 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h64 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h65 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h66 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h67 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h68 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h69 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h6a :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h6b :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h6c :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h6d :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h6e :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h6f :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h70 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h71 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h72 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h73 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h74 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h75 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h76 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h77 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h78 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h79 :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h7a :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h7b :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h7c :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h7d :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h7e :
		rl_a20_t4_t1 = RG_rl_203 ;
	7'h7f :
		rl_a20_t4_t1 = RG_rl_203 ;
	default :
		rl_a20_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a20_t4_t1 or rl_a20_t5 or FF_i )
	begin
	rl_a20_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a20_t4 = ( ( { 9{ FF_i } } & rl_a20_t5 )
		| ( { 9{ rl_a20_t4_c1 } } & rl_a20_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_204 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h01 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h02 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h03 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h04 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h05 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h06 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h07 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h08 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h09 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h0a :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h0b :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h0c :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h0d :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h0e :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h0f :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h10 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h11 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h12 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h13 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h14 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h15 :
		rl_a21_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h16 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h17 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h18 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h19 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h1a :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h1b :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h1c :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h1d :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h1e :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h1f :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h20 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h21 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h22 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h23 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h24 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h25 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h26 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h27 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h28 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h29 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h2a :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h2b :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h2c :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h2d :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h2e :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h2f :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h30 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h31 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h32 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h33 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h34 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h35 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h36 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h37 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h38 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h39 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h3a :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h3b :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h3c :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h3d :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h3e :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h3f :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h40 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h41 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h42 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h43 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h44 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h45 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h46 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h47 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h48 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h49 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h4a :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h4b :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h4c :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h4d :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h4e :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h4f :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h50 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h51 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h52 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h53 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h54 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h55 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h56 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h57 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h58 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h59 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h5a :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h5b :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h5c :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h5d :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h5e :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h5f :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h60 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h61 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h62 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h63 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h64 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h65 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h66 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h67 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h68 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h69 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h6a :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h6b :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h6c :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h6d :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h6e :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h6f :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h70 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h71 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h72 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h73 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h74 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h75 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h76 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h77 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h78 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h79 :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h7a :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h7b :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h7c :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h7d :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h7e :
		rl_a21_t4_t1 = RG_rl_204 ;
	7'h7f :
		rl_a21_t4_t1 = RG_rl_204 ;
	default :
		rl_a21_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a21_t4_t1 or rl_a21_t5 or FF_i )
	begin
	rl_a21_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a21_t4 = ( ( { 9{ FF_i } } & rl_a21_t5 )
		| ( { 9{ rl_a21_t4_c1 } } & rl_a21_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_205 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h01 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h02 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h03 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h04 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h05 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h06 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h07 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h08 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h09 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h0a :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h0b :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h0c :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h0d :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h0e :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h0f :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h10 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h11 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h12 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h13 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h14 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h15 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h16 :
		rl_a22_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h17 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h18 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h19 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h1a :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h1b :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h1c :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h1d :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h1e :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h1f :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h20 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h21 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h22 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h23 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h24 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h25 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h26 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h27 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h28 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h29 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h2a :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h2b :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h2c :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h2d :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h2e :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h2f :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h30 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h31 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h32 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h33 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h34 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h35 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h36 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h37 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h38 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h39 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h3a :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h3b :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h3c :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h3d :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h3e :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h3f :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h40 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h41 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h42 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h43 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h44 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h45 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h46 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h47 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h48 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h49 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h4a :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h4b :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h4c :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h4d :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h4e :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h4f :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h50 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h51 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h52 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h53 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h54 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h55 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h56 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h57 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h58 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h59 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h5a :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h5b :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h5c :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h5d :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h5e :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h5f :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h60 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h61 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h62 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h63 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h64 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h65 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h66 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h67 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h68 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h69 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h6a :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h6b :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h6c :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h6d :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h6e :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h6f :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h70 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h71 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h72 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h73 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h74 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h75 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h76 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h77 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h78 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h79 :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h7a :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h7b :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h7c :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h7d :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h7e :
		rl_a22_t4_t1 = RG_rl_205 ;
	7'h7f :
		rl_a22_t4_t1 = RG_rl_205 ;
	default :
		rl_a22_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a22_t4_t1 or rl_a22_t5 or FF_i )
	begin
	rl_a22_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a22_t4 = ( ( { 9{ FF_i } } & rl_a22_t5 )
		| ( { 9{ rl_a22_t4_c1 } } & rl_a22_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_206 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h01 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h02 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h03 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h04 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h05 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h06 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h07 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h08 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h09 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h0a :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h0b :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h0c :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h0d :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h0e :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h0f :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h10 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h11 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h12 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h13 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h14 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h15 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h16 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h17 :
		rl_a23_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h18 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h19 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h1a :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h1b :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h1c :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h1d :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h1e :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h1f :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h20 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h21 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h22 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h23 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h24 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h25 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h26 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h27 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h28 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h29 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h2a :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h2b :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h2c :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h2d :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h2e :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h2f :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h30 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h31 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h32 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h33 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h34 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h35 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h36 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h37 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h38 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h39 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h3a :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h3b :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h3c :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h3d :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h3e :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h3f :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h40 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h41 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h42 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h43 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h44 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h45 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h46 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h47 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h48 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h49 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h4a :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h4b :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h4c :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h4d :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h4e :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h4f :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h50 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h51 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h52 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h53 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h54 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h55 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h56 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h57 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h58 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h59 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h5a :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h5b :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h5c :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h5d :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h5e :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h5f :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h60 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h61 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h62 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h63 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h64 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h65 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h66 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h67 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h68 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h69 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h6a :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h6b :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h6c :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h6d :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h6e :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h6f :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h70 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h71 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h72 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h73 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h74 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h75 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h76 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h77 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h78 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h79 :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h7a :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h7b :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h7c :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h7d :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h7e :
		rl_a23_t4_t1 = RG_rl_206 ;
	7'h7f :
		rl_a23_t4_t1 = RG_rl_206 ;
	default :
		rl_a23_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a23_t4_t1 or rl_a23_t5 or FF_i )
	begin
	rl_a23_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a23_t4 = ( ( { 9{ FF_i } } & rl_a23_t5 )
		| ( { 9{ rl_a23_t4_c1 } } & rl_a23_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_207 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h01 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h02 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h03 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h04 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h05 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h06 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h07 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h08 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h09 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h0a :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h0b :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h0c :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h0d :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h0e :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h0f :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h10 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h11 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h12 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h13 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h14 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h15 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h16 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h17 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h18 :
		rl_a24_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h19 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h1a :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h1b :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h1c :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h1d :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h1e :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h1f :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h20 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h21 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h22 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h23 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h24 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h25 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h26 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h27 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h28 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h29 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h2a :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h2b :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h2c :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h2d :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h2e :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h2f :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h30 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h31 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h32 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h33 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h34 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h35 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h36 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h37 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h38 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h39 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h3a :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h3b :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h3c :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h3d :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h3e :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h3f :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h40 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h41 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h42 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h43 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h44 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h45 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h46 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h47 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h48 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h49 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h4a :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h4b :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h4c :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h4d :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h4e :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h4f :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h50 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h51 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h52 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h53 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h54 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h55 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h56 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h57 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h58 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h59 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h5a :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h5b :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h5c :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h5d :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h5e :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h5f :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h60 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h61 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h62 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h63 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h64 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h65 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h66 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h67 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h68 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h69 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h6a :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h6b :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h6c :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h6d :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h6e :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h6f :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h70 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h71 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h72 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h73 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h74 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h75 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h76 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h77 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h78 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h79 :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h7a :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h7b :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h7c :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h7d :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h7e :
		rl_a24_t4_t1 = RG_rl_207 ;
	7'h7f :
		rl_a24_t4_t1 = RG_rl_207 ;
	default :
		rl_a24_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a24_t4_t1 or rl_a24_t5 or FF_i )
	begin
	rl_a24_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a24_t4 = ( ( { 9{ FF_i } } & rl_a24_t5 )
		| ( { 9{ rl_a24_t4_c1 } } & rl_a24_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_208 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h01 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h02 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h03 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h04 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h05 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h06 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h07 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h08 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h09 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h0a :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h0b :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h0c :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h0d :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h0e :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h0f :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h10 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h11 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h12 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h13 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h14 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h15 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h16 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h17 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h18 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h19 :
		rl_a25_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h1a :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h1b :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h1c :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h1d :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h1e :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h1f :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h20 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h21 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h22 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h23 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h24 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h25 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h26 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h27 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h28 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h29 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h2a :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h2b :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h2c :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h2d :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h2e :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h2f :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h30 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h31 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h32 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h33 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h34 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h35 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h36 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h37 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h38 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h39 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h3a :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h3b :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h3c :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h3d :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h3e :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h3f :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h40 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h41 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h42 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h43 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h44 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h45 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h46 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h47 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h48 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h49 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h4a :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h4b :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h4c :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h4d :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h4e :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h4f :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h50 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h51 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h52 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h53 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h54 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h55 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h56 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h57 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h58 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h59 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h5a :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h5b :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h5c :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h5d :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h5e :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h5f :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h60 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h61 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h62 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h63 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h64 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h65 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h66 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h67 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h68 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h69 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h6a :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h6b :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h6c :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h6d :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h6e :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h6f :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h70 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h71 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h72 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h73 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h74 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h75 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h76 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h77 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h78 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h79 :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h7a :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h7b :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h7c :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h7d :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h7e :
		rl_a25_t4_t1 = RG_rl_208 ;
	7'h7f :
		rl_a25_t4_t1 = RG_rl_208 ;
	default :
		rl_a25_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a25_t4_t1 or rl_a25_t5 or FF_i )
	begin
	rl_a25_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a25_t4 = ( ( { 9{ FF_i } } & rl_a25_t5 )
		| ( { 9{ rl_a25_t4_c1 } } & rl_a25_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_209 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h01 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h02 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h03 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h04 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h05 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h06 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h07 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h08 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h09 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h0a :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h0b :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h0c :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h0d :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h0e :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h0f :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h10 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h11 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h12 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h13 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h14 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h15 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h16 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h17 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h18 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h19 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h1a :
		rl_a26_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h1b :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h1c :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h1d :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h1e :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h1f :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h20 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h21 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h22 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h23 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h24 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h25 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h26 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h27 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h28 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h29 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h2a :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h2b :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h2c :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h2d :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h2e :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h2f :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h30 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h31 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h32 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h33 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h34 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h35 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h36 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h37 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h38 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h39 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h3a :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h3b :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h3c :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h3d :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h3e :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h3f :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h40 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h41 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h42 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h43 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h44 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h45 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h46 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h47 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h48 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h49 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h4a :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h4b :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h4c :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h4d :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h4e :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h4f :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h50 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h51 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h52 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h53 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h54 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h55 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h56 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h57 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h58 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h59 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h5a :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h5b :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h5c :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h5d :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h5e :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h5f :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h60 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h61 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h62 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h63 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h64 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h65 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h66 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h67 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h68 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h69 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h6a :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h6b :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h6c :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h6d :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h6e :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h6f :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h70 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h71 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h72 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h73 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h74 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h75 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h76 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h77 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h78 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h79 :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h7a :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h7b :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h7c :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h7d :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h7e :
		rl_a26_t4_t1 = RG_rl_209 ;
	7'h7f :
		rl_a26_t4_t1 = RG_rl_209 ;
	default :
		rl_a26_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a26_t4_t1 or rl_a26_t5 or FF_i )
	begin
	rl_a26_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a26_t4 = ( ( { 9{ FF_i } } & rl_a26_t5 )
		| ( { 9{ rl_a26_t4_c1 } } & rl_a26_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_210 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h01 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h02 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h03 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h04 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h05 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h06 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h07 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h08 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h09 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h0a :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h0b :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h0c :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h0d :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h0e :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h0f :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h10 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h11 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h12 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h13 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h14 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h15 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h16 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h17 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h18 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h19 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h1a :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h1b :
		rl_a27_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h1c :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h1d :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h1e :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h1f :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h20 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h21 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h22 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h23 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h24 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h25 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h26 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h27 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h28 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h29 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h2a :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h2b :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h2c :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h2d :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h2e :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h2f :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h30 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h31 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h32 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h33 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h34 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h35 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h36 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h37 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h38 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h39 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h3a :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h3b :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h3c :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h3d :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h3e :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h3f :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h40 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h41 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h42 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h43 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h44 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h45 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h46 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h47 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h48 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h49 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h4a :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h4b :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h4c :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h4d :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h4e :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h4f :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h50 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h51 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h52 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h53 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h54 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h55 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h56 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h57 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h58 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h59 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h5a :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h5b :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h5c :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h5d :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h5e :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h5f :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h60 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h61 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h62 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h63 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h64 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h65 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h66 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h67 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h68 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h69 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h6a :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h6b :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h6c :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h6d :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h6e :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h6f :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h70 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h71 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h72 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h73 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h74 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h75 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h76 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h77 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h78 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h79 :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h7a :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h7b :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h7c :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h7d :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h7e :
		rl_a27_t4_t1 = RG_rl_210 ;
	7'h7f :
		rl_a27_t4_t1 = RG_rl_210 ;
	default :
		rl_a27_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a27_t4_t1 or rl_a27_t5 or FF_i )
	begin
	rl_a27_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a27_t4 = ( ( { 9{ FF_i } } & rl_a27_t5 )
		| ( { 9{ rl_a27_t4_c1 } } & rl_a27_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_211 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h01 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h02 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h03 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h04 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h05 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h06 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h07 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h08 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h09 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h0a :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h0b :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h0c :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h0d :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h0e :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h0f :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h10 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h11 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h12 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h13 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h14 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h15 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h16 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h17 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h18 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h19 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h1a :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h1b :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h1c :
		rl_a28_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h1d :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h1e :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h1f :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h20 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h21 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h22 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h23 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h24 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h25 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h26 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h27 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h28 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h29 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h2a :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h2b :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h2c :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h2d :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h2e :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h2f :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h30 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h31 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h32 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h33 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h34 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h35 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h36 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h37 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h38 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h39 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h3a :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h3b :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h3c :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h3d :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h3e :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h3f :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h40 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h41 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h42 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h43 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h44 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h45 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h46 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h47 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h48 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h49 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h4a :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h4b :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h4c :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h4d :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h4e :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h4f :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h50 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h51 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h52 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h53 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h54 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h55 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h56 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h57 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h58 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h59 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h5a :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h5b :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h5c :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h5d :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h5e :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h5f :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h60 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h61 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h62 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h63 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h64 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h65 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h66 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h67 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h68 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h69 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h6a :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h6b :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h6c :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h6d :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h6e :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h6f :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h70 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h71 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h72 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h73 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h74 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h75 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h76 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h77 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h78 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h79 :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h7a :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h7b :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h7c :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h7d :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h7e :
		rl_a28_t4_t1 = RG_rl_211 ;
	7'h7f :
		rl_a28_t4_t1 = RG_rl_211 ;
	default :
		rl_a28_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a28_t4_t1 or rl_a28_t5 or FF_i )
	begin
	rl_a28_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a28_t4 = ( ( { 9{ FF_i } } & rl_a28_t5 )
		| ( { 9{ rl_a28_t4_c1 } } & rl_a28_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_212 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h01 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h02 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h03 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h04 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h05 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h06 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h07 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h08 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h09 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h0a :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h0b :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h0c :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h0d :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h0e :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h0f :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h10 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h11 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h12 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h13 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h14 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h15 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h16 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h17 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h18 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h19 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h1a :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h1b :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h1c :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h1d :
		rl_a29_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h1e :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h1f :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h20 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h21 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h22 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h23 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h24 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h25 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h26 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h27 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h28 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h29 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h2a :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h2b :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h2c :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h2d :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h2e :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h2f :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h30 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h31 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h32 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h33 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h34 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h35 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h36 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h37 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h38 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h39 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h3a :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h3b :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h3c :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h3d :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h3e :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h3f :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h40 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h41 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h42 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h43 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h44 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h45 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h46 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h47 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h48 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h49 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h4a :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h4b :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h4c :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h4d :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h4e :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h4f :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h50 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h51 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h52 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h53 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h54 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h55 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h56 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h57 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h58 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h59 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h5a :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h5b :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h5c :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h5d :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h5e :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h5f :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h60 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h61 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h62 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h63 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h64 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h65 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h66 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h67 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h68 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h69 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h6a :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h6b :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h6c :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h6d :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h6e :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h6f :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h70 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h71 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h72 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h73 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h74 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h75 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h76 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h77 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h78 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h79 :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h7a :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h7b :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h7c :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h7d :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h7e :
		rl_a29_t4_t1 = RG_rl_212 ;
	7'h7f :
		rl_a29_t4_t1 = RG_rl_212 ;
	default :
		rl_a29_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a29_t4_t1 or rl_a29_t5 or FF_i )
	begin
	rl_a29_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a29_t4 = ( ( { 9{ FF_i } } & rl_a29_t5 )
		| ( { 9{ rl_a29_t4_c1 } } & rl_a29_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_213 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h01 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h02 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h03 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h04 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h05 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h06 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h07 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h08 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h09 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h0a :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h0b :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h0c :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h0d :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h0e :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h0f :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h10 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h11 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h12 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h13 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h14 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h15 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h16 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h17 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h18 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h19 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h1a :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h1b :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h1c :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h1d :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h1e :
		rl_a30_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h1f :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h20 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h21 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h22 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h23 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h24 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h25 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h26 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h27 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h28 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h29 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h2a :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h2b :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h2c :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h2d :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h2e :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h2f :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h30 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h31 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h32 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h33 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h34 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h35 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h36 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h37 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h38 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h39 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h3a :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h3b :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h3c :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h3d :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h3e :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h3f :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h40 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h41 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h42 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h43 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h44 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h45 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h46 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h47 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h48 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h49 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h4a :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h4b :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h4c :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h4d :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h4e :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h4f :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h50 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h51 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h52 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h53 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h54 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h55 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h56 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h57 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h58 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h59 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h5a :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h5b :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h5c :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h5d :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h5e :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h5f :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h60 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h61 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h62 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h63 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h64 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h65 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h66 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h67 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h68 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h69 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h6a :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h6b :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h6c :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h6d :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h6e :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h6f :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h70 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h71 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h72 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h73 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h74 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h75 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h76 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h77 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h78 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h79 :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h7a :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h7b :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h7c :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h7d :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h7e :
		rl_a30_t4_t1 = RG_rl_213 ;
	7'h7f :
		rl_a30_t4_t1 = RG_rl_213 ;
	default :
		rl_a30_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a30_t4_t1 or rl_a30_t5 or FF_i )
	begin
	rl_a30_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a30_t4 = ( ( { 9{ FF_i } } & rl_a30_t5 )
		| ( { 9{ rl_a30_t4_c1 } } & rl_a30_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_214 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h01 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h02 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h03 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h04 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h05 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h06 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h07 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h08 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h09 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h0a :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h0b :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h0c :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h0d :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h0e :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h0f :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h10 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h11 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h12 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h13 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h14 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h15 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h16 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h17 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h18 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h19 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h1a :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h1b :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h1c :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h1d :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h1e :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h1f :
		rl_a31_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h20 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h21 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h22 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h23 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h24 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h25 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h26 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h27 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h28 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h29 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h2a :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h2b :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h2c :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h2d :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h2e :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h2f :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h30 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h31 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h32 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h33 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h34 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h35 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h36 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h37 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h38 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h39 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h3a :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h3b :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h3c :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h3d :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h3e :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h3f :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h40 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h41 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h42 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h43 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h44 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h45 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h46 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h47 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h48 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h49 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h4a :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h4b :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h4c :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h4d :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h4e :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h4f :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h50 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h51 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h52 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h53 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h54 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h55 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h56 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h57 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h58 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h59 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h5a :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h5b :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h5c :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h5d :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h5e :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h5f :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h60 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h61 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h62 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h63 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h64 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h65 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h66 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h67 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h68 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h69 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h6a :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h6b :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h6c :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h6d :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h6e :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h6f :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h70 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h71 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h72 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h73 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h74 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h75 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h76 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h77 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h78 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h79 :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h7a :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h7b :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h7c :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h7d :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h7e :
		rl_a31_t4_t1 = RG_rl_214 ;
	7'h7f :
		rl_a31_t4_t1 = RG_rl_214 ;
	default :
		rl_a31_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a31_t4_t1 or rl_a31_t5 or FF_i )
	begin
	rl_a31_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a31_t4 = ( ( { 9{ FF_i } } & rl_a31_t5 )
		| ( { 9{ rl_a31_t4_c1 } } & rl_a31_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_215 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h01 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h02 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h03 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h04 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h05 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h06 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h07 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h08 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h09 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h0a :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h0b :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h0c :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h0d :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h0e :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h0f :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h10 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h11 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h12 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h13 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h14 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h15 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h16 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h17 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h18 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h19 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h1a :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h1b :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h1c :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h1d :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h1e :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h1f :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h20 :
		rl_a32_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h21 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h22 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h23 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h24 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h25 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h26 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h27 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h28 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h29 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h2a :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h2b :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h2c :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h2d :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h2e :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h2f :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h30 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h31 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h32 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h33 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h34 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h35 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h36 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h37 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h38 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h39 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h3a :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h3b :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h3c :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h3d :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h3e :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h3f :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h40 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h41 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h42 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h43 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h44 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h45 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h46 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h47 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h48 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h49 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h4a :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h4b :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h4c :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h4d :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h4e :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h4f :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h50 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h51 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h52 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h53 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h54 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h55 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h56 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h57 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h58 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h59 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h5a :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h5b :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h5c :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h5d :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h5e :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h5f :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h60 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h61 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h62 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h63 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h64 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h65 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h66 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h67 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h68 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h69 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h6a :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h6b :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h6c :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h6d :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h6e :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h6f :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h70 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h71 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h72 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h73 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h74 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h75 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h76 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h77 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h78 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h79 :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h7a :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h7b :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h7c :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h7d :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h7e :
		rl_a32_t4_t1 = RG_rl_215 ;
	7'h7f :
		rl_a32_t4_t1 = RG_rl_215 ;
	default :
		rl_a32_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a32_t4_t1 or rl_a32_t5 or FF_i )
	begin
	rl_a32_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a32_t4 = ( ( { 9{ FF_i } } & rl_a32_t5 )
		| ( { 9{ rl_a32_t4_c1 } } & rl_a32_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_216 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h01 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h02 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h03 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h04 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h05 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h06 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h07 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h08 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h09 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h0a :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h0b :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h0c :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h0d :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h0e :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h0f :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h10 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h11 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h12 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h13 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h14 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h15 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h16 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h17 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h18 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h19 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h1a :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h1b :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h1c :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h1d :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h1e :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h1f :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h20 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h21 :
		rl_a33_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h22 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h23 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h24 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h25 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h26 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h27 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h28 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h29 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h2a :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h2b :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h2c :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h2d :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h2e :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h2f :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h30 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h31 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h32 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h33 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h34 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h35 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h36 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h37 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h38 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h39 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h3a :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h3b :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h3c :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h3d :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h3e :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h3f :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h40 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h41 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h42 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h43 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h44 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h45 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h46 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h47 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h48 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h49 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h4a :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h4b :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h4c :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h4d :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h4e :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h4f :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h50 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h51 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h52 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h53 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h54 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h55 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h56 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h57 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h58 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h59 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h5a :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h5b :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h5c :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h5d :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h5e :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h5f :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h60 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h61 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h62 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h63 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h64 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h65 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h66 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h67 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h68 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h69 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h6a :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h6b :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h6c :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h6d :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h6e :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h6f :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h70 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h71 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h72 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h73 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h74 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h75 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h76 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h77 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h78 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h79 :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h7a :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h7b :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h7c :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h7d :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h7e :
		rl_a33_t4_t1 = RG_rl_216 ;
	7'h7f :
		rl_a33_t4_t1 = RG_rl_216 ;
	default :
		rl_a33_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a33_t4_t1 or rl_a33_t5 or FF_i )
	begin
	rl_a33_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a33_t4 = ( ( { 9{ FF_i } } & rl_a33_t5 )
		| ( { 9{ rl_a33_t4_c1 } } & rl_a33_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_217 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h01 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h02 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h03 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h04 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h05 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h06 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h07 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h08 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h09 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h0a :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h0b :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h0c :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h0d :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h0e :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h0f :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h10 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h11 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h12 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h13 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h14 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h15 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h16 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h17 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h18 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h19 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h1a :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h1b :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h1c :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h1d :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h1e :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h1f :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h20 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h21 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h22 :
		rl_a34_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h23 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h24 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h25 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h26 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h27 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h28 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h29 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h2a :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h2b :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h2c :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h2d :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h2e :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h2f :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h30 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h31 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h32 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h33 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h34 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h35 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h36 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h37 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h38 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h39 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h3a :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h3b :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h3c :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h3d :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h3e :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h3f :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h40 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h41 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h42 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h43 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h44 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h45 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h46 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h47 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h48 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h49 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h4a :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h4b :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h4c :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h4d :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h4e :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h4f :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h50 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h51 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h52 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h53 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h54 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h55 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h56 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h57 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h58 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h59 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h5a :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h5b :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h5c :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h5d :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h5e :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h5f :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h60 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h61 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h62 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h63 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h64 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h65 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h66 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h67 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h68 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h69 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h6a :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h6b :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h6c :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h6d :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h6e :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h6f :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h70 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h71 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h72 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h73 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h74 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h75 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h76 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h77 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h78 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h79 :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h7a :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h7b :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h7c :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h7d :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h7e :
		rl_a34_t4_t1 = RG_rl_217 ;
	7'h7f :
		rl_a34_t4_t1 = RG_rl_217 ;
	default :
		rl_a34_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a34_t4_t1 or rl_a34_t5 or FF_i )
	begin
	rl_a34_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a34_t4 = ( ( { 9{ FF_i } } & rl_a34_t5 )
		| ( { 9{ rl_a34_t4_c1 } } & rl_a34_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_218 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h01 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h02 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h03 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h04 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h05 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h06 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h07 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h08 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h09 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h0a :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h0b :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h0c :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h0d :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h0e :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h0f :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h10 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h11 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h12 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h13 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h14 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h15 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h16 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h17 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h18 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h19 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h1a :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h1b :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h1c :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h1d :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h1e :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h1f :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h20 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h21 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h22 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h23 :
		rl_a35_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h24 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h25 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h26 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h27 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h28 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h29 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h2a :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h2b :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h2c :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h2d :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h2e :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h2f :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h30 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h31 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h32 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h33 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h34 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h35 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h36 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h37 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h38 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h39 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h3a :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h3b :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h3c :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h3d :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h3e :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h3f :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h40 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h41 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h42 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h43 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h44 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h45 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h46 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h47 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h48 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h49 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h4a :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h4b :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h4c :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h4d :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h4e :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h4f :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h50 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h51 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h52 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h53 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h54 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h55 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h56 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h57 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h58 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h59 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h5a :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h5b :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h5c :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h5d :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h5e :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h5f :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h60 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h61 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h62 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h63 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h64 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h65 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h66 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h67 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h68 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h69 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h6a :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h6b :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h6c :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h6d :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h6e :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h6f :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h70 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h71 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h72 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h73 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h74 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h75 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h76 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h77 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h78 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h79 :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h7a :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h7b :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h7c :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h7d :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h7e :
		rl_a35_t4_t1 = RG_rl_218 ;
	7'h7f :
		rl_a35_t4_t1 = RG_rl_218 ;
	default :
		rl_a35_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a35_t4_t1 or rl_a35_t5 or FF_i )
	begin
	rl_a35_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a35_t4 = ( ( { 9{ FF_i } } & rl_a35_t5 )
		| ( { 9{ rl_a35_t4_c1 } } & rl_a35_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_219 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h01 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h02 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h03 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h04 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h05 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h06 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h07 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h08 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h09 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h0a :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h0b :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h0c :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h0d :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h0e :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h0f :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h10 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h11 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h12 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h13 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h14 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h15 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h16 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h17 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h18 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h19 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h1a :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h1b :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h1c :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h1d :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h1e :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h1f :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h20 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h21 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h22 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h23 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h24 :
		rl_a36_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h25 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h26 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h27 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h28 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h29 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h2a :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h2b :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h2c :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h2d :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h2e :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h2f :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h30 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h31 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h32 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h33 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h34 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h35 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h36 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h37 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h38 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h39 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h3a :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h3b :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h3c :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h3d :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h3e :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h3f :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h40 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h41 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h42 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h43 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h44 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h45 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h46 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h47 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h48 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h49 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h4a :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h4b :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h4c :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h4d :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h4e :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h4f :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h50 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h51 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h52 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h53 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h54 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h55 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h56 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h57 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h58 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h59 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h5a :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h5b :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h5c :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h5d :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h5e :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h5f :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h60 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h61 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h62 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h63 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h64 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h65 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h66 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h67 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h68 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h69 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h6a :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h6b :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h6c :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h6d :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h6e :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h6f :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h70 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h71 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h72 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h73 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h74 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h75 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h76 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h77 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h78 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h79 :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h7a :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h7b :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h7c :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h7d :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h7e :
		rl_a36_t4_t1 = RG_rl_219 ;
	7'h7f :
		rl_a36_t4_t1 = RG_rl_219 ;
	default :
		rl_a36_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a36_t4_t1 or rl_a36_t5 or FF_i )
	begin
	rl_a36_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a36_t4 = ( ( { 9{ FF_i } } & rl_a36_t5 )
		| ( { 9{ rl_a36_t4_c1 } } & rl_a36_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_220 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h01 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h02 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h03 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h04 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h05 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h06 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h07 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h08 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h09 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h0a :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h0b :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h0c :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h0d :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h0e :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h0f :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h10 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h11 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h12 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h13 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h14 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h15 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h16 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h17 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h18 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h19 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h1a :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h1b :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h1c :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h1d :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h1e :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h1f :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h20 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h21 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h22 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h23 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h24 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h25 :
		rl_a37_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h26 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h27 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h28 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h29 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h2a :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h2b :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h2c :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h2d :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h2e :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h2f :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h30 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h31 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h32 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h33 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h34 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h35 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h36 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h37 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h38 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h39 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h3a :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h3b :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h3c :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h3d :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h3e :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h3f :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h40 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h41 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h42 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h43 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h44 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h45 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h46 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h47 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h48 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h49 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h4a :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h4b :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h4c :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h4d :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h4e :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h4f :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h50 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h51 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h52 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h53 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h54 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h55 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h56 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h57 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h58 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h59 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h5a :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h5b :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h5c :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h5d :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h5e :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h5f :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h60 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h61 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h62 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h63 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h64 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h65 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h66 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h67 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h68 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h69 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h6a :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h6b :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h6c :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h6d :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h6e :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h6f :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h70 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h71 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h72 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h73 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h74 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h75 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h76 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h77 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h78 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h79 :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h7a :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h7b :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h7c :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h7d :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h7e :
		rl_a37_t4_t1 = RG_rl_220 ;
	7'h7f :
		rl_a37_t4_t1 = RG_rl_220 ;
	default :
		rl_a37_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a37_t4_t1 or rl_a37_t5 or FF_i )
	begin
	rl_a37_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a37_t4 = ( ( { 9{ FF_i } } & rl_a37_t5 )
		| ( { 9{ rl_a37_t4_c1 } } & rl_a37_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_221 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h01 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h02 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h03 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h04 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h05 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h06 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h07 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h08 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h09 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h0a :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h0b :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h0c :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h0d :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h0e :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h0f :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h10 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h11 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h12 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h13 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h14 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h15 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h16 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h17 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h18 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h19 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h1a :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h1b :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h1c :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h1d :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h1e :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h1f :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h20 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h21 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h22 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h23 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h24 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h25 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h26 :
		rl_a38_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h27 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h28 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h29 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h2a :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h2b :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h2c :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h2d :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h2e :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h2f :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h30 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h31 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h32 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h33 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h34 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h35 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h36 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h37 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h38 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h39 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h3a :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h3b :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h3c :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h3d :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h3e :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h3f :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h40 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h41 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h42 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h43 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h44 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h45 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h46 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h47 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h48 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h49 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h4a :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h4b :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h4c :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h4d :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h4e :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h4f :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h50 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h51 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h52 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h53 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h54 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h55 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h56 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h57 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h58 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h59 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h5a :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h5b :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h5c :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h5d :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h5e :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h5f :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h60 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h61 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h62 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h63 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h64 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h65 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h66 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h67 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h68 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h69 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h6a :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h6b :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h6c :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h6d :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h6e :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h6f :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h70 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h71 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h72 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h73 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h74 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h75 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h76 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h77 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h78 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h79 :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h7a :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h7b :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h7c :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h7d :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h7e :
		rl_a38_t4_t1 = RG_rl_221 ;
	7'h7f :
		rl_a38_t4_t1 = RG_rl_221 ;
	default :
		rl_a38_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a38_t4_t1 or rl_a38_t5 or FF_i )
	begin
	rl_a38_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a38_t4 = ( ( { 9{ FF_i } } & rl_a38_t5 )
		| ( { 9{ rl_a38_t4_c1 } } & rl_a38_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_222 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h01 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h02 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h03 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h04 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h05 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h06 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h07 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h08 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h09 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h0a :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h0b :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h0c :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h0d :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h0e :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h0f :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h10 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h11 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h12 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h13 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h14 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h15 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h16 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h17 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h18 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h19 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h1a :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h1b :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h1c :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h1d :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h1e :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h1f :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h20 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h21 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h22 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h23 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h24 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h25 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h26 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h27 :
		rl_a39_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h28 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h29 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h2a :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h2b :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h2c :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h2d :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h2e :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h2f :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h30 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h31 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h32 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h33 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h34 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h35 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h36 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h37 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h38 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h39 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h3a :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h3b :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h3c :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h3d :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h3e :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h3f :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h40 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h41 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h42 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h43 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h44 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h45 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h46 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h47 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h48 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h49 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h4a :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h4b :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h4c :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h4d :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h4e :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h4f :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h50 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h51 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h52 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h53 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h54 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h55 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h56 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h57 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h58 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h59 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h5a :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h5b :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h5c :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h5d :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h5e :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h5f :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h60 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h61 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h62 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h63 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h64 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h65 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h66 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h67 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h68 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h69 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h6a :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h6b :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h6c :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h6d :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h6e :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h6f :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h70 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h71 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h72 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h73 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h74 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h75 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h76 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h77 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h78 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h79 :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h7a :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h7b :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h7c :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h7d :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h7e :
		rl_a39_t4_t1 = RG_rl_222 ;
	7'h7f :
		rl_a39_t4_t1 = RG_rl_222 ;
	default :
		rl_a39_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a39_t4_t1 or rl_a39_t5 or FF_i )
	begin
	rl_a39_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a39_t4 = ( ( { 9{ FF_i } } & rl_a39_t5 )
		| ( { 9{ rl_a39_t4_c1 } } & rl_a39_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_223 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h01 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h02 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h03 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h04 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h05 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h06 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h07 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h08 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h09 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h0a :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h0b :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h0c :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h0d :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h0e :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h0f :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h10 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h11 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h12 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h13 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h14 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h15 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h16 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h17 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h18 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h19 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h1a :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h1b :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h1c :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h1d :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h1e :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h1f :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h20 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h21 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h22 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h23 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h24 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h25 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h26 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h27 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h28 :
		rl_a40_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h29 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h2a :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h2b :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h2c :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h2d :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h2e :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h2f :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h30 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h31 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h32 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h33 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h34 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h35 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h36 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h37 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h38 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h39 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h3a :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h3b :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h3c :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h3d :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h3e :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h3f :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h40 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h41 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h42 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h43 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h44 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h45 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h46 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h47 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h48 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h49 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h4a :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h4b :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h4c :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h4d :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h4e :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h4f :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h50 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h51 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h52 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h53 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h54 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h55 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h56 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h57 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h58 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h59 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h5a :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h5b :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h5c :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h5d :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h5e :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h5f :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h60 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h61 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h62 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h63 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h64 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h65 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h66 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h67 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h68 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h69 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h6a :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h6b :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h6c :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h6d :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h6e :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h6f :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h70 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h71 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h72 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h73 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h74 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h75 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h76 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h77 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h78 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h79 :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h7a :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h7b :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h7c :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h7d :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h7e :
		rl_a40_t4_t1 = RG_rl_223 ;
	7'h7f :
		rl_a40_t4_t1 = RG_rl_223 ;
	default :
		rl_a40_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a40_t4_t1 or rl_a40_t5 or FF_i )
	begin
	rl_a40_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a40_t4 = ( ( { 9{ FF_i } } & rl_a40_t5 )
		| ( { 9{ rl_a40_t4_c1 } } & rl_a40_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_224 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h01 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h02 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h03 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h04 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h05 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h06 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h07 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h08 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h09 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h0a :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h0b :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h0c :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h0d :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h0e :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h0f :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h10 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h11 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h12 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h13 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h14 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h15 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h16 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h17 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h18 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h19 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h1a :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h1b :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h1c :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h1d :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h1e :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h1f :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h20 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h21 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h22 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h23 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h24 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h25 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h26 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h27 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h28 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h29 :
		rl_a41_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h2a :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h2b :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h2c :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h2d :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h2e :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h2f :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h30 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h31 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h32 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h33 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h34 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h35 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h36 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h37 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h38 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h39 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h3a :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h3b :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h3c :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h3d :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h3e :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h3f :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h40 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h41 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h42 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h43 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h44 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h45 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h46 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h47 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h48 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h49 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h4a :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h4b :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h4c :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h4d :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h4e :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h4f :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h50 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h51 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h52 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h53 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h54 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h55 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h56 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h57 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h58 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h59 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h5a :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h5b :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h5c :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h5d :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h5e :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h5f :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h60 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h61 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h62 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h63 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h64 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h65 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h66 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h67 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h68 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h69 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h6a :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h6b :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h6c :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h6d :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h6e :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h6f :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h70 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h71 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h72 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h73 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h74 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h75 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h76 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h77 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h78 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h79 :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h7a :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h7b :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h7c :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h7d :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h7e :
		rl_a41_t4_t1 = RG_rl_224 ;
	7'h7f :
		rl_a41_t4_t1 = RG_rl_224 ;
	default :
		rl_a41_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a41_t4_t1 or rl_a41_t5 or FF_i )
	begin
	rl_a41_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a41_t4 = ( ( { 9{ FF_i } } & rl_a41_t5 )
		| ( { 9{ rl_a41_t4_c1 } } & rl_a41_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_225 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h01 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h02 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h03 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h04 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h05 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h06 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h07 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h08 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h09 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h0a :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h0b :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h0c :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h0d :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h0e :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h0f :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h10 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h11 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h12 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h13 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h14 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h15 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h16 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h17 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h18 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h19 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h1a :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h1b :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h1c :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h1d :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h1e :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h1f :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h20 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h21 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h22 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h23 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h24 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h25 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h26 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h27 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h28 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h29 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h2a :
		rl_a42_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h2b :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h2c :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h2d :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h2e :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h2f :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h30 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h31 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h32 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h33 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h34 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h35 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h36 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h37 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h38 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h39 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h3a :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h3b :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h3c :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h3d :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h3e :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h3f :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h40 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h41 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h42 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h43 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h44 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h45 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h46 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h47 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h48 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h49 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h4a :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h4b :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h4c :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h4d :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h4e :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h4f :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h50 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h51 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h52 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h53 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h54 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h55 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h56 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h57 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h58 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h59 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h5a :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h5b :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h5c :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h5d :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h5e :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h5f :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h60 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h61 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h62 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h63 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h64 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h65 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h66 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h67 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h68 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h69 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h6a :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h6b :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h6c :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h6d :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h6e :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h6f :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h70 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h71 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h72 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h73 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h74 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h75 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h76 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h77 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h78 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h79 :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h7a :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h7b :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h7c :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h7d :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h7e :
		rl_a42_t4_t1 = RG_rl_225 ;
	7'h7f :
		rl_a42_t4_t1 = RG_rl_225 ;
	default :
		rl_a42_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a42_t4_t1 or rl_a42_t5 or FF_i )
	begin
	rl_a42_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a42_t4 = ( ( { 9{ FF_i } } & rl_a42_t5 )
		| ( { 9{ rl_a42_t4_c1 } } & rl_a42_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_226 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h01 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h02 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h03 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h04 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h05 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h06 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h07 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h08 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h09 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h0a :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h0b :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h0c :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h0d :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h0e :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h0f :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h10 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h11 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h12 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h13 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h14 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h15 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h16 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h17 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h18 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h19 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h1a :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h1b :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h1c :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h1d :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h1e :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h1f :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h20 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h21 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h22 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h23 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h24 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h25 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h26 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h27 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h28 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h29 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h2a :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h2b :
		rl_a43_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h2c :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h2d :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h2e :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h2f :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h30 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h31 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h32 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h33 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h34 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h35 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h36 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h37 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h38 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h39 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h3a :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h3b :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h3c :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h3d :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h3e :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h3f :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h40 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h41 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h42 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h43 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h44 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h45 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h46 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h47 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h48 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h49 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h4a :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h4b :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h4c :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h4d :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h4e :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h4f :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h50 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h51 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h52 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h53 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h54 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h55 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h56 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h57 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h58 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h59 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h5a :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h5b :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h5c :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h5d :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h5e :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h5f :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h60 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h61 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h62 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h63 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h64 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h65 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h66 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h67 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h68 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h69 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h6a :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h6b :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h6c :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h6d :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h6e :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h6f :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h70 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h71 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h72 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h73 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h74 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h75 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h76 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h77 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h78 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h79 :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h7a :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h7b :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h7c :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h7d :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h7e :
		rl_a43_t4_t1 = RG_rl_226 ;
	7'h7f :
		rl_a43_t4_t1 = RG_rl_226 ;
	default :
		rl_a43_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a43_t4_t1 or rl_a43_t5 or FF_i )
	begin
	rl_a43_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a43_t4 = ( ( { 9{ FF_i } } & rl_a43_t5 )
		| ( { 9{ rl_a43_t4_c1 } } & rl_a43_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_227 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h01 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h02 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h03 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h04 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h05 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h06 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h07 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h08 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h09 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h0a :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h0b :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h0c :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h0d :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h0e :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h0f :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h10 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h11 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h12 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h13 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h14 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h15 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h16 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h17 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h18 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h19 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h1a :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h1b :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h1c :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h1d :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h1e :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h1f :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h20 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h21 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h22 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h23 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h24 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h25 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h26 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h27 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h28 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h29 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h2a :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h2b :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h2c :
		rl_a44_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h2d :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h2e :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h2f :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h30 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h31 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h32 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h33 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h34 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h35 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h36 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h37 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h38 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h39 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h3a :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h3b :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h3c :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h3d :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h3e :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h3f :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h40 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h41 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h42 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h43 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h44 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h45 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h46 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h47 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h48 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h49 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h4a :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h4b :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h4c :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h4d :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h4e :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h4f :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h50 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h51 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h52 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h53 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h54 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h55 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h56 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h57 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h58 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h59 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h5a :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h5b :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h5c :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h5d :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h5e :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h5f :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h60 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h61 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h62 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h63 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h64 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h65 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h66 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h67 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h68 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h69 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h6a :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h6b :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h6c :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h6d :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h6e :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h6f :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h70 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h71 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h72 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h73 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h74 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h75 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h76 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h77 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h78 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h79 :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h7a :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h7b :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h7c :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h7d :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h7e :
		rl_a44_t4_t1 = RG_rl_227 ;
	7'h7f :
		rl_a44_t4_t1 = RG_rl_227 ;
	default :
		rl_a44_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a44_t4_t1 or rl_a44_t5 or FF_i )
	begin
	rl_a44_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a44_t4 = ( ( { 9{ FF_i } } & rl_a44_t5 )
		| ( { 9{ rl_a44_t4_c1 } } & rl_a44_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_228 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h01 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h02 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h03 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h04 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h05 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h06 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h07 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h08 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h09 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h0a :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h0b :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h0c :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h0d :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h0e :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h0f :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h10 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h11 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h12 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h13 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h14 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h15 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h16 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h17 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h18 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h19 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h1a :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h1b :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h1c :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h1d :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h1e :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h1f :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h20 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h21 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h22 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h23 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h24 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h25 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h26 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h27 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h28 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h29 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h2a :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h2b :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h2c :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h2d :
		rl_a45_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h2e :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h2f :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h30 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h31 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h32 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h33 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h34 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h35 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h36 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h37 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h38 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h39 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h3a :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h3b :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h3c :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h3d :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h3e :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h3f :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h40 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h41 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h42 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h43 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h44 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h45 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h46 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h47 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h48 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h49 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h4a :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h4b :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h4c :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h4d :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h4e :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h4f :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h50 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h51 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h52 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h53 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h54 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h55 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h56 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h57 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h58 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h59 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h5a :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h5b :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h5c :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h5d :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h5e :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h5f :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h60 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h61 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h62 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h63 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h64 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h65 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h66 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h67 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h68 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h69 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h6a :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h6b :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h6c :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h6d :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h6e :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h6f :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h70 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h71 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h72 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h73 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h74 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h75 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h76 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h77 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h78 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h79 :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h7a :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h7b :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h7c :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h7d :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h7e :
		rl_a45_t4_t1 = RG_rl_228 ;
	7'h7f :
		rl_a45_t4_t1 = RG_rl_228 ;
	default :
		rl_a45_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a45_t4_t1 or rl_a45_t5 or FF_i )
	begin
	rl_a45_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a45_t4 = ( ( { 9{ FF_i } } & rl_a45_t5 )
		| ( { 9{ rl_a45_t4_c1 } } & rl_a45_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_229 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h01 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h02 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h03 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h04 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h05 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h06 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h07 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h08 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h09 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h0a :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h0b :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h0c :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h0d :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h0e :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h0f :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h10 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h11 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h12 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h13 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h14 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h15 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h16 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h17 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h18 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h19 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h1a :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h1b :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h1c :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h1d :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h1e :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h1f :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h20 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h21 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h22 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h23 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h24 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h25 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h26 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h27 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h28 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h29 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h2a :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h2b :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h2c :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h2d :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h2e :
		rl_a46_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h2f :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h30 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h31 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h32 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h33 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h34 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h35 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h36 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h37 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h38 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h39 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h3a :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h3b :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h3c :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h3d :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h3e :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h3f :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h40 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h41 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h42 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h43 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h44 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h45 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h46 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h47 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h48 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h49 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h4a :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h4b :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h4c :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h4d :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h4e :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h4f :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h50 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h51 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h52 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h53 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h54 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h55 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h56 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h57 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h58 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h59 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h5a :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h5b :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h5c :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h5d :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h5e :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h5f :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h60 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h61 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h62 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h63 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h64 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h65 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h66 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h67 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h68 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h69 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h6a :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h6b :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h6c :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h6d :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h6e :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h6f :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h70 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h71 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h72 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h73 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h74 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h75 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h76 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h77 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h78 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h79 :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h7a :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h7b :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h7c :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h7d :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h7e :
		rl_a46_t4_t1 = RG_rl_229 ;
	7'h7f :
		rl_a46_t4_t1 = RG_rl_229 ;
	default :
		rl_a46_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a46_t4_t1 or rl_a46_t5 or FF_i )
	begin
	rl_a46_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a46_t4 = ( ( { 9{ FF_i } } & rl_a46_t5 )
		| ( { 9{ rl_a46_t4_c1 } } & rl_a46_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_230 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h01 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h02 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h03 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h04 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h05 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h06 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h07 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h08 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h09 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h0a :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h0b :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h0c :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h0d :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h0e :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h0f :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h10 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h11 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h12 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h13 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h14 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h15 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h16 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h17 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h18 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h19 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h1a :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h1b :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h1c :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h1d :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h1e :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h1f :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h20 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h21 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h22 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h23 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h24 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h25 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h26 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h27 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h28 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h29 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h2a :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h2b :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h2c :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h2d :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h2e :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h2f :
		rl_a47_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h30 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h31 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h32 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h33 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h34 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h35 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h36 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h37 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h38 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h39 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h3a :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h3b :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h3c :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h3d :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h3e :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h3f :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h40 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h41 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h42 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h43 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h44 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h45 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h46 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h47 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h48 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h49 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h4a :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h4b :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h4c :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h4d :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h4e :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h4f :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h50 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h51 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h52 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h53 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h54 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h55 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h56 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h57 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h58 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h59 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h5a :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h5b :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h5c :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h5d :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h5e :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h5f :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h60 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h61 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h62 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h63 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h64 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h65 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h66 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h67 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h68 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h69 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h6a :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h6b :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h6c :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h6d :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h6e :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h6f :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h70 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h71 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h72 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h73 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h74 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h75 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h76 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h77 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h78 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h79 :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h7a :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h7b :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h7c :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h7d :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h7e :
		rl_a47_t4_t1 = RG_rl_230 ;
	7'h7f :
		rl_a47_t4_t1 = RG_rl_230 ;
	default :
		rl_a47_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a47_t4_t1 or rl_a47_t5 or FF_i )
	begin
	rl_a47_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a47_t4 = ( ( { 9{ FF_i } } & rl_a47_t5 )
		| ( { 9{ rl_a47_t4_c1 } } & rl_a47_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_231 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h01 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h02 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h03 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h04 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h05 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h06 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h07 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h08 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h09 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h0a :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h0b :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h0c :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h0d :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h0e :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h0f :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h10 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h11 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h12 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h13 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h14 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h15 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h16 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h17 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h18 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h19 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h1a :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h1b :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h1c :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h1d :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h1e :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h1f :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h20 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h21 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h22 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h23 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h24 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h25 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h26 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h27 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h28 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h29 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h2a :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h2b :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h2c :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h2d :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h2e :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h2f :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h30 :
		rl_a48_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h31 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h32 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h33 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h34 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h35 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h36 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h37 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h38 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h39 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h3a :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h3b :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h3c :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h3d :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h3e :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h3f :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h40 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h41 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h42 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h43 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h44 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h45 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h46 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h47 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h48 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h49 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h4a :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h4b :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h4c :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h4d :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h4e :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h4f :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h50 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h51 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h52 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h53 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h54 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h55 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h56 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h57 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h58 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h59 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h5a :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h5b :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h5c :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h5d :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h5e :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h5f :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h60 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h61 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h62 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h63 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h64 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h65 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h66 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h67 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h68 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h69 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h6a :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h6b :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h6c :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h6d :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h6e :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h6f :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h70 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h71 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h72 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h73 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h74 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h75 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h76 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h77 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h78 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h79 :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h7a :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h7b :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h7c :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h7d :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h7e :
		rl_a48_t4_t1 = RG_rl_231 ;
	7'h7f :
		rl_a48_t4_t1 = RG_rl_231 ;
	default :
		rl_a48_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a48_t4_t1 or rl_a48_t5 or FF_i )
	begin
	rl_a48_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a48_t4 = ( ( { 9{ FF_i } } & rl_a48_t5 )
		| ( { 9{ rl_a48_t4_c1 } } & rl_a48_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_232 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h01 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h02 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h03 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h04 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h05 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h06 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h07 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h08 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h09 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h0a :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h0b :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h0c :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h0d :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h0e :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h0f :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h10 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h11 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h12 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h13 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h14 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h15 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h16 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h17 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h18 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h19 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h1a :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h1b :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h1c :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h1d :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h1e :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h1f :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h20 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h21 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h22 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h23 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h24 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h25 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h26 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h27 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h28 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h29 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h2a :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h2b :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h2c :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h2d :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h2e :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h2f :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h30 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h31 :
		rl_a49_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h32 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h33 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h34 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h35 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h36 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h37 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h38 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h39 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h3a :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h3b :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h3c :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h3d :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h3e :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h3f :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h40 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h41 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h42 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h43 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h44 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h45 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h46 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h47 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h48 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h49 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h4a :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h4b :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h4c :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h4d :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h4e :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h4f :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h50 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h51 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h52 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h53 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h54 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h55 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h56 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h57 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h58 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h59 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h5a :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h5b :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h5c :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h5d :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h5e :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h5f :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h60 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h61 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h62 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h63 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h64 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h65 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h66 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h67 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h68 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h69 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h6a :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h6b :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h6c :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h6d :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h6e :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h6f :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h70 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h71 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h72 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h73 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h74 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h75 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h76 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h77 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h78 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h79 :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h7a :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h7b :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h7c :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h7d :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h7e :
		rl_a49_t4_t1 = RG_rl_232 ;
	7'h7f :
		rl_a49_t4_t1 = RG_rl_232 ;
	default :
		rl_a49_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a49_t4_t1 or rl_a49_t5 or FF_i )
	begin
	rl_a49_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a49_t4 = ( ( { 9{ FF_i } } & rl_a49_t5 )
		| ( { 9{ rl_a49_t4_c1 } } & rl_a49_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_233 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h01 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h02 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h03 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h04 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h05 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h06 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h07 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h08 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h09 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h0a :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h0b :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h0c :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h0d :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h0e :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h0f :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h10 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h11 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h12 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h13 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h14 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h15 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h16 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h17 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h18 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h19 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h1a :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h1b :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h1c :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h1d :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h1e :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h1f :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h20 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h21 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h22 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h23 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h24 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h25 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h26 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h27 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h28 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h29 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h2a :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h2b :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h2c :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h2d :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h2e :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h2f :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h30 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h31 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h32 :
		rl_a50_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h33 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h34 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h35 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h36 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h37 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h38 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h39 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h3a :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h3b :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h3c :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h3d :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h3e :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h3f :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h40 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h41 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h42 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h43 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h44 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h45 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h46 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h47 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h48 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h49 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h4a :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h4b :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h4c :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h4d :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h4e :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h4f :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h50 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h51 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h52 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h53 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h54 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h55 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h56 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h57 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h58 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h59 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h5a :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h5b :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h5c :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h5d :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h5e :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h5f :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h60 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h61 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h62 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h63 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h64 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h65 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h66 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h67 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h68 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h69 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h6a :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h6b :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h6c :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h6d :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h6e :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h6f :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h70 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h71 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h72 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h73 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h74 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h75 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h76 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h77 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h78 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h79 :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h7a :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h7b :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h7c :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h7d :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h7e :
		rl_a50_t4_t1 = RG_rl_233 ;
	7'h7f :
		rl_a50_t4_t1 = RG_rl_233 ;
	default :
		rl_a50_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a50_t4_t1 or rl_a50_t5 or FF_i )
	begin
	rl_a50_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a50_t4 = ( ( { 9{ FF_i } } & rl_a50_t5 )
		| ( { 9{ rl_a50_t4_c1 } } & rl_a50_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_234 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h01 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h02 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h03 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h04 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h05 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h06 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h07 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h08 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h09 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h0a :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h0b :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h0c :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h0d :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h0e :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h0f :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h10 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h11 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h12 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h13 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h14 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h15 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h16 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h17 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h18 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h19 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h1a :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h1b :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h1c :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h1d :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h1e :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h1f :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h20 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h21 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h22 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h23 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h24 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h25 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h26 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h27 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h28 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h29 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h2a :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h2b :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h2c :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h2d :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h2e :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h2f :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h30 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h31 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h32 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h33 :
		rl_a51_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h34 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h35 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h36 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h37 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h38 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h39 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h3a :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h3b :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h3c :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h3d :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h3e :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h3f :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h40 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h41 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h42 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h43 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h44 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h45 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h46 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h47 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h48 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h49 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h4a :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h4b :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h4c :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h4d :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h4e :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h4f :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h50 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h51 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h52 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h53 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h54 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h55 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h56 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h57 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h58 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h59 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h5a :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h5b :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h5c :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h5d :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h5e :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h5f :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h60 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h61 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h62 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h63 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h64 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h65 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h66 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h67 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h68 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h69 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h6a :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h6b :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h6c :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h6d :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h6e :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h6f :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h70 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h71 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h72 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h73 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h74 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h75 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h76 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h77 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h78 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h79 :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h7a :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h7b :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h7c :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h7d :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h7e :
		rl_a51_t4_t1 = RG_rl_234 ;
	7'h7f :
		rl_a51_t4_t1 = RG_rl_234 ;
	default :
		rl_a51_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a51_t4_t1 or rl_a51_t5 or FF_i )
	begin
	rl_a51_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a51_t4 = ( ( { 9{ FF_i } } & rl_a51_t5 )
		| ( { 9{ rl_a51_t4_c1 } } & rl_a51_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_235 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h01 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h02 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h03 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h04 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h05 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h06 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h07 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h08 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h09 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h0a :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h0b :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h0c :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h0d :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h0e :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h0f :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h10 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h11 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h12 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h13 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h14 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h15 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h16 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h17 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h18 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h19 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h1a :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h1b :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h1c :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h1d :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h1e :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h1f :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h20 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h21 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h22 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h23 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h24 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h25 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h26 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h27 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h28 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h29 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h2a :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h2b :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h2c :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h2d :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h2e :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h2f :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h30 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h31 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h32 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h33 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h34 :
		rl_a52_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h35 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h36 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h37 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h38 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h39 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h3a :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h3b :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h3c :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h3d :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h3e :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h3f :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h40 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h41 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h42 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h43 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h44 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h45 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h46 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h47 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h48 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h49 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h4a :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h4b :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h4c :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h4d :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h4e :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h4f :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h50 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h51 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h52 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h53 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h54 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h55 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h56 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h57 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h58 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h59 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h5a :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h5b :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h5c :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h5d :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h5e :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h5f :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h60 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h61 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h62 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h63 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h64 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h65 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h66 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h67 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h68 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h69 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h6a :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h6b :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h6c :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h6d :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h6e :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h6f :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h70 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h71 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h72 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h73 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h74 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h75 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h76 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h77 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h78 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h79 :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h7a :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h7b :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h7c :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h7d :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h7e :
		rl_a52_t4_t1 = RG_rl_235 ;
	7'h7f :
		rl_a52_t4_t1 = RG_rl_235 ;
	default :
		rl_a52_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a52_t4_t1 or rl_a52_t5 or FF_i )
	begin
	rl_a52_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a52_t4 = ( ( { 9{ FF_i } } & rl_a52_t5 )
		| ( { 9{ rl_a52_t4_c1 } } & rl_a52_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_236 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h01 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h02 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h03 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h04 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h05 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h06 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h07 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h08 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h09 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h0a :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h0b :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h0c :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h0d :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h0e :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h0f :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h10 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h11 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h12 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h13 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h14 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h15 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h16 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h17 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h18 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h19 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h1a :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h1b :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h1c :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h1d :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h1e :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h1f :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h20 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h21 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h22 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h23 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h24 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h25 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h26 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h27 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h28 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h29 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h2a :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h2b :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h2c :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h2d :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h2e :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h2f :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h30 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h31 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h32 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h33 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h34 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h35 :
		rl_a53_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h36 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h37 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h38 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h39 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h3a :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h3b :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h3c :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h3d :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h3e :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h3f :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h40 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h41 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h42 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h43 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h44 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h45 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h46 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h47 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h48 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h49 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h4a :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h4b :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h4c :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h4d :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h4e :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h4f :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h50 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h51 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h52 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h53 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h54 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h55 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h56 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h57 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h58 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h59 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h5a :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h5b :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h5c :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h5d :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h5e :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h5f :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h60 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h61 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h62 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h63 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h64 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h65 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h66 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h67 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h68 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h69 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h6a :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h6b :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h6c :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h6d :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h6e :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h6f :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h70 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h71 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h72 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h73 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h74 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h75 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h76 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h77 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h78 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h79 :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h7a :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h7b :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h7c :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h7d :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h7e :
		rl_a53_t4_t1 = RG_rl_236 ;
	7'h7f :
		rl_a53_t4_t1 = RG_rl_236 ;
	default :
		rl_a53_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a53_t4_t1 or rl_a53_t5 or FF_i )
	begin
	rl_a53_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a53_t4 = ( ( { 9{ FF_i } } & rl_a53_t5 )
		| ( { 9{ rl_a53_t4_c1 } } & rl_a53_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_237 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h01 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h02 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h03 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h04 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h05 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h06 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h07 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h08 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h09 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h0a :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h0b :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h0c :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h0d :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h0e :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h0f :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h10 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h11 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h12 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h13 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h14 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h15 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h16 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h17 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h18 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h19 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h1a :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h1b :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h1c :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h1d :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h1e :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h1f :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h20 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h21 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h22 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h23 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h24 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h25 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h26 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h27 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h28 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h29 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h2a :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h2b :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h2c :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h2d :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h2e :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h2f :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h30 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h31 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h32 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h33 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h34 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h35 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h36 :
		rl_a54_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h37 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h38 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h39 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h3a :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h3b :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h3c :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h3d :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h3e :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h3f :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h40 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h41 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h42 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h43 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h44 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h45 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h46 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h47 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h48 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h49 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h4a :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h4b :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h4c :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h4d :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h4e :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h4f :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h50 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h51 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h52 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h53 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h54 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h55 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h56 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h57 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h58 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h59 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h5a :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h5b :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h5c :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h5d :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h5e :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h5f :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h60 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h61 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h62 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h63 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h64 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h65 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h66 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h67 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h68 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h69 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h6a :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h6b :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h6c :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h6d :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h6e :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h6f :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h70 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h71 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h72 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h73 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h74 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h75 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h76 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h77 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h78 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h79 :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h7a :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h7b :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h7c :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h7d :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h7e :
		rl_a54_t4_t1 = RG_rl_237 ;
	7'h7f :
		rl_a54_t4_t1 = RG_rl_237 ;
	default :
		rl_a54_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a54_t4_t1 or rl_a54_t5 or FF_i )
	begin
	rl_a54_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a54_t4 = ( ( { 9{ FF_i } } & rl_a54_t5 )
		| ( { 9{ rl_a54_t4_c1 } } & rl_a54_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_238 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h01 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h02 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h03 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h04 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h05 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h06 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h07 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h08 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h09 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h0a :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h0b :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h0c :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h0d :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h0e :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h0f :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h10 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h11 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h12 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h13 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h14 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h15 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h16 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h17 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h18 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h19 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h1a :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h1b :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h1c :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h1d :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h1e :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h1f :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h20 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h21 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h22 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h23 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h24 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h25 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h26 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h27 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h28 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h29 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h2a :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h2b :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h2c :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h2d :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h2e :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h2f :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h30 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h31 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h32 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h33 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h34 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h35 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h36 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h37 :
		rl_a55_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h38 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h39 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h3a :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h3b :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h3c :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h3d :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h3e :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h3f :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h40 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h41 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h42 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h43 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h44 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h45 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h46 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h47 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h48 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h49 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h4a :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h4b :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h4c :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h4d :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h4e :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h4f :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h50 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h51 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h52 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h53 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h54 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h55 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h56 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h57 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h58 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h59 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h5a :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h5b :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h5c :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h5d :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h5e :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h5f :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h60 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h61 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h62 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h63 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h64 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h65 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h66 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h67 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h68 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h69 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h6a :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h6b :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h6c :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h6d :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h6e :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h6f :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h70 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h71 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h72 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h73 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h74 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h75 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h76 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h77 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h78 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h79 :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h7a :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h7b :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h7c :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h7d :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h7e :
		rl_a55_t4_t1 = RG_rl_238 ;
	7'h7f :
		rl_a55_t4_t1 = RG_rl_238 ;
	default :
		rl_a55_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a55_t4_t1 or rl_a55_t5 or FF_i )
	begin
	rl_a55_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a55_t4 = ( ( { 9{ FF_i } } & rl_a55_t5 )
		| ( { 9{ rl_a55_t4_c1 } } & rl_a55_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_239 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h01 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h02 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h03 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h04 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h05 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h06 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h07 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h08 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h09 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h0a :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h0b :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h0c :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h0d :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h0e :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h0f :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h10 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h11 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h12 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h13 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h14 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h15 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h16 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h17 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h18 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h19 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h1a :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h1b :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h1c :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h1d :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h1e :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h1f :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h20 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h21 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h22 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h23 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h24 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h25 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h26 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h27 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h28 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h29 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h2a :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h2b :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h2c :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h2d :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h2e :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h2f :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h30 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h31 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h32 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h33 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h34 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h35 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h36 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h37 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h38 :
		rl_a56_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h39 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h3a :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h3b :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h3c :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h3d :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h3e :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h3f :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h40 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h41 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h42 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h43 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h44 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h45 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h46 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h47 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h48 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h49 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h4a :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h4b :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h4c :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h4d :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h4e :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h4f :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h50 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h51 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h52 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h53 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h54 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h55 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h56 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h57 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h58 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h59 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h5a :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h5b :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h5c :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h5d :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h5e :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h5f :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h60 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h61 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h62 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h63 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h64 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h65 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h66 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h67 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h68 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h69 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h6a :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h6b :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h6c :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h6d :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h6e :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h6f :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h70 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h71 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h72 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h73 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h74 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h75 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h76 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h77 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h78 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h79 :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h7a :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h7b :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h7c :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h7d :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h7e :
		rl_a56_t4_t1 = RG_rl_239 ;
	7'h7f :
		rl_a56_t4_t1 = RG_rl_239 ;
	default :
		rl_a56_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a56_t4_t1 or rl_a56_t5 or FF_i )
	begin
	rl_a56_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a56_t4 = ( ( { 9{ FF_i } } & rl_a56_t5 )
		| ( { 9{ rl_a56_t4_c1 } } & rl_a56_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_240 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h01 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h02 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h03 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h04 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h05 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h06 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h07 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h08 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h09 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h0a :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h0b :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h0c :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h0d :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h0e :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h0f :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h10 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h11 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h12 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h13 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h14 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h15 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h16 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h17 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h18 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h19 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h1a :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h1b :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h1c :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h1d :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h1e :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h1f :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h20 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h21 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h22 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h23 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h24 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h25 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h26 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h27 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h28 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h29 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h2a :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h2b :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h2c :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h2d :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h2e :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h2f :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h30 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h31 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h32 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h33 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h34 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h35 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h36 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h37 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h38 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h39 :
		rl_a57_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h3a :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h3b :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h3c :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h3d :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h3e :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h3f :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h40 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h41 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h42 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h43 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h44 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h45 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h46 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h47 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h48 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h49 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h4a :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h4b :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h4c :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h4d :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h4e :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h4f :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h50 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h51 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h52 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h53 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h54 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h55 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h56 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h57 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h58 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h59 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h5a :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h5b :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h5c :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h5d :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h5e :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h5f :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h60 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h61 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h62 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h63 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h64 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h65 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h66 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h67 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h68 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h69 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h6a :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h6b :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h6c :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h6d :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h6e :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h6f :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h70 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h71 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h72 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h73 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h74 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h75 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h76 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h77 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h78 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h79 :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h7a :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h7b :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h7c :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h7d :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h7e :
		rl_a57_t4_t1 = RG_rl_240 ;
	7'h7f :
		rl_a57_t4_t1 = RG_rl_240 ;
	default :
		rl_a57_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a57_t4_t1 or rl_a57_t5 or FF_i )
	begin
	rl_a57_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a57_t4 = ( ( { 9{ FF_i } } & rl_a57_t5 )
		| ( { 9{ rl_a57_t4_c1 } } & rl_a57_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_241 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h01 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h02 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h03 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h04 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h05 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h06 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h07 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h08 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h09 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h0a :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h0b :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h0c :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h0d :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h0e :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h0f :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h10 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h11 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h12 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h13 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h14 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h15 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h16 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h17 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h18 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h19 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h1a :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h1b :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h1c :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h1d :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h1e :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h1f :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h20 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h21 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h22 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h23 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h24 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h25 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h26 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h27 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h28 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h29 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h2a :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h2b :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h2c :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h2d :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h2e :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h2f :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h30 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h31 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h32 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h33 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h34 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h35 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h36 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h37 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h38 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h39 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h3a :
		rl_a58_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h3b :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h3c :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h3d :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h3e :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h3f :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h40 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h41 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h42 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h43 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h44 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h45 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h46 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h47 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h48 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h49 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h4a :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h4b :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h4c :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h4d :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h4e :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h4f :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h50 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h51 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h52 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h53 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h54 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h55 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h56 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h57 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h58 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h59 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h5a :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h5b :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h5c :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h5d :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h5e :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h5f :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h60 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h61 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h62 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h63 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h64 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h65 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h66 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h67 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h68 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h69 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h6a :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h6b :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h6c :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h6d :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h6e :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h6f :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h70 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h71 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h72 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h73 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h74 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h75 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h76 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h77 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h78 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h79 :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h7a :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h7b :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h7c :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h7d :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h7e :
		rl_a58_t4_t1 = RG_rl_241 ;
	7'h7f :
		rl_a58_t4_t1 = RG_rl_241 ;
	default :
		rl_a58_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a58_t4_t1 or rl_a58_t5 or FF_i )
	begin
	rl_a58_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a58_t4 = ( ( { 9{ FF_i } } & rl_a58_t5 )
		| ( { 9{ rl_a58_t4_c1 } } & rl_a58_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h01 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h02 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h03 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h04 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h05 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h06 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h07 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h08 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h09 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h0a :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h0b :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h0c :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h0d :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h0e :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h0f :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h10 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h11 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h12 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h13 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h14 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h15 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h16 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h17 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h18 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h19 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h1a :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h1b :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h1c :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h1d :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h1e :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h1f :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h20 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h21 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h22 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h23 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h24 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h25 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h26 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h27 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h28 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h29 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h2a :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h2b :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h2c :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h2d :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h2e :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h2f :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h30 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h31 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h32 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h33 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h34 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h35 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h36 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h37 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h38 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h39 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h3a :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h3b :
		rl_a59_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h3c :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h3d :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h3e :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h3f :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h40 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h41 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h42 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h43 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h44 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h45 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h46 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h47 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h48 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h49 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h4a :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h4b :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h4c :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h4d :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h4e :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h4f :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h50 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h51 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h52 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h53 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h54 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h55 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h56 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h57 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h58 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h59 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h5a :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h5b :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h5c :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h5d :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h5e :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h5f :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h60 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h61 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h62 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h63 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h64 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h65 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h66 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h67 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h68 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h69 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h6a :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h6b :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h6c :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h6d :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h6e :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h6f :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h70 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h71 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h72 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h73 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h74 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h75 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h76 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h77 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h78 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h79 :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h7a :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h7b :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h7c :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h7d :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h7e :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	7'h7f :
		rl_a59_t4_t1 = RG_quantized_block_rl ;
	default :
		rl_a59_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a59_t4_t1 or rl_a59_t5 or FF_i )
	begin
	rl_a59_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a59_t4 = ( ( { 9{ FF_i } } & rl_a59_t5 )
		| ( { 9{ rl_a59_t4_c1 } } & rl_a59_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_1 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h01 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h02 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h03 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h04 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h05 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h06 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h07 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h08 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h09 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h0a :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h0b :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h0c :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h0d :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h0e :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h0f :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h10 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h11 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h12 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h13 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h14 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h15 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h16 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h17 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h18 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h19 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h1a :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h1b :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h1c :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h1d :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h1e :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h1f :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h20 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h21 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h22 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h23 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h24 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h25 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h26 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h27 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h28 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h29 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h2a :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h2b :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h2c :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h2d :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h2e :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h2f :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h30 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h31 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h32 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h33 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h34 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h35 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h36 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h37 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h38 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h39 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h3a :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h3b :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h3c :
		rl_a60_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h3d :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h3e :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h3f :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h40 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h41 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h42 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h43 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h44 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h45 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h46 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h47 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h48 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h49 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h4a :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h4b :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h4c :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h4d :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h4e :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h4f :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h50 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h51 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h52 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h53 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h54 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h55 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h56 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h57 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h58 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h59 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h5a :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h5b :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h5c :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h5d :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h5e :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h5f :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h60 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h61 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h62 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h63 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h64 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h65 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h66 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h67 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h68 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h69 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h6a :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h6b :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h6c :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h6d :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h6e :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h6f :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h70 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h71 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h72 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h73 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h74 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h75 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h76 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h77 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h78 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h79 :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h7a :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h7b :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h7c :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h7d :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h7e :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	7'h7f :
		rl_a60_t4_t1 = RG_quantized_block_rl_1 ;
	default :
		rl_a60_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a60_t4_t1 or rl_a60_t5 or FF_i )
	begin
	rl_a60_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a60_t4 = ( ( { 9{ FF_i } } & rl_a60_t5 )
		| ( { 9{ rl_a60_t4_c1 } } & rl_a60_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_2 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h01 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h02 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h03 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h04 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h05 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h06 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h07 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h08 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h09 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h0a :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h0b :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h0c :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h0d :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h0e :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h0f :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h10 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h11 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h12 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h13 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h14 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h15 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h16 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h17 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h18 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h19 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h1a :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h1b :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h1c :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h1d :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h1e :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h1f :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h20 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h21 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h22 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h23 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h24 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h25 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h26 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h27 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h28 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h29 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h2a :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h2b :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h2c :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h2d :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h2e :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h2f :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h30 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h31 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h32 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h33 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h34 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h35 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h36 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h37 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h38 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h39 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h3a :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h3b :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h3c :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h3d :
		rl_a61_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h3e :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h3f :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h40 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h41 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h42 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h43 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h44 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h45 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h46 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h47 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h48 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h49 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h4a :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h4b :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h4c :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h4d :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h4e :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h4f :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h50 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h51 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h52 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h53 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h54 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h55 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h56 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h57 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h58 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h59 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h5a :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h5b :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h5c :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h5d :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h5e :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h5f :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h60 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h61 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h62 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h63 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h64 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h65 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h66 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h67 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h68 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h69 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h6a :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h6b :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h6c :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h6d :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h6e :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h6f :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h70 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h71 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h72 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h73 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h74 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h75 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h76 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h77 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h78 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h79 :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h7a :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h7b :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h7c :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h7d :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h7e :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	7'h7f :
		rl_a61_t4_t1 = RG_quantized_block_rl_2 ;
	default :
		rl_a61_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a61_t4_t1 or rl_a61_t5 or FF_i )
	begin
	rl_a61_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a61_t4 = ( ( { 9{ FF_i } } & rl_a61_t5 )
		| ( { 9{ rl_a61_t4_c1 } } & rl_a61_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_3 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h01 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h02 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h03 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h04 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h05 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h06 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h07 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h08 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h09 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h0a :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h0b :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h0c :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h0d :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h0e :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h0f :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h10 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h11 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h12 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h13 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h14 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h15 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h16 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h17 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h18 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h19 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h1a :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h1b :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h1c :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h1d :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h1e :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h1f :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h20 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h21 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h22 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h23 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h24 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h25 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h26 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h27 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h28 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h29 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h2a :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h2b :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h2c :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h2d :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h2e :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h2f :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h30 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h31 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h32 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h33 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h34 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h35 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h36 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h37 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h38 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h39 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h3a :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h3b :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h3c :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h3d :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h3e :
		rl_a62_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h3f :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h40 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h41 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h42 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h43 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h44 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h45 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h46 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h47 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h48 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h49 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h4a :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h4b :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h4c :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h4d :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h4e :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h4f :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h50 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h51 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h52 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h53 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h54 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h55 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h56 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h57 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h58 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h59 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h5a :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h5b :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h5c :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h5d :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h5e :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h5f :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h60 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h61 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h62 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h63 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h64 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h65 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h66 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h67 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h68 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h69 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h6a :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h6b :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h6c :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h6d :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h6e :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h6f :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h70 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h71 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h72 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h73 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h74 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h75 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h76 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h77 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h78 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h79 :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h7a :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h7b :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h7c :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h7d :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h7e :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	7'h7f :
		rl_a62_t4_t1 = RG_quantized_block_rl_3 ;
	default :
		rl_a62_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a62_t4_t1 or rl_a62_t5 or FF_i )
	begin
	rl_a62_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a62_t4 = ( ( { 9{ FF_i } } & rl_a62_t5 )
		| ( { 9{ rl_a62_t4_c1 } } & rl_a62_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_4 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h01 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h02 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h03 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h04 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h05 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h06 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h07 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h08 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h09 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h0a :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h0b :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h0c :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h0d :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h0e :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h0f :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h10 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h11 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h12 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h13 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h14 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h15 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h16 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h17 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h18 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h19 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h1a :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h1b :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h1c :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h1d :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h1e :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h1f :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h20 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h21 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h22 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h23 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h24 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h25 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h26 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h27 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h28 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h29 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h2a :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h2b :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h2c :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h2d :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h2e :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h2f :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h30 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h31 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h32 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h33 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h34 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h35 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h36 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h37 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h38 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h39 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h3a :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h3b :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h3c :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h3d :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h3e :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h3f :
		rl_a63_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h40 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h41 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h42 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h43 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h44 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h45 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h46 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h47 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h48 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h49 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h4a :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h4b :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h4c :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h4d :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h4e :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h4f :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h50 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h51 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h52 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h53 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h54 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h55 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h56 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h57 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h58 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h59 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h5a :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h5b :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h5c :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h5d :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h5e :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h5f :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h60 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h61 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h62 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h63 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h64 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h65 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h66 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h67 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h68 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h69 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h6a :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h6b :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h6c :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h6d :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h6e :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h6f :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h70 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h71 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h72 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h73 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h74 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h75 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h76 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h77 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h78 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h79 :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h7a :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h7b :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h7c :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h7d :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h7e :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	7'h7f :
		rl_a63_t4_t1 = RG_quantized_block_rl_4 ;
	default :
		rl_a63_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a63_t4_t1 or rl_a63_t5 or FF_i )
	begin
	rl_a63_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a63_t4 = ( ( { 9{ FF_i } } & rl_a63_t5 )
		| ( { 9{ rl_a63_t4_c1 } } & rl_a63_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_5 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h01 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h02 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h03 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h04 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h05 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h06 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h07 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h08 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h09 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h0a :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h0b :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h0c :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h0d :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h0e :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h0f :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h10 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h11 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h12 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h13 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h14 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h15 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h16 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h17 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h18 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h19 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h1a :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h1b :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h1c :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h1d :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h1e :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h1f :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h20 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h21 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h22 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h23 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h24 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h25 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h26 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h27 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h28 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h29 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h2a :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h2b :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h2c :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h2d :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h2e :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h2f :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h30 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h31 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h32 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h33 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h34 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h35 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h36 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h37 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h38 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h39 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h3a :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h3b :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h3c :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h3d :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h3e :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h3f :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h40 :
		rl_a64_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h41 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h42 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h43 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h44 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h45 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h46 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h47 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h48 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h49 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h4a :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h4b :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h4c :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h4d :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h4e :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h4f :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h50 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h51 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h52 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h53 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h54 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h55 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h56 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h57 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h58 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h59 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h5a :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h5b :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h5c :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h5d :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h5e :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h5f :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h60 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h61 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h62 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h63 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h64 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h65 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h66 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h67 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h68 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h69 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h6a :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h6b :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h6c :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h6d :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h6e :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h6f :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h70 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h71 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h72 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h73 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h74 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h75 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h76 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h77 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h78 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h79 :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h7a :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h7b :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h7c :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h7d :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h7e :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	7'h7f :
		rl_a64_t4_t1 = RG_quantized_block_rl_5 ;
	default :
		rl_a64_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a64_t4_t1 or rl_a64_t5 or FF_i )
	begin
	rl_a64_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a64_t4 = ( ( { 9{ FF_i } } & rl_a64_t5 )
		| ( { 9{ rl_a64_t4_c1 } } & rl_a64_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_6 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h01 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h02 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h03 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h04 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h05 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h06 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h07 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h08 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h09 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h0a :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h0b :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h0c :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h0d :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h0e :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h0f :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h10 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h11 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h12 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h13 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h14 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h15 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h16 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h17 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h18 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h19 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h1a :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h1b :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h1c :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h1d :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h1e :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h1f :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h20 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h21 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h22 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h23 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h24 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h25 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h26 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h27 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h28 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h29 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h2a :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h2b :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h2c :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h2d :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h2e :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h2f :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h30 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h31 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h32 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h33 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h34 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h35 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h36 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h37 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h38 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h39 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h3a :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h3b :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h3c :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h3d :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h3e :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h3f :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h40 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h41 :
		rl_a65_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h42 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h43 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h44 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h45 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h46 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h47 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h48 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h49 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h4a :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h4b :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h4c :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h4d :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h4e :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h4f :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h50 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h51 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h52 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h53 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h54 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h55 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h56 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h57 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h58 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h59 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h5a :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h5b :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h5c :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h5d :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h5e :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h5f :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h60 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h61 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h62 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h63 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h64 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h65 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h66 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h67 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h68 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h69 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h6a :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h6b :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h6c :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h6d :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h6e :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h6f :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h70 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h71 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h72 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h73 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h74 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h75 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h76 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h77 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h78 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h79 :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h7a :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h7b :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h7c :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h7d :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h7e :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	7'h7f :
		rl_a65_t4_t1 = RG_quantized_block_rl_6 ;
	default :
		rl_a65_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a65_t4_t1 or rl_a65_t5 or FF_i )
	begin
	rl_a65_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a65_t4 = ( ( { 9{ FF_i } } & rl_a65_t5 )
		| ( { 9{ rl_a65_t4_c1 } } & rl_a65_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_7 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h01 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h02 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h03 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h04 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h05 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h06 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h07 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h08 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h09 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h0a :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h0b :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h0c :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h0d :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h0e :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h0f :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h10 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h11 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h12 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h13 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h14 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h15 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h16 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h17 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h18 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h19 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h1a :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h1b :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h1c :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h1d :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h1e :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h1f :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h20 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h21 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h22 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h23 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h24 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h25 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h26 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h27 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h28 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h29 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h2a :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h2b :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h2c :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h2d :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h2e :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h2f :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h30 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h31 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h32 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h33 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h34 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h35 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h36 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h37 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h38 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h39 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h3a :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h3b :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h3c :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h3d :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h3e :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h3f :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h40 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h41 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h42 :
		rl_a66_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h43 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h44 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h45 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h46 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h47 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h48 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h49 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h4a :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h4b :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h4c :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h4d :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h4e :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h4f :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h50 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h51 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h52 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h53 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h54 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h55 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h56 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h57 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h58 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h59 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h5a :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h5b :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h5c :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h5d :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h5e :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h5f :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h60 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h61 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h62 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h63 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h64 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h65 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h66 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h67 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h68 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h69 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h6a :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h6b :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h6c :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h6d :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h6e :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h6f :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h70 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h71 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h72 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h73 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h74 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h75 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h76 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h77 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h78 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h79 :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h7a :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h7b :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h7c :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h7d :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h7e :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	7'h7f :
		rl_a66_t4_t1 = RG_quantized_block_rl_7 ;
	default :
		rl_a66_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a66_t4_t1 or rl_a66_t5 or FF_i )
	begin
	rl_a66_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a66_t4 = ( ( { 9{ FF_i } } & rl_a66_t5 )
		| ( { 9{ rl_a66_t4_c1 } } & rl_a66_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_8 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h01 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h02 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h03 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h04 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h05 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h06 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h07 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h08 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h09 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h0a :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h0b :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h0c :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h0d :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h0e :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h0f :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h10 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h11 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h12 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h13 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h14 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h15 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h16 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h17 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h18 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h19 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h1a :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h1b :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h1c :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h1d :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h1e :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h1f :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h20 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h21 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h22 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h23 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h24 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h25 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h26 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h27 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h28 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h29 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h2a :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h2b :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h2c :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h2d :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h2e :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h2f :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h30 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h31 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h32 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h33 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h34 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h35 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h36 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h37 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h38 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h39 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h3a :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h3b :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h3c :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h3d :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h3e :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h3f :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h40 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h41 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h42 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h43 :
		rl_a67_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h44 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h45 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h46 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h47 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h48 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h49 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h4a :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h4b :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h4c :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h4d :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h4e :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h4f :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h50 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h51 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h52 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h53 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h54 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h55 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h56 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h57 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h58 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h59 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h5a :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h5b :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h5c :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h5d :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h5e :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h5f :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h60 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h61 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h62 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h63 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h64 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h65 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h66 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h67 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h68 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h69 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h6a :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h6b :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h6c :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h6d :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h6e :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h6f :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h70 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h71 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h72 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h73 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h74 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h75 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h76 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h77 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h78 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h79 :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h7a :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h7b :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h7c :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h7d :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h7e :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	7'h7f :
		rl_a67_t4_t1 = RG_quantized_block_rl_8 ;
	default :
		rl_a67_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a67_t4_t1 or rl_a67_t5 or FF_i )
	begin
	rl_a67_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a67_t4 = ( ( { 9{ FF_i } } & rl_a67_t5 )
		| ( { 9{ rl_a67_t4_c1 } } & rl_a67_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_9 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h01 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h02 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h03 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h04 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h05 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h06 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h07 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h08 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h09 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h0a :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h0b :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h0c :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h0d :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h0e :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h0f :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h10 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h11 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h12 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h13 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h14 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h15 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h16 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h17 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h18 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h19 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h1a :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h1b :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h1c :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h1d :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h1e :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h1f :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h20 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h21 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h22 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h23 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h24 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h25 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h26 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h27 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h28 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h29 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h2a :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h2b :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h2c :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h2d :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h2e :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h2f :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h30 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h31 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h32 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h33 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h34 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h35 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h36 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h37 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h38 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h39 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h3a :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h3b :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h3c :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h3d :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h3e :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h3f :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h40 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h41 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h42 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h43 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h44 :
		rl_a68_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h45 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h46 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h47 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h48 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h49 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h4a :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h4b :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h4c :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h4d :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h4e :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h4f :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h50 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h51 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h52 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h53 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h54 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h55 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h56 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h57 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h58 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h59 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h5a :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h5b :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h5c :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h5d :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h5e :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h5f :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h60 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h61 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h62 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h63 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h64 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h65 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h66 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h67 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h68 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h69 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h6a :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h6b :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h6c :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h6d :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h6e :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h6f :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h70 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h71 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h72 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h73 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h74 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h75 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h76 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h77 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h78 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h79 :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h7a :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h7b :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h7c :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h7d :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h7e :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	7'h7f :
		rl_a68_t4_t1 = RG_quantized_block_rl_9 ;
	default :
		rl_a68_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a68_t4_t1 or rl_a68_t5 or FF_i )
	begin
	rl_a68_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a68_t4 = ( ( { 9{ FF_i } } & rl_a68_t5 )
		| ( { 9{ rl_a68_t4_c1 } } & rl_a68_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_10 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h01 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h02 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h03 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h04 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h05 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h06 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h07 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h08 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h09 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h0a :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h0b :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h0c :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h0d :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h0e :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h0f :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h10 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h11 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h12 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h13 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h14 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h15 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h16 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h17 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h18 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h19 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h1a :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h1b :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h1c :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h1d :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h1e :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h1f :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h20 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h21 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h22 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h23 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h24 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h25 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h26 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h27 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h28 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h29 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h2a :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h2b :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h2c :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h2d :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h2e :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h2f :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h30 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h31 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h32 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h33 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h34 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h35 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h36 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h37 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h38 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h39 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h3a :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h3b :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h3c :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h3d :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h3e :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h3f :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h40 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h41 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h42 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h43 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h44 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h45 :
		rl_a69_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h46 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h47 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h48 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h49 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h4a :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h4b :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h4c :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h4d :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h4e :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h4f :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h50 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h51 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h52 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h53 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h54 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h55 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h56 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h57 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h58 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h59 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h5a :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h5b :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h5c :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h5d :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h5e :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h5f :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h60 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h61 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h62 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h63 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h64 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h65 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h66 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h67 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h68 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h69 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h6a :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h6b :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h6c :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h6d :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h6e :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h6f :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h70 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h71 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h72 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h73 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h74 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h75 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h76 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h77 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h78 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h79 :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h7a :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h7b :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h7c :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h7d :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h7e :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	7'h7f :
		rl_a69_t4_t1 = RG_quantized_block_rl_10 ;
	default :
		rl_a69_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a69_t4_t1 or rl_a69_t5 or FF_i )
	begin
	rl_a69_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a69_t4 = ( ( { 9{ FF_i } } & rl_a69_t5 )
		| ( { 9{ rl_a69_t4_c1 } } & rl_a69_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_11 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h01 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h02 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h03 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h04 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h05 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h06 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h07 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h08 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h09 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h0a :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h0b :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h0c :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h0d :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h0e :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h0f :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h10 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h11 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h12 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h13 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h14 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h15 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h16 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h17 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h18 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h19 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h1a :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h1b :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h1c :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h1d :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h1e :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h1f :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h20 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h21 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h22 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h23 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h24 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h25 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h26 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h27 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h28 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h29 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h2a :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h2b :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h2c :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h2d :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h2e :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h2f :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h30 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h31 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h32 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h33 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h34 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h35 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h36 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h37 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h38 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h39 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h3a :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h3b :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h3c :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h3d :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h3e :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h3f :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h40 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h41 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h42 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h43 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h44 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h45 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h46 :
		rl_a70_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h47 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h48 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h49 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h4a :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h4b :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h4c :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h4d :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h4e :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h4f :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h50 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h51 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h52 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h53 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h54 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h55 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h56 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h57 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h58 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h59 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h5a :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h5b :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h5c :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h5d :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h5e :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h5f :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h60 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h61 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h62 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h63 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h64 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h65 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h66 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h67 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h68 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h69 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h6a :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h6b :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h6c :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h6d :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h6e :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h6f :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h70 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h71 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h72 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h73 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h74 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h75 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h76 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h77 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h78 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h79 :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h7a :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h7b :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h7c :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h7d :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h7e :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	7'h7f :
		rl_a70_t4_t1 = RG_quantized_block_rl_11 ;
	default :
		rl_a70_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a70_t4_t1 or rl_a70_t5 or FF_i )
	begin
	rl_a70_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a70_t4 = ( ( { 9{ FF_i } } & rl_a70_t5 )
		| ( { 9{ rl_a70_t4_c1 } } & rl_a70_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_12 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h01 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h02 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h03 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h04 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h05 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h06 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h07 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h08 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h09 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h0a :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h0b :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h0c :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h0d :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h0e :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h0f :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h10 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h11 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h12 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h13 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h14 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h15 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h16 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h17 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h18 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h19 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h1a :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h1b :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h1c :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h1d :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h1e :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h1f :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h20 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h21 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h22 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h23 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h24 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h25 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h26 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h27 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h28 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h29 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h2a :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h2b :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h2c :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h2d :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h2e :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h2f :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h30 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h31 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h32 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h33 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h34 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h35 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h36 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h37 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h38 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h39 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h3a :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h3b :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h3c :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h3d :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h3e :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h3f :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h40 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h41 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h42 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h43 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h44 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h45 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h46 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h47 :
		rl_a71_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h48 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h49 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h4a :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h4b :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h4c :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h4d :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h4e :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h4f :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h50 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h51 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h52 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h53 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h54 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h55 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h56 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h57 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h58 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h59 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h5a :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h5b :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h5c :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h5d :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h5e :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h5f :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h60 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h61 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h62 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h63 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h64 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h65 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h66 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h67 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h68 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h69 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h6a :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h6b :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h6c :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h6d :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h6e :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h6f :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h70 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h71 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h72 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h73 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h74 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h75 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h76 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h77 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h78 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h79 :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h7a :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h7b :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h7c :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h7d :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h7e :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	7'h7f :
		rl_a71_t4_t1 = RG_quantized_block_rl_12 ;
	default :
		rl_a71_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a71_t4_t1 or rl_a71_t5 or FF_i )
	begin
	rl_a71_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a71_t4 = ( ( { 9{ FF_i } } & rl_a71_t5 )
		| ( { 9{ rl_a71_t4_c1 } } & rl_a71_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_13 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h01 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h02 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h03 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h04 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h05 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h06 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h07 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h08 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h09 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h0a :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h0b :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h0c :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h0d :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h0e :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h0f :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h10 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h11 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h12 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h13 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h14 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h15 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h16 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h17 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h18 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h19 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h1a :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h1b :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h1c :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h1d :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h1e :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h1f :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h20 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h21 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h22 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h23 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h24 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h25 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h26 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h27 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h28 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h29 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h2a :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h2b :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h2c :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h2d :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h2e :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h2f :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h30 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h31 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h32 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h33 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h34 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h35 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h36 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h37 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h38 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h39 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h3a :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h3b :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h3c :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h3d :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h3e :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h3f :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h40 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h41 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h42 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h43 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h44 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h45 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h46 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h47 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h48 :
		rl_a72_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h49 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h4a :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h4b :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h4c :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h4d :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h4e :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h4f :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h50 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h51 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h52 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h53 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h54 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h55 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h56 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h57 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h58 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h59 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h5a :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h5b :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h5c :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h5d :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h5e :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h5f :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h60 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h61 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h62 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h63 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h64 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h65 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h66 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h67 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h68 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h69 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h6a :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h6b :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h6c :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h6d :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h6e :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h6f :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h70 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h71 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h72 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h73 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h74 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h75 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h76 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h77 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h78 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h79 :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h7a :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h7b :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h7c :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h7d :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h7e :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	7'h7f :
		rl_a72_t4_t1 = RG_quantized_block_rl_13 ;
	default :
		rl_a72_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a72_t4_t1 or rl_a72_t5 or FF_i )
	begin
	rl_a72_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a72_t4 = ( ( { 9{ FF_i } } & rl_a72_t5 )
		| ( { 9{ rl_a72_t4_c1 } } & rl_a72_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_14 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h01 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h02 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h03 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h04 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h05 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h06 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h07 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h08 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h09 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h0a :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h0b :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h0c :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h0d :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h0e :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h0f :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h10 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h11 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h12 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h13 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h14 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h15 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h16 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h17 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h18 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h19 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h1a :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h1b :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h1c :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h1d :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h1e :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h1f :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h20 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h21 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h22 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h23 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h24 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h25 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h26 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h27 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h28 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h29 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h2a :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h2b :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h2c :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h2d :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h2e :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h2f :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h30 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h31 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h32 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h33 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h34 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h35 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h36 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h37 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h38 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h39 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h3a :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h3b :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h3c :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h3d :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h3e :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h3f :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h40 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h41 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h42 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h43 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h44 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h45 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h46 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h47 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h48 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h49 :
		rl_a73_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h4a :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h4b :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h4c :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h4d :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h4e :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h4f :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h50 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h51 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h52 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h53 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h54 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h55 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h56 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h57 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h58 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h59 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h5a :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h5b :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h5c :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h5d :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h5e :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h5f :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h60 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h61 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h62 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h63 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h64 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h65 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h66 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h67 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h68 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h69 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h6a :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h6b :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h6c :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h6d :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h6e :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h6f :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h70 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h71 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h72 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h73 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h74 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h75 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h76 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h77 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h78 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h79 :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h7a :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h7b :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h7c :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h7d :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h7e :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	7'h7f :
		rl_a73_t4_t1 = RG_quantized_block_rl_14 ;
	default :
		rl_a73_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a73_t4_t1 or rl_a73_t5 or FF_i )
	begin
	rl_a73_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a73_t4 = ( ( { 9{ FF_i } } & rl_a73_t5 )
		| ( { 9{ rl_a73_t4_c1 } } & rl_a73_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_15 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h01 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h02 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h03 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h04 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h05 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h06 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h07 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h08 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h09 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h0a :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h0b :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h0c :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h0d :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h0e :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h0f :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h10 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h11 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h12 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h13 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h14 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h15 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h16 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h17 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h18 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h19 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h1a :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h1b :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h1c :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h1d :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h1e :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h1f :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h20 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h21 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h22 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h23 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h24 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h25 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h26 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h27 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h28 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h29 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h2a :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h2b :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h2c :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h2d :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h2e :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h2f :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h30 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h31 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h32 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h33 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h34 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h35 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h36 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h37 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h38 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h39 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h3a :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h3b :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h3c :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h3d :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h3e :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h3f :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h40 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h41 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h42 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h43 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h44 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h45 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h46 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h47 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h48 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h49 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h4a :
		rl_a74_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h4b :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h4c :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h4d :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h4e :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h4f :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h50 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h51 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h52 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h53 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h54 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h55 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h56 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h57 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h58 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h59 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h5a :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h5b :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h5c :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h5d :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h5e :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h5f :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h60 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h61 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h62 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h63 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h64 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h65 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h66 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h67 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h68 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h69 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h6a :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h6b :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h6c :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h6d :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h6e :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h6f :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h70 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h71 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h72 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h73 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h74 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h75 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h76 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h77 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h78 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h79 :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h7a :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h7b :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h7c :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h7d :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h7e :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	7'h7f :
		rl_a74_t4_t1 = RG_quantized_block_rl_15 ;
	default :
		rl_a74_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a74_t4_t1 or rl_a74_t5 or FF_i )
	begin
	rl_a74_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a74_t4 = ( ( { 9{ FF_i } } & rl_a74_t5 )
		| ( { 9{ rl_a74_t4_c1 } } & rl_a74_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_16 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h01 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h02 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h03 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h04 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h05 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h06 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h07 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h08 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h09 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h0a :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h0b :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h0c :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h0d :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h0e :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h0f :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h10 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h11 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h12 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h13 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h14 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h15 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h16 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h17 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h18 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h19 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h1a :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h1b :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h1c :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h1d :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h1e :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h1f :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h20 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h21 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h22 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h23 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h24 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h25 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h26 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h27 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h28 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h29 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h2a :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h2b :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h2c :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h2d :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h2e :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h2f :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h30 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h31 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h32 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h33 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h34 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h35 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h36 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h37 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h38 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h39 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h3a :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h3b :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h3c :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h3d :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h3e :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h3f :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h40 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h41 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h42 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h43 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h44 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h45 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h46 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h47 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h48 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h49 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h4a :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h4b :
		rl_a75_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h4c :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h4d :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h4e :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h4f :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h50 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h51 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h52 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h53 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h54 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h55 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h56 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h57 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h58 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h59 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h5a :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h5b :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h5c :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h5d :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h5e :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h5f :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h60 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h61 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h62 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h63 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h64 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h65 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h66 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h67 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h68 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h69 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h6a :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h6b :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h6c :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h6d :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h6e :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h6f :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h70 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h71 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h72 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h73 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h74 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h75 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h76 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h77 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h78 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h79 :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h7a :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h7b :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h7c :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h7d :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h7e :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	7'h7f :
		rl_a75_t4_t1 = RG_quantized_block_rl_16 ;
	default :
		rl_a75_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a75_t4_t1 or rl_a75_t5 or FF_i )
	begin
	rl_a75_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a75_t4 = ( ( { 9{ FF_i } } & rl_a75_t5 )
		| ( { 9{ rl_a75_t4_c1 } } & rl_a75_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_17 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h01 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h02 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h03 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h04 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h05 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h06 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h07 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h08 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h09 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h0a :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h0b :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h0c :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h0d :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h0e :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h0f :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h10 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h11 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h12 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h13 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h14 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h15 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h16 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h17 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h18 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h19 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h1a :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h1b :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h1c :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h1d :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h1e :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h1f :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h20 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h21 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h22 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h23 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h24 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h25 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h26 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h27 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h28 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h29 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h2a :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h2b :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h2c :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h2d :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h2e :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h2f :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h30 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h31 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h32 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h33 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h34 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h35 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h36 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h37 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h38 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h39 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h3a :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h3b :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h3c :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h3d :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h3e :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h3f :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h40 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h41 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h42 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h43 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h44 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h45 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h46 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h47 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h48 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h49 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h4a :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h4b :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h4c :
		rl_a76_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h4d :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h4e :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h4f :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h50 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h51 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h52 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h53 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h54 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h55 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h56 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h57 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h58 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h59 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h5a :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h5b :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h5c :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h5d :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h5e :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h5f :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h60 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h61 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h62 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h63 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h64 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h65 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h66 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h67 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h68 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h69 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h6a :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h6b :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h6c :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h6d :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h6e :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h6f :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h70 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h71 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h72 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h73 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h74 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h75 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h76 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h77 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h78 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h79 :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h7a :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h7b :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h7c :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h7d :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h7e :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	7'h7f :
		rl_a76_t4_t1 = RG_quantized_block_rl_17 ;
	default :
		rl_a76_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a76_t4_t1 or rl_a76_t5 or FF_i )
	begin
	rl_a76_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a76_t4 = ( ( { 9{ FF_i } } & rl_a76_t5 )
		| ( { 9{ rl_a76_t4_c1 } } & rl_a76_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_18 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h01 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h02 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h03 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h04 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h05 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h06 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h07 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h08 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h09 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h0a :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h0b :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h0c :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h0d :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h0e :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h0f :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h10 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h11 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h12 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h13 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h14 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h15 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h16 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h17 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h18 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h19 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h1a :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h1b :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h1c :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h1d :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h1e :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h1f :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h20 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h21 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h22 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h23 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h24 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h25 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h26 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h27 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h28 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h29 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h2a :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h2b :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h2c :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h2d :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h2e :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h2f :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h30 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h31 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h32 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h33 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h34 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h35 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h36 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h37 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h38 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h39 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h3a :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h3b :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h3c :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h3d :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h3e :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h3f :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h40 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h41 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h42 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h43 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h44 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h45 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h46 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h47 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h48 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h49 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h4a :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h4b :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h4c :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h4d :
		rl_a77_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h4e :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h4f :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h50 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h51 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h52 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h53 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h54 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h55 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h56 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h57 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h58 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h59 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h5a :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h5b :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h5c :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h5d :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h5e :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h5f :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h60 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h61 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h62 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h63 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h64 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h65 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h66 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h67 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h68 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h69 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h6a :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h6b :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h6c :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h6d :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h6e :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h6f :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h70 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h71 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h72 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h73 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h74 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h75 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h76 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h77 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h78 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h79 :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h7a :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h7b :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h7c :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h7d :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h7e :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	7'h7f :
		rl_a77_t4_t1 = RG_quantized_block_rl_18 ;
	default :
		rl_a77_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a77_t4_t1 or rl_a77_t5 or FF_i )
	begin
	rl_a77_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a77_t4 = ( ( { 9{ FF_i } } & rl_a77_t5 )
		| ( { 9{ rl_a77_t4_c1 } } & rl_a77_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_19 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h01 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h02 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h03 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h04 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h05 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h06 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h07 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h08 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h09 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h0a :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h0b :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h0c :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h0d :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h0e :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h0f :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h10 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h11 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h12 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h13 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h14 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h15 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h16 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h17 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h18 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h19 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h1a :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h1b :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h1c :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h1d :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h1e :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h1f :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h20 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h21 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h22 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h23 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h24 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h25 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h26 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h27 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h28 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h29 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h2a :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h2b :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h2c :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h2d :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h2e :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h2f :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h30 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h31 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h32 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h33 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h34 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h35 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h36 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h37 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h38 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h39 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h3a :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h3b :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h3c :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h3d :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h3e :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h3f :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h40 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h41 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h42 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h43 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h44 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h45 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h46 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h47 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h48 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h49 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h4a :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h4b :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h4c :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h4d :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h4e :
		rl_a78_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h4f :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h50 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h51 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h52 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h53 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h54 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h55 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h56 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h57 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h58 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h59 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h5a :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h5b :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h5c :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h5d :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h5e :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h5f :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h60 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h61 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h62 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h63 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h64 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h65 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h66 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h67 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h68 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h69 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h6a :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h6b :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h6c :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h6d :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h6e :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h6f :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h70 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h71 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h72 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h73 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h74 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h75 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h76 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h77 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h78 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h79 :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h7a :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h7b :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h7c :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h7d :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h7e :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	7'h7f :
		rl_a78_t4_t1 = RG_quantized_block_rl_19 ;
	default :
		rl_a78_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a78_t4_t1 or rl_a78_t5 or FF_i )
	begin
	rl_a78_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a78_t4 = ( ( { 9{ FF_i } } & rl_a78_t5 )
		| ( { 9{ rl_a78_t4_c1 } } & rl_a78_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_20 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h01 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h02 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h03 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h04 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h05 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h06 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h07 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h08 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h09 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h0a :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h0b :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h0c :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h0d :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h0e :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h0f :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h10 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h11 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h12 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h13 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h14 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h15 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h16 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h17 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h18 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h19 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h1a :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h1b :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h1c :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h1d :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h1e :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h1f :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h20 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h21 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h22 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h23 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h24 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h25 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h26 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h27 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h28 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h29 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h2a :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h2b :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h2c :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h2d :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h2e :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h2f :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h30 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h31 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h32 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h33 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h34 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h35 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h36 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h37 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h38 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h39 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h3a :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h3b :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h3c :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h3d :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h3e :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h3f :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h40 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h41 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h42 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h43 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h44 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h45 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h46 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h47 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h48 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h49 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h4a :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h4b :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h4c :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h4d :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h4e :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h4f :
		rl_a79_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h50 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h51 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h52 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h53 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h54 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h55 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h56 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h57 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h58 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h59 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h5a :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h5b :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h5c :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h5d :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h5e :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h5f :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h60 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h61 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h62 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h63 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h64 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h65 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h66 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h67 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h68 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h69 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h6a :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h6b :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h6c :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h6d :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h6e :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h6f :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h70 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h71 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h72 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h73 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h74 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h75 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h76 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h77 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h78 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h79 :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h7a :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h7b :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h7c :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h7d :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h7e :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	7'h7f :
		rl_a79_t4_t1 = RG_quantized_block_rl_20 ;
	default :
		rl_a79_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a79_t4_t1 or rl_a79_t5 or FF_i )
	begin
	rl_a79_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a79_t4 = ( ( { 9{ FF_i } } & rl_a79_t5 )
		| ( { 9{ rl_a79_t4_c1 } } & rl_a79_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_21 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h01 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h02 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h03 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h04 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h05 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h06 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h07 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h08 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h09 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h0a :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h0b :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h0c :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h0d :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h0e :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h0f :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h10 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h11 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h12 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h13 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h14 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h15 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h16 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h17 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h18 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h19 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h1a :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h1b :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h1c :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h1d :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h1e :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h1f :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h20 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h21 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h22 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h23 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h24 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h25 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h26 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h27 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h28 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h29 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h2a :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h2b :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h2c :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h2d :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h2e :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h2f :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h30 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h31 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h32 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h33 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h34 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h35 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h36 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h37 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h38 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h39 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h3a :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h3b :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h3c :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h3d :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h3e :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h3f :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h40 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h41 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h42 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h43 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h44 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h45 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h46 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h47 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h48 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h49 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h4a :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h4b :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h4c :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h4d :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h4e :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h4f :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h50 :
		rl_a80_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h51 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h52 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h53 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h54 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h55 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h56 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h57 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h58 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h59 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h5a :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h5b :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h5c :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h5d :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h5e :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h5f :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h60 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h61 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h62 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h63 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h64 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h65 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h66 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h67 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h68 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h69 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h6a :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h6b :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h6c :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h6d :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h6e :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h6f :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h70 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h71 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h72 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h73 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h74 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h75 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h76 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h77 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h78 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h79 :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h7a :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h7b :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h7c :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h7d :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h7e :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	7'h7f :
		rl_a80_t4_t1 = RG_quantized_block_rl_21 ;
	default :
		rl_a80_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a80_t4_t1 or rl_a80_t5 or FF_i )
	begin
	rl_a80_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a80_t4 = ( ( { 9{ FF_i } } & rl_a80_t5 )
		| ( { 9{ rl_a80_t4_c1 } } & rl_a80_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_22 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h01 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h02 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h03 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h04 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h05 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h06 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h07 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h08 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h09 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h0a :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h0b :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h0c :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h0d :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h0e :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h0f :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h10 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h11 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h12 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h13 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h14 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h15 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h16 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h17 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h18 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h19 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h1a :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h1b :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h1c :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h1d :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h1e :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h1f :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h20 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h21 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h22 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h23 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h24 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h25 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h26 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h27 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h28 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h29 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h2a :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h2b :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h2c :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h2d :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h2e :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h2f :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h30 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h31 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h32 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h33 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h34 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h35 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h36 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h37 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h38 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h39 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h3a :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h3b :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h3c :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h3d :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h3e :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h3f :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h40 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h41 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h42 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h43 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h44 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h45 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h46 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h47 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h48 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h49 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h4a :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h4b :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h4c :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h4d :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h4e :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h4f :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h50 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h51 :
		rl_a81_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h52 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h53 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h54 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h55 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h56 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h57 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h58 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h59 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h5a :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h5b :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h5c :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h5d :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h5e :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h5f :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h60 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h61 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h62 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h63 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h64 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h65 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h66 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h67 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h68 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h69 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h6a :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h6b :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h6c :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h6d :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h6e :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h6f :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h70 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h71 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h72 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h73 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h74 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h75 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h76 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h77 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h78 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h79 :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h7a :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h7b :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h7c :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h7d :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h7e :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	7'h7f :
		rl_a81_t4_t1 = RG_quantized_block_rl_22 ;
	default :
		rl_a81_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a81_t4_t1 or rl_a81_t5 or FF_i )
	begin
	rl_a81_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a81_t4 = ( ( { 9{ FF_i } } & rl_a81_t5 )
		| ( { 9{ rl_a81_t4_c1 } } & rl_a81_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_23 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h01 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h02 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h03 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h04 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h05 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h06 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h07 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h08 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h09 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h0a :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h0b :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h0c :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h0d :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h0e :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h0f :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h10 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h11 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h12 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h13 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h14 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h15 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h16 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h17 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h18 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h19 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h1a :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h1b :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h1c :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h1d :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h1e :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h1f :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h20 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h21 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h22 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h23 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h24 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h25 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h26 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h27 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h28 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h29 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h2a :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h2b :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h2c :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h2d :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h2e :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h2f :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h30 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h31 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h32 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h33 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h34 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h35 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h36 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h37 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h38 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h39 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h3a :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h3b :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h3c :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h3d :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h3e :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h3f :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h40 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h41 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h42 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h43 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h44 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h45 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h46 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h47 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h48 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h49 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h4a :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h4b :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h4c :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h4d :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h4e :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h4f :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h50 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h51 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h52 :
		rl_a82_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h53 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h54 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h55 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h56 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h57 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h58 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h59 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h5a :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h5b :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h5c :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h5d :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h5e :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h5f :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h60 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h61 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h62 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h63 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h64 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h65 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h66 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h67 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h68 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h69 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h6a :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h6b :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h6c :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h6d :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h6e :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h6f :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h70 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h71 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h72 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h73 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h74 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h75 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h76 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h77 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h78 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h79 :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h7a :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h7b :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h7c :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h7d :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h7e :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	7'h7f :
		rl_a82_t4_t1 = RG_quantized_block_rl_23 ;
	default :
		rl_a82_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a82_t4_t1 or rl_a82_t5 or FF_i )
	begin
	rl_a82_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a82_t4 = ( ( { 9{ FF_i } } & rl_a82_t5 )
		| ( { 9{ rl_a82_t4_c1 } } & rl_a82_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_24 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h01 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h02 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h03 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h04 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h05 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h06 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h07 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h08 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h09 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h0a :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h0b :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h0c :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h0d :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h0e :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h0f :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h10 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h11 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h12 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h13 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h14 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h15 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h16 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h17 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h18 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h19 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h1a :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h1b :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h1c :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h1d :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h1e :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h1f :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h20 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h21 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h22 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h23 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h24 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h25 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h26 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h27 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h28 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h29 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h2a :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h2b :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h2c :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h2d :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h2e :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h2f :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h30 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h31 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h32 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h33 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h34 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h35 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h36 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h37 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h38 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h39 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h3a :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h3b :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h3c :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h3d :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h3e :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h3f :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h40 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h41 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h42 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h43 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h44 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h45 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h46 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h47 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h48 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h49 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h4a :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h4b :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h4c :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h4d :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h4e :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h4f :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h50 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h51 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h52 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h53 :
		rl_a83_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h54 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h55 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h56 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h57 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h58 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h59 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h5a :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h5b :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h5c :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h5d :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h5e :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h5f :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h60 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h61 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h62 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h63 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h64 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h65 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h66 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h67 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h68 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h69 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h6a :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h6b :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h6c :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h6d :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h6e :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h6f :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h70 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h71 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h72 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h73 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h74 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h75 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h76 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h77 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h78 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h79 :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h7a :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h7b :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h7c :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h7d :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h7e :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	7'h7f :
		rl_a83_t4_t1 = RG_quantized_block_rl_24 ;
	default :
		rl_a83_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a83_t4_t1 or rl_a83_t5 or FF_i )
	begin
	rl_a83_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a83_t4 = ( ( { 9{ FF_i } } & rl_a83_t5 )
		| ( { 9{ rl_a83_t4_c1 } } & rl_a83_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_25 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h01 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h02 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h03 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h04 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h05 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h06 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h07 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h08 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h09 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h0a :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h0b :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h0c :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h0d :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h0e :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h0f :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h10 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h11 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h12 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h13 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h14 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h15 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h16 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h17 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h18 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h19 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h1a :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h1b :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h1c :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h1d :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h1e :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h1f :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h20 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h21 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h22 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h23 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h24 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h25 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h26 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h27 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h28 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h29 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h2a :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h2b :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h2c :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h2d :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h2e :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h2f :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h30 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h31 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h32 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h33 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h34 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h35 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h36 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h37 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h38 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h39 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h3a :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h3b :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h3c :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h3d :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h3e :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h3f :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h40 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h41 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h42 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h43 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h44 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h45 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h46 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h47 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h48 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h49 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h4a :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h4b :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h4c :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h4d :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h4e :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h4f :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h50 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h51 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h52 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h53 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h54 :
		rl_a84_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h55 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h56 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h57 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h58 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h59 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h5a :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h5b :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h5c :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h5d :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h5e :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h5f :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h60 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h61 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h62 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h63 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h64 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h65 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h66 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h67 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h68 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h69 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h6a :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h6b :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h6c :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h6d :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h6e :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h6f :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h70 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h71 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h72 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h73 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h74 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h75 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h76 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h77 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h78 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h79 :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h7a :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h7b :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h7c :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h7d :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h7e :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	7'h7f :
		rl_a84_t4_t1 = RG_quantized_block_rl_25 ;
	default :
		rl_a84_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a84_t4_t1 or rl_a84_t5 or FF_i )
	begin
	rl_a84_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a84_t4 = ( ( { 9{ FF_i } } & rl_a84_t5 )
		| ( { 9{ rl_a84_t4_c1 } } & rl_a84_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_26 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h01 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h02 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h03 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h04 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h05 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h06 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h07 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h08 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h09 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h0a :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h0b :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h0c :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h0d :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h0e :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h0f :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h10 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h11 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h12 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h13 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h14 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h15 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h16 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h17 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h18 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h19 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h1a :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h1b :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h1c :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h1d :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h1e :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h1f :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h20 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h21 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h22 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h23 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h24 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h25 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h26 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h27 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h28 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h29 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h2a :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h2b :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h2c :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h2d :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h2e :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h2f :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h30 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h31 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h32 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h33 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h34 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h35 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h36 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h37 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h38 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h39 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h3a :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h3b :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h3c :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h3d :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h3e :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h3f :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h40 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h41 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h42 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h43 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h44 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h45 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h46 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h47 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h48 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h49 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h4a :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h4b :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h4c :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h4d :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h4e :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h4f :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h50 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h51 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h52 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h53 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h54 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h55 :
		rl_a85_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h56 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h57 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h58 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h59 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h5a :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h5b :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h5c :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h5d :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h5e :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h5f :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h60 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h61 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h62 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h63 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h64 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h65 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h66 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h67 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h68 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h69 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h6a :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h6b :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h6c :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h6d :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h6e :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h6f :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h70 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h71 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h72 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h73 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h74 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h75 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h76 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h77 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h78 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h79 :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h7a :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h7b :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h7c :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h7d :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h7e :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	7'h7f :
		rl_a85_t4_t1 = RG_quantized_block_rl_26 ;
	default :
		rl_a85_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a85_t4_t1 or rl_a85_t5 or FF_i )
	begin
	rl_a85_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a85_t4 = ( ( { 9{ FF_i } } & rl_a85_t5 )
		| ( { 9{ rl_a85_t4_c1 } } & rl_a85_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_27 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h01 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h02 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h03 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h04 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h05 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h06 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h07 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h08 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h09 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h0a :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h0b :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h0c :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h0d :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h0e :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h0f :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h10 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h11 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h12 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h13 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h14 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h15 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h16 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h17 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h18 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h19 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h1a :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h1b :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h1c :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h1d :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h1e :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h1f :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h20 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h21 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h22 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h23 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h24 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h25 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h26 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h27 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h28 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h29 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h2a :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h2b :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h2c :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h2d :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h2e :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h2f :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h30 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h31 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h32 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h33 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h34 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h35 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h36 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h37 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h38 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h39 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h3a :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h3b :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h3c :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h3d :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h3e :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h3f :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h40 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h41 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h42 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h43 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h44 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h45 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h46 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h47 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h48 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h49 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h4a :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h4b :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h4c :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h4d :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h4e :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h4f :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h50 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h51 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h52 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h53 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h54 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h55 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h56 :
		rl_a86_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h57 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h58 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h59 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h5a :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h5b :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h5c :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h5d :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h5e :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h5f :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h60 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h61 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h62 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h63 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h64 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h65 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h66 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h67 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h68 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h69 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h6a :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h6b :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h6c :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h6d :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h6e :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h6f :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h70 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h71 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h72 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h73 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h74 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h75 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h76 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h77 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h78 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h79 :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h7a :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h7b :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h7c :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h7d :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h7e :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	7'h7f :
		rl_a86_t4_t1 = RG_quantized_block_rl_27 ;
	default :
		rl_a86_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a86_t4_t1 or rl_a86_t5 or FF_i )
	begin
	rl_a86_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a86_t4 = ( ( { 9{ FF_i } } & rl_a86_t5 )
		| ( { 9{ rl_a86_t4_c1 } } & rl_a86_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_28 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h01 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h02 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h03 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h04 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h05 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h06 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h07 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h08 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h09 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h0a :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h0b :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h0c :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h0d :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h0e :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h0f :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h10 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h11 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h12 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h13 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h14 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h15 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h16 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h17 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h18 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h19 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h1a :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h1b :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h1c :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h1d :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h1e :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h1f :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h20 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h21 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h22 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h23 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h24 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h25 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h26 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h27 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h28 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h29 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h2a :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h2b :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h2c :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h2d :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h2e :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h2f :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h30 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h31 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h32 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h33 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h34 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h35 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h36 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h37 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h38 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h39 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h3a :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h3b :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h3c :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h3d :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h3e :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h3f :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h40 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h41 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h42 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h43 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h44 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h45 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h46 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h47 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h48 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h49 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h4a :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h4b :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h4c :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h4d :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h4e :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h4f :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h50 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h51 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h52 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h53 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h54 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h55 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h56 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h57 :
		rl_a87_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h58 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h59 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h5a :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h5b :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h5c :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h5d :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h5e :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h5f :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h60 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h61 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h62 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h63 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h64 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h65 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h66 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h67 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h68 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h69 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h6a :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h6b :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h6c :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h6d :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h6e :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h6f :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h70 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h71 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h72 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h73 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h74 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h75 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h76 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h77 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h78 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h79 :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h7a :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h7b :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h7c :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h7d :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h7e :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	7'h7f :
		rl_a87_t4_t1 = RG_quantized_block_rl_28 ;
	default :
		rl_a87_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a87_t4_t1 or rl_a87_t5 or FF_i )
	begin
	rl_a87_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a87_t4 = ( ( { 9{ FF_i } } & rl_a87_t5 )
		| ( { 9{ rl_a87_t4_c1 } } & rl_a87_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_29 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h01 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h02 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h03 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h04 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h05 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h06 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h07 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h08 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h09 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h0a :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h0b :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h0c :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h0d :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h0e :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h0f :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h10 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h11 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h12 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h13 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h14 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h15 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h16 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h17 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h18 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h19 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h1a :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h1b :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h1c :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h1d :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h1e :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h1f :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h20 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h21 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h22 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h23 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h24 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h25 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h26 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h27 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h28 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h29 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h2a :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h2b :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h2c :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h2d :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h2e :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h2f :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h30 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h31 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h32 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h33 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h34 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h35 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h36 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h37 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h38 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h39 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h3a :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h3b :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h3c :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h3d :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h3e :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h3f :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h40 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h41 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h42 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h43 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h44 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h45 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h46 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h47 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h48 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h49 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h4a :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h4b :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h4c :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h4d :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h4e :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h4f :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h50 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h51 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h52 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h53 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h54 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h55 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h56 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h57 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h58 :
		rl_a88_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h59 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h5a :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h5b :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h5c :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h5d :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h5e :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h5f :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h60 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h61 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h62 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h63 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h64 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h65 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h66 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h67 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h68 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h69 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h6a :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h6b :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h6c :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h6d :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h6e :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h6f :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h70 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h71 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h72 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h73 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h74 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h75 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h76 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h77 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h78 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h79 :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h7a :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h7b :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h7c :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h7d :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h7e :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	7'h7f :
		rl_a88_t4_t1 = RG_quantized_block_rl_29 ;
	default :
		rl_a88_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a88_t4_t1 or rl_a88_t5 or FF_i )
	begin
	rl_a88_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a88_t4 = ( ( { 9{ FF_i } } & rl_a88_t5 )
		| ( { 9{ rl_a88_t4_c1 } } & rl_a88_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_30 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h01 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h02 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h03 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h04 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h05 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h06 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h07 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h08 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h09 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h0a :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h0b :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h0c :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h0d :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h0e :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h0f :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h10 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h11 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h12 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h13 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h14 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h15 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h16 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h17 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h18 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h19 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h1a :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h1b :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h1c :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h1d :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h1e :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h1f :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h20 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h21 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h22 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h23 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h24 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h25 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h26 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h27 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h28 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h29 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h2a :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h2b :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h2c :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h2d :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h2e :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h2f :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h30 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h31 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h32 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h33 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h34 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h35 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h36 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h37 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h38 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h39 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h3a :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h3b :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h3c :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h3d :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h3e :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h3f :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h40 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h41 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h42 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h43 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h44 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h45 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h46 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h47 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h48 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h49 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h4a :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h4b :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h4c :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h4d :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h4e :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h4f :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h50 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h51 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h52 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h53 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h54 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h55 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h56 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h57 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h58 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h59 :
		rl_a89_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h5a :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h5b :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h5c :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h5d :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h5e :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h5f :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h60 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h61 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h62 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h63 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h64 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h65 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h66 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h67 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h68 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h69 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h6a :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h6b :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h6c :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h6d :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h6e :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h6f :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h70 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h71 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h72 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h73 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h74 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h75 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h76 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h77 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h78 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h79 :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h7a :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h7b :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h7c :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h7d :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h7e :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	7'h7f :
		rl_a89_t4_t1 = RG_quantized_block_rl_30 ;
	default :
		rl_a89_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a89_t4_t1 or rl_a89_t5 or FF_i )
	begin
	rl_a89_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a89_t4 = ( ( { 9{ FF_i } } & rl_a89_t5 )
		| ( { 9{ rl_a89_t4_c1 } } & rl_a89_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_31 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h01 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h02 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h03 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h04 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h05 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h06 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h07 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h08 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h09 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h0a :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h0b :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h0c :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h0d :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h0e :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h0f :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h10 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h11 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h12 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h13 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h14 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h15 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h16 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h17 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h18 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h19 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h1a :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h1b :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h1c :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h1d :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h1e :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h1f :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h20 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h21 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h22 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h23 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h24 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h25 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h26 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h27 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h28 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h29 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h2a :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h2b :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h2c :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h2d :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h2e :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h2f :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h30 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h31 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h32 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h33 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h34 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h35 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h36 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h37 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h38 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h39 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h3a :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h3b :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h3c :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h3d :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h3e :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h3f :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h40 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h41 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h42 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h43 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h44 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h45 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h46 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h47 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h48 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h49 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h4a :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h4b :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h4c :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h4d :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h4e :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h4f :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h50 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h51 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h52 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h53 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h54 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h55 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h56 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h57 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h58 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h59 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h5a :
		rl_a90_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h5b :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h5c :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h5d :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h5e :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h5f :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h60 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h61 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h62 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h63 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h64 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h65 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h66 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h67 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h68 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h69 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h6a :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h6b :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h6c :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h6d :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h6e :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h6f :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h70 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h71 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h72 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h73 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h74 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h75 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h76 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h77 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h78 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h79 :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h7a :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h7b :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h7c :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h7d :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h7e :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	7'h7f :
		rl_a90_t4_t1 = RG_quantized_block_rl_31 ;
	default :
		rl_a90_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a90_t4_t1 or rl_a90_t5 or FF_i )
	begin
	rl_a90_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a90_t4 = ( ( { 9{ FF_i } } & rl_a90_t5 )
		| ( { 9{ rl_a90_t4_c1 } } & rl_a90_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_32 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h01 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h02 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h03 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h04 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h05 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h06 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h07 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h08 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h09 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h0a :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h0b :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h0c :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h0d :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h0e :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h0f :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h10 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h11 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h12 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h13 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h14 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h15 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h16 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h17 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h18 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h19 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h1a :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h1b :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h1c :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h1d :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h1e :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h1f :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h20 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h21 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h22 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h23 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h24 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h25 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h26 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h27 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h28 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h29 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h2a :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h2b :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h2c :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h2d :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h2e :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h2f :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h30 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h31 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h32 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h33 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h34 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h35 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h36 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h37 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h38 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h39 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h3a :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h3b :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h3c :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h3d :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h3e :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h3f :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h40 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h41 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h42 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h43 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h44 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h45 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h46 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h47 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h48 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h49 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h4a :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h4b :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h4c :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h4d :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h4e :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h4f :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h50 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h51 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h52 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h53 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h54 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h55 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h56 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h57 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h58 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h59 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h5a :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h5b :
		rl_a91_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h5c :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h5d :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h5e :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h5f :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h60 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h61 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h62 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h63 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h64 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h65 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h66 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h67 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h68 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h69 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h6a :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h6b :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h6c :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h6d :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h6e :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h6f :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h70 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h71 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h72 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h73 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h74 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h75 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h76 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h77 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h78 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h79 :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h7a :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h7b :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h7c :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h7d :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h7e :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	7'h7f :
		rl_a91_t4_t1 = RG_quantized_block_rl_32 ;
	default :
		rl_a91_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a91_t4_t1 or rl_a91_t5 or FF_i )
	begin
	rl_a91_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a91_t4 = ( ( { 9{ FF_i } } & rl_a91_t5 )
		| ( { 9{ rl_a91_t4_c1 } } & rl_a91_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_33 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h01 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h02 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h03 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h04 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h05 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h06 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h07 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h08 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h09 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h0a :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h0b :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h0c :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h0d :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h0e :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h0f :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h10 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h11 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h12 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h13 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h14 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h15 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h16 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h17 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h18 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h19 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h1a :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h1b :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h1c :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h1d :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h1e :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h1f :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h20 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h21 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h22 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h23 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h24 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h25 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h26 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h27 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h28 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h29 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h2a :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h2b :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h2c :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h2d :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h2e :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h2f :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h30 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h31 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h32 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h33 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h34 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h35 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h36 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h37 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h38 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h39 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h3a :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h3b :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h3c :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h3d :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h3e :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h3f :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h40 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h41 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h42 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h43 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h44 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h45 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h46 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h47 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h48 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h49 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h4a :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h4b :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h4c :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h4d :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h4e :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h4f :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h50 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h51 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h52 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h53 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h54 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h55 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h56 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h57 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h58 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h59 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h5a :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h5b :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h5c :
		rl_a92_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h5d :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h5e :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h5f :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h60 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h61 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h62 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h63 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h64 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h65 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h66 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h67 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h68 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h69 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h6a :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h6b :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h6c :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h6d :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h6e :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h6f :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h70 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h71 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h72 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h73 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h74 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h75 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h76 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h77 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h78 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h79 :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h7a :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h7b :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h7c :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h7d :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h7e :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	7'h7f :
		rl_a92_t4_t1 = RG_quantized_block_rl_33 ;
	default :
		rl_a92_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a92_t4_t1 or rl_a92_t5 or FF_i )
	begin
	rl_a92_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a92_t4 = ( ( { 9{ FF_i } } & rl_a92_t5 )
		| ( { 9{ rl_a92_t4_c1 } } & rl_a92_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_34 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h01 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h02 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h03 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h04 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h05 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h06 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h07 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h08 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h09 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h0a :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h0b :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h0c :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h0d :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h0e :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h0f :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h10 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h11 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h12 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h13 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h14 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h15 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h16 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h17 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h18 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h19 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h1a :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h1b :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h1c :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h1d :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h1e :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h1f :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h20 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h21 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h22 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h23 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h24 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h25 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h26 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h27 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h28 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h29 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h2a :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h2b :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h2c :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h2d :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h2e :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h2f :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h30 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h31 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h32 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h33 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h34 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h35 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h36 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h37 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h38 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h39 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h3a :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h3b :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h3c :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h3d :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h3e :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h3f :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h40 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h41 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h42 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h43 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h44 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h45 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h46 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h47 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h48 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h49 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h4a :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h4b :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h4c :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h4d :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h4e :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h4f :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h50 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h51 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h52 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h53 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h54 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h55 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h56 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h57 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h58 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h59 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h5a :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h5b :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h5c :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h5d :
		rl_a93_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h5e :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h5f :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h60 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h61 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h62 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h63 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h64 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h65 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h66 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h67 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h68 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h69 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h6a :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h6b :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h6c :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h6d :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h6e :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h6f :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h70 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h71 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h72 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h73 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h74 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h75 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h76 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h77 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h78 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h79 :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h7a :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h7b :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h7c :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h7d :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h7e :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	7'h7f :
		rl_a93_t4_t1 = RG_quantized_block_rl_34 ;
	default :
		rl_a93_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a93_t4_t1 or rl_a93_t5 or FF_i )
	begin
	rl_a93_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a93_t4 = ( ( { 9{ FF_i } } & rl_a93_t5 )
		| ( { 9{ rl_a93_t4_c1 } } & rl_a93_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_35 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h01 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h02 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h03 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h04 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h05 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h06 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h07 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h08 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h09 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h0a :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h0b :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h0c :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h0d :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h0e :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h0f :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h10 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h11 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h12 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h13 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h14 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h15 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h16 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h17 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h18 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h19 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h1a :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h1b :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h1c :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h1d :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h1e :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h1f :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h20 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h21 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h22 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h23 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h24 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h25 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h26 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h27 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h28 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h29 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h2a :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h2b :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h2c :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h2d :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h2e :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h2f :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h30 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h31 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h32 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h33 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h34 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h35 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h36 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h37 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h38 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h39 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h3a :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h3b :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h3c :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h3d :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h3e :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h3f :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h40 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h41 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h42 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h43 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h44 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h45 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h46 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h47 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h48 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h49 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h4a :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h4b :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h4c :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h4d :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h4e :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h4f :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h50 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h51 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h52 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h53 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h54 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h55 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h56 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h57 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h58 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h59 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h5a :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h5b :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h5c :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h5d :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h5e :
		rl_a94_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h5f :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h60 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h61 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h62 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h63 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h64 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h65 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h66 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h67 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h68 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h69 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h6a :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h6b :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h6c :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h6d :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h6e :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h6f :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h70 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h71 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h72 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h73 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h74 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h75 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h76 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h77 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h78 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h79 :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h7a :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h7b :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h7c :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h7d :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h7e :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	7'h7f :
		rl_a94_t4_t1 = RG_quantized_block_rl_35 ;
	default :
		rl_a94_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a94_t4_t1 or rl_a94_t5 or FF_i )
	begin
	rl_a94_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a94_t4 = ( ( { 9{ FF_i } } & rl_a94_t5 )
		| ( { 9{ rl_a94_t4_c1 } } & rl_a94_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_36 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h01 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h02 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h03 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h04 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h05 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h06 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h07 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h08 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h09 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h0a :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h0b :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h0c :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h0d :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h0e :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h0f :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h10 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h11 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h12 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h13 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h14 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h15 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h16 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h17 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h18 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h19 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h1a :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h1b :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h1c :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h1d :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h1e :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h1f :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h20 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h21 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h22 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h23 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h24 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h25 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h26 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h27 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h28 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h29 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h2a :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h2b :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h2c :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h2d :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h2e :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h2f :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h30 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h31 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h32 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h33 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h34 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h35 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h36 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h37 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h38 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h39 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h3a :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h3b :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h3c :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h3d :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h3e :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h3f :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h40 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h41 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h42 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h43 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h44 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h45 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h46 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h47 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h48 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h49 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h4a :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h4b :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h4c :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h4d :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h4e :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h4f :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h50 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h51 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h52 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h53 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h54 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h55 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h56 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h57 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h58 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h59 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h5a :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h5b :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h5c :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h5d :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h5e :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h5f :
		rl_a95_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h60 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h61 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h62 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h63 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h64 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h65 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h66 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h67 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h68 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h69 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h6a :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h6b :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h6c :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h6d :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h6e :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h6f :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h70 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h71 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h72 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h73 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h74 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h75 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h76 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h77 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h78 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h79 :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h7a :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h7b :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h7c :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h7d :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h7e :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	7'h7f :
		rl_a95_t4_t1 = RG_quantized_block_rl_36 ;
	default :
		rl_a95_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a95_t4_t1 or rl_a95_t5 or FF_i )
	begin
	rl_a95_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a95_t4 = ( ( { 9{ FF_i } } & rl_a95_t5 )
		| ( { 9{ rl_a95_t4_c1 } } & rl_a95_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_37 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h01 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h02 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h03 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h04 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h05 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h06 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h07 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h08 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h09 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h0a :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h0b :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h0c :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h0d :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h0e :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h0f :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h10 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h11 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h12 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h13 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h14 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h15 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h16 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h17 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h18 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h19 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h1a :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h1b :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h1c :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h1d :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h1e :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h1f :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h20 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h21 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h22 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h23 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h24 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h25 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h26 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h27 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h28 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h29 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h2a :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h2b :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h2c :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h2d :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h2e :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h2f :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h30 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h31 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h32 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h33 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h34 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h35 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h36 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h37 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h38 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h39 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h3a :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h3b :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h3c :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h3d :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h3e :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h3f :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h40 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h41 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h42 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h43 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h44 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h45 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h46 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h47 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h48 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h49 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h4a :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h4b :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h4c :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h4d :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h4e :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h4f :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h50 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h51 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h52 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h53 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h54 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h55 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h56 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h57 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h58 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h59 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h5a :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h5b :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h5c :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h5d :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h5e :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h5f :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h60 :
		rl_a96_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h61 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h62 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h63 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h64 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h65 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h66 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h67 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h68 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h69 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h6a :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h6b :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h6c :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h6d :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h6e :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h6f :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h70 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h71 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h72 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h73 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h74 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h75 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h76 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h77 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h78 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h79 :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h7a :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h7b :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h7c :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h7d :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h7e :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	7'h7f :
		rl_a96_t4_t1 = RG_quantized_block_rl_37 ;
	default :
		rl_a96_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a96_t4_t1 or rl_a96_t5 or FF_i )
	begin
	rl_a96_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a96_t4 = ( ( { 9{ FF_i } } & rl_a96_t5 )
		| ( { 9{ rl_a96_t4_c1 } } & rl_a96_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_38 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h01 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h02 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h03 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h04 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h05 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h06 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h07 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h08 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h09 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h0a :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h0b :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h0c :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h0d :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h0e :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h0f :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h10 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h11 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h12 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h13 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h14 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h15 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h16 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h17 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h18 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h19 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h1a :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h1b :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h1c :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h1d :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h1e :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h1f :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h20 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h21 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h22 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h23 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h24 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h25 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h26 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h27 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h28 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h29 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h2a :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h2b :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h2c :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h2d :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h2e :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h2f :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h30 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h31 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h32 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h33 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h34 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h35 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h36 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h37 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h38 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h39 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h3a :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h3b :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h3c :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h3d :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h3e :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h3f :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h40 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h41 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h42 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h43 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h44 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h45 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h46 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h47 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h48 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h49 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h4a :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h4b :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h4c :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h4d :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h4e :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h4f :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h50 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h51 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h52 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h53 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h54 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h55 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h56 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h57 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h58 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h59 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h5a :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h5b :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h5c :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h5d :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h5e :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h5f :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h60 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h61 :
		rl_a97_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h62 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h63 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h64 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h65 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h66 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h67 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h68 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h69 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h6a :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h6b :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h6c :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h6d :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h6e :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h6f :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h70 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h71 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h72 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h73 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h74 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h75 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h76 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h77 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h78 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h79 :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h7a :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h7b :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h7c :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h7d :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h7e :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	7'h7f :
		rl_a97_t4_t1 = RG_quantized_block_rl_38 ;
	default :
		rl_a97_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a97_t4_t1 or rl_a97_t5 or FF_i )
	begin
	rl_a97_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a97_t4 = ( ( { 9{ FF_i } } & rl_a97_t5 )
		| ( { 9{ rl_a97_t4_c1 } } & rl_a97_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_39 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h01 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h02 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h03 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h04 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h05 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h06 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h07 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h08 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h09 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h0a :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h0b :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h0c :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h0d :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h0e :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h0f :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h10 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h11 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h12 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h13 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h14 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h15 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h16 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h17 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h18 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h19 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h1a :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h1b :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h1c :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h1d :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h1e :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h1f :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h20 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h21 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h22 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h23 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h24 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h25 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h26 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h27 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h28 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h29 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h2a :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h2b :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h2c :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h2d :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h2e :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h2f :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h30 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h31 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h32 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h33 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h34 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h35 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h36 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h37 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h38 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h39 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h3a :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h3b :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h3c :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h3d :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h3e :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h3f :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h40 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h41 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h42 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h43 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h44 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h45 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h46 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h47 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h48 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h49 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h4a :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h4b :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h4c :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h4d :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h4e :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h4f :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h50 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h51 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h52 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h53 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h54 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h55 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h56 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h57 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h58 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h59 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h5a :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h5b :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h5c :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h5d :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h5e :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h5f :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h60 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h61 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h62 :
		rl_a98_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h63 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h64 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h65 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h66 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h67 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h68 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h69 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h6a :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h6b :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h6c :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h6d :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h6e :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h6f :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h70 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h71 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h72 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h73 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h74 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h75 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h76 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h77 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h78 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h79 :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h7a :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h7b :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h7c :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h7d :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h7e :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	7'h7f :
		rl_a98_t4_t1 = RG_quantized_block_rl_39 ;
	default :
		rl_a98_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a98_t4_t1 or rl_a98_t5 or FF_i )
	begin
	rl_a98_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a98_t4 = ( ( { 9{ FF_i } } & rl_a98_t5 )
		| ( { 9{ rl_a98_t4_c1 } } & rl_a98_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_40 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h01 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h02 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h03 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h04 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h05 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h06 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h07 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h08 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h09 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h0a :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h0b :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h0c :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h0d :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h0e :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h0f :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h10 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h11 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h12 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h13 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h14 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h15 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h16 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h17 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h18 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h19 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h1a :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h1b :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h1c :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h1d :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h1e :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h1f :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h20 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h21 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h22 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h23 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h24 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h25 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h26 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h27 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h28 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h29 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h2a :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h2b :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h2c :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h2d :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h2e :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h2f :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h30 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h31 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h32 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h33 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h34 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h35 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h36 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h37 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h38 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h39 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h3a :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h3b :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h3c :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h3d :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h3e :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h3f :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h40 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h41 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h42 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h43 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h44 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h45 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h46 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h47 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h48 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h49 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h4a :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h4b :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h4c :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h4d :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h4e :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h4f :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h50 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h51 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h52 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h53 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h54 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h55 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h56 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h57 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h58 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h59 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h5a :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h5b :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h5c :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h5d :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h5e :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h5f :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h60 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h61 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h62 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h63 :
		rl_a99_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h64 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h65 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h66 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h67 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h68 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h69 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h6a :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h6b :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h6c :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h6d :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h6e :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h6f :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h70 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h71 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h72 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h73 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h74 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h75 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h76 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h77 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h78 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h79 :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h7a :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h7b :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h7c :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h7d :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h7e :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	7'h7f :
		rl_a99_t4_t1 = RG_quantized_block_rl_40 ;
	default :
		rl_a99_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a99_t4_t1 or rl_a99_t5 or FF_i )
	begin
	rl_a99_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a99_t4 = ( ( { 9{ FF_i } } & rl_a99_t5 )
		| ( { 9{ rl_a99_t4_c1 } } & rl_a99_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_41 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h01 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h02 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h03 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h04 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h05 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h06 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h07 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h08 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h09 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h0a :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h0b :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h0c :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h0d :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h0e :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h0f :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h10 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h11 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h12 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h13 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h14 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h15 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h16 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h17 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h18 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h19 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h1a :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h1b :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h1c :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h1d :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h1e :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h1f :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h20 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h21 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h22 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h23 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h24 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h25 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h26 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h27 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h28 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h29 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h2a :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h2b :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h2c :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h2d :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h2e :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h2f :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h30 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h31 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h32 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h33 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h34 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h35 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h36 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h37 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h38 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h39 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h3a :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h3b :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h3c :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h3d :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h3e :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h3f :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h40 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h41 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h42 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h43 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h44 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h45 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h46 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h47 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h48 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h49 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h4a :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h4b :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h4c :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h4d :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h4e :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h4f :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h50 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h51 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h52 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h53 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h54 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h55 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h56 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h57 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h58 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h59 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h5a :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h5b :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h5c :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h5d :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h5e :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h5f :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h60 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h61 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h62 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h63 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h64 :
		rl_a100_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h65 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h66 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h67 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h68 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h69 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h6a :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h6b :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h6c :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h6d :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h6e :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h6f :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h70 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h71 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h72 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h73 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h74 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h75 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h76 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h77 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h78 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h79 :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h7a :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h7b :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h7c :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h7d :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h7e :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	7'h7f :
		rl_a100_t4_t1 = RG_quantized_block_rl_41 ;
	default :
		rl_a100_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a100_t4_t1 or rl_a100_t5 or FF_i )
	begin
	rl_a100_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a100_t4 = ( ( { 9{ FF_i } } & rl_a100_t5 )
		| ( { 9{ rl_a100_t4_c1 } } & rl_a100_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_42 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h01 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h02 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h03 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h04 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h05 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h06 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h07 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h08 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h09 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h0a :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h0b :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h0c :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h0d :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h0e :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h0f :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h10 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h11 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h12 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h13 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h14 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h15 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h16 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h17 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h18 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h19 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h1a :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h1b :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h1c :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h1d :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h1e :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h1f :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h20 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h21 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h22 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h23 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h24 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h25 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h26 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h27 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h28 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h29 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h2a :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h2b :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h2c :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h2d :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h2e :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h2f :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h30 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h31 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h32 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h33 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h34 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h35 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h36 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h37 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h38 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h39 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h3a :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h3b :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h3c :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h3d :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h3e :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h3f :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h40 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h41 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h42 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h43 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h44 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h45 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h46 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h47 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h48 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h49 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h4a :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h4b :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h4c :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h4d :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h4e :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h4f :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h50 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h51 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h52 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h53 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h54 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h55 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h56 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h57 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h58 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h59 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h5a :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h5b :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h5c :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h5d :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h5e :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h5f :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h60 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h61 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h62 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h63 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h64 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h65 :
		rl_a101_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h66 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h67 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h68 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h69 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h6a :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h6b :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h6c :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h6d :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h6e :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h6f :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h70 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h71 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h72 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h73 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h74 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h75 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h76 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h77 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h78 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h79 :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h7a :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h7b :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h7c :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h7d :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h7e :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	7'h7f :
		rl_a101_t4_t1 = RG_quantized_block_rl_42 ;
	default :
		rl_a101_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a101_t4_t1 or rl_a101_t5 or FF_i )
	begin
	rl_a101_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a101_t4 = ( ( { 9{ FF_i } } & rl_a101_t5 )
		| ( { 9{ rl_a101_t4_c1 } } & rl_a101_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_43 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h01 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h02 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h03 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h04 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h05 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h06 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h07 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h08 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h09 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h0a :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h0b :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h0c :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h0d :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h0e :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h0f :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h10 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h11 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h12 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h13 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h14 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h15 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h16 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h17 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h18 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h19 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h1a :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h1b :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h1c :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h1d :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h1e :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h1f :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h20 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h21 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h22 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h23 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h24 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h25 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h26 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h27 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h28 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h29 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h2a :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h2b :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h2c :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h2d :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h2e :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h2f :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h30 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h31 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h32 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h33 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h34 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h35 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h36 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h37 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h38 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h39 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h3a :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h3b :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h3c :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h3d :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h3e :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h3f :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h40 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h41 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h42 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h43 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h44 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h45 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h46 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h47 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h48 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h49 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h4a :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h4b :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h4c :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h4d :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h4e :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h4f :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h50 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h51 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h52 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h53 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h54 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h55 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h56 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h57 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h58 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h59 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h5a :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h5b :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h5c :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h5d :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h5e :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h5f :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h60 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h61 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h62 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h63 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h64 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h65 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h66 :
		rl_a102_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h67 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h68 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h69 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h6a :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h6b :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h6c :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h6d :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h6e :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h6f :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h70 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h71 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h72 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h73 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h74 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h75 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h76 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h77 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h78 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h79 :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h7a :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h7b :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h7c :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h7d :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h7e :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	7'h7f :
		rl_a102_t4_t1 = RG_quantized_block_rl_43 ;
	default :
		rl_a102_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a102_t4_t1 or rl_a102_t5 or FF_i )
	begin
	rl_a102_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a102_t4 = ( ( { 9{ FF_i } } & rl_a102_t5 )
		| ( { 9{ rl_a102_t4_c1 } } & rl_a102_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_44 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h01 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h02 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h03 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h04 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h05 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h06 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h07 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h08 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h09 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h0a :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h0b :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h0c :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h0d :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h0e :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h0f :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h10 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h11 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h12 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h13 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h14 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h15 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h16 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h17 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h18 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h19 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h1a :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h1b :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h1c :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h1d :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h1e :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h1f :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h20 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h21 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h22 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h23 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h24 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h25 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h26 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h27 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h28 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h29 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h2a :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h2b :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h2c :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h2d :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h2e :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h2f :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h30 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h31 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h32 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h33 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h34 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h35 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h36 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h37 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h38 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h39 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h3a :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h3b :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h3c :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h3d :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h3e :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h3f :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h40 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h41 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h42 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h43 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h44 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h45 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h46 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h47 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h48 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h49 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h4a :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h4b :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h4c :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h4d :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h4e :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h4f :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h50 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h51 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h52 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h53 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h54 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h55 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h56 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h57 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h58 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h59 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h5a :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h5b :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h5c :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h5d :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h5e :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h5f :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h60 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h61 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h62 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h63 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h64 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h65 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h66 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h67 :
		rl_a103_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h68 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h69 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h6a :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h6b :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h6c :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h6d :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h6e :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h6f :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h70 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h71 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h72 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h73 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h74 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h75 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h76 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h77 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h78 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h79 :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h7a :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h7b :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h7c :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h7d :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h7e :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	7'h7f :
		rl_a103_t4_t1 = RG_quantized_block_rl_44 ;
	default :
		rl_a103_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a103_t4_t1 or rl_a103_t5 or FF_i )
	begin
	rl_a103_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a103_t4 = ( ( { 9{ FF_i } } & rl_a103_t5 )
		| ( { 9{ rl_a103_t4_c1 } } & rl_a103_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_45 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h01 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h02 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h03 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h04 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h05 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h06 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h07 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h08 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h09 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h0a :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h0b :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h0c :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h0d :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h0e :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h0f :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h10 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h11 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h12 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h13 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h14 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h15 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h16 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h17 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h18 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h19 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h1a :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h1b :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h1c :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h1d :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h1e :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h1f :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h20 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h21 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h22 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h23 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h24 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h25 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h26 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h27 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h28 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h29 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h2a :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h2b :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h2c :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h2d :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h2e :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h2f :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h30 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h31 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h32 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h33 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h34 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h35 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h36 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h37 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h38 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h39 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h3a :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h3b :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h3c :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h3d :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h3e :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h3f :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h40 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h41 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h42 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h43 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h44 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h45 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h46 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h47 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h48 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h49 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h4a :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h4b :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h4c :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h4d :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h4e :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h4f :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h50 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h51 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h52 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h53 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h54 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h55 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h56 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h57 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h58 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h59 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h5a :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h5b :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h5c :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h5d :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h5e :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h5f :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h60 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h61 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h62 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h63 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h64 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h65 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h66 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h67 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h68 :
		rl_a104_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h69 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h6a :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h6b :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h6c :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h6d :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h6e :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h6f :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h70 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h71 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h72 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h73 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h74 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h75 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h76 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h77 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h78 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h79 :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h7a :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h7b :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h7c :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h7d :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h7e :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	7'h7f :
		rl_a104_t4_t1 = RG_quantized_block_rl_45 ;
	default :
		rl_a104_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a104_t4_t1 or rl_a104_t5 or FF_i )
	begin
	rl_a104_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a104_t4 = ( ( { 9{ FF_i } } & rl_a104_t5 )
		| ( { 9{ rl_a104_t4_c1 } } & rl_a104_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_46 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h01 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h02 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h03 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h04 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h05 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h06 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h07 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h08 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h09 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h0a :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h0b :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h0c :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h0d :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h0e :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h0f :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h10 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h11 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h12 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h13 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h14 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h15 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h16 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h17 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h18 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h19 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h1a :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h1b :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h1c :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h1d :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h1e :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h1f :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h20 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h21 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h22 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h23 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h24 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h25 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h26 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h27 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h28 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h29 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h2a :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h2b :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h2c :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h2d :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h2e :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h2f :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h30 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h31 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h32 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h33 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h34 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h35 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h36 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h37 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h38 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h39 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h3a :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h3b :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h3c :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h3d :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h3e :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h3f :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h40 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h41 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h42 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h43 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h44 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h45 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h46 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h47 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h48 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h49 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h4a :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h4b :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h4c :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h4d :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h4e :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h4f :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h50 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h51 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h52 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h53 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h54 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h55 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h56 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h57 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h58 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h59 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h5a :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h5b :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h5c :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h5d :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h5e :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h5f :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h60 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h61 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h62 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h63 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h64 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h65 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h66 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h67 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h68 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h69 :
		rl_a105_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h6a :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h6b :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h6c :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h6d :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h6e :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h6f :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h70 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h71 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h72 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h73 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h74 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h75 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h76 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h77 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h78 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h79 :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h7a :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h7b :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h7c :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h7d :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h7e :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	7'h7f :
		rl_a105_t4_t1 = RG_quantized_block_rl_46 ;
	default :
		rl_a105_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a105_t4_t1 or rl_a105_t5 or FF_i )
	begin
	rl_a105_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a105_t4 = ( ( { 9{ FF_i } } & rl_a105_t5 )
		| ( { 9{ rl_a105_t4_c1 } } & rl_a105_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_47 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h01 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h02 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h03 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h04 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h05 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h06 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h07 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h08 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h09 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h0a :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h0b :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h0c :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h0d :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h0e :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h0f :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h10 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h11 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h12 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h13 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h14 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h15 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h16 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h17 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h18 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h19 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h1a :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h1b :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h1c :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h1d :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h1e :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h1f :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h20 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h21 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h22 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h23 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h24 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h25 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h26 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h27 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h28 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h29 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h2a :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h2b :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h2c :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h2d :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h2e :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h2f :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h30 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h31 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h32 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h33 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h34 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h35 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h36 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h37 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h38 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h39 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h3a :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h3b :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h3c :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h3d :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h3e :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h3f :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h40 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h41 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h42 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h43 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h44 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h45 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h46 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h47 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h48 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h49 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h4a :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h4b :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h4c :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h4d :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h4e :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h4f :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h50 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h51 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h52 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h53 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h54 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h55 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h56 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h57 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h58 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h59 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h5a :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h5b :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h5c :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h5d :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h5e :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h5f :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h60 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h61 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h62 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h63 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h64 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h65 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h66 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h67 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h68 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h69 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h6a :
		rl_a106_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h6b :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h6c :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h6d :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h6e :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h6f :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h70 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h71 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h72 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h73 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h74 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h75 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h76 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h77 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h78 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h79 :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h7a :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h7b :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h7c :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h7d :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h7e :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	7'h7f :
		rl_a106_t4_t1 = RG_quantized_block_rl_47 ;
	default :
		rl_a106_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a106_t4_t1 or rl_a106_t5 or FF_i )
	begin
	rl_a106_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a106_t4 = ( ( { 9{ FF_i } } & rl_a106_t5 )
		| ( { 9{ rl_a106_t4_c1 } } & rl_a106_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_48 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h01 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h02 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h03 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h04 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h05 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h06 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h07 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h08 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h09 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h0a :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h0b :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h0c :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h0d :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h0e :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h0f :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h10 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h11 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h12 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h13 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h14 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h15 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h16 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h17 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h18 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h19 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h1a :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h1b :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h1c :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h1d :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h1e :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h1f :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h20 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h21 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h22 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h23 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h24 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h25 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h26 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h27 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h28 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h29 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h2a :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h2b :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h2c :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h2d :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h2e :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h2f :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h30 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h31 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h32 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h33 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h34 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h35 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h36 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h37 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h38 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h39 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h3a :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h3b :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h3c :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h3d :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h3e :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h3f :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h40 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h41 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h42 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h43 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h44 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h45 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h46 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h47 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h48 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h49 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h4a :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h4b :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h4c :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h4d :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h4e :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h4f :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h50 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h51 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h52 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h53 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h54 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h55 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h56 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h57 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h58 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h59 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h5a :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h5b :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h5c :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h5d :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h5e :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h5f :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h60 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h61 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h62 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h63 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h64 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h65 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h66 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h67 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h68 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h69 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h6a :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h6b :
		rl_a107_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h6c :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h6d :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h6e :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h6f :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h70 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h71 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h72 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h73 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h74 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h75 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h76 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h77 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h78 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h79 :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h7a :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h7b :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h7c :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h7d :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h7e :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	7'h7f :
		rl_a107_t4_t1 = RG_quantized_block_rl_48 ;
	default :
		rl_a107_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a107_t4_t1 or rl_a107_t5 or FF_i )
	begin
	rl_a107_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a107_t4 = ( ( { 9{ FF_i } } & rl_a107_t5 )
		| ( { 9{ rl_a107_t4_c1 } } & rl_a107_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_49 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h01 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h02 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h03 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h04 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h05 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h06 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h07 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h08 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h09 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h0a :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h0b :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h0c :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h0d :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h0e :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h0f :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h10 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h11 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h12 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h13 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h14 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h15 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h16 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h17 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h18 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h19 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h1a :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h1b :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h1c :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h1d :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h1e :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h1f :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h20 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h21 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h22 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h23 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h24 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h25 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h26 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h27 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h28 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h29 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h2a :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h2b :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h2c :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h2d :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h2e :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h2f :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h30 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h31 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h32 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h33 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h34 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h35 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h36 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h37 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h38 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h39 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h3a :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h3b :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h3c :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h3d :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h3e :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h3f :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h40 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h41 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h42 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h43 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h44 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h45 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h46 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h47 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h48 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h49 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h4a :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h4b :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h4c :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h4d :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h4e :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h4f :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h50 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h51 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h52 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h53 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h54 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h55 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h56 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h57 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h58 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h59 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h5a :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h5b :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h5c :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h5d :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h5e :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h5f :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h60 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h61 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h62 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h63 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h64 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h65 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h66 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h67 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h68 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h69 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h6a :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h6b :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h6c :
		rl_a108_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h6d :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h6e :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h6f :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h70 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h71 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h72 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h73 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h74 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h75 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h76 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h77 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h78 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h79 :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h7a :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h7b :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h7c :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h7d :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h7e :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	7'h7f :
		rl_a108_t4_t1 = RG_quantized_block_rl_49 ;
	default :
		rl_a108_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a108_t4_t1 or rl_a108_t5 or FF_i )
	begin
	rl_a108_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a108_t4 = ( ( { 9{ FF_i } } & rl_a108_t5 )
		| ( { 9{ rl_a108_t4_c1 } } & rl_a108_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_50 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h01 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h02 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h03 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h04 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h05 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h06 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h07 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h08 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h09 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h0a :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h0b :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h0c :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h0d :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h0e :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h0f :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h10 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h11 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h12 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h13 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h14 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h15 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h16 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h17 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h18 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h19 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h1a :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h1b :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h1c :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h1d :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h1e :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h1f :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h20 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h21 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h22 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h23 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h24 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h25 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h26 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h27 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h28 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h29 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h2a :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h2b :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h2c :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h2d :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h2e :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h2f :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h30 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h31 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h32 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h33 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h34 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h35 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h36 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h37 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h38 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h39 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h3a :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h3b :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h3c :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h3d :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h3e :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h3f :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h40 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h41 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h42 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h43 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h44 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h45 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h46 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h47 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h48 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h49 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h4a :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h4b :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h4c :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h4d :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h4e :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h4f :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h50 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h51 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h52 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h53 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h54 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h55 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h56 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h57 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h58 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h59 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h5a :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h5b :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h5c :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h5d :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h5e :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h5f :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h60 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h61 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h62 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h63 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h64 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h65 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h66 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h67 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h68 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h69 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h6a :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h6b :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h6c :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h6d :
		rl_a109_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h6e :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h6f :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h70 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h71 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h72 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h73 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h74 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h75 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h76 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h77 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h78 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h79 :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h7a :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h7b :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h7c :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h7d :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h7e :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	7'h7f :
		rl_a109_t4_t1 = RG_quantized_block_rl_50 ;
	default :
		rl_a109_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a109_t4_t1 or rl_a109_t5 or FF_i )
	begin
	rl_a109_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a109_t4 = ( ( { 9{ FF_i } } & rl_a109_t5 )
		| ( { 9{ rl_a109_t4_c1 } } & rl_a109_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_51 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h01 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h02 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h03 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h04 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h05 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h06 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h07 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h08 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h09 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h0a :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h0b :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h0c :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h0d :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h0e :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h0f :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h10 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h11 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h12 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h13 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h14 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h15 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h16 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h17 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h18 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h19 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h1a :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h1b :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h1c :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h1d :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h1e :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h1f :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h20 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h21 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h22 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h23 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h24 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h25 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h26 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h27 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h28 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h29 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h2a :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h2b :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h2c :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h2d :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h2e :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h2f :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h30 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h31 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h32 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h33 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h34 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h35 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h36 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h37 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h38 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h39 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h3a :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h3b :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h3c :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h3d :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h3e :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h3f :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h40 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h41 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h42 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h43 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h44 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h45 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h46 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h47 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h48 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h49 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h4a :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h4b :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h4c :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h4d :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h4e :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h4f :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h50 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h51 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h52 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h53 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h54 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h55 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h56 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h57 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h58 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h59 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h5a :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h5b :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h5c :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h5d :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h5e :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h5f :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h60 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h61 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h62 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h63 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h64 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h65 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h66 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h67 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h68 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h69 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h6a :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h6b :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h6c :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h6d :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h6e :
		rl_a110_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h6f :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h70 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h71 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h72 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h73 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h74 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h75 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h76 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h77 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h78 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h79 :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h7a :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h7b :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h7c :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h7d :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h7e :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	7'h7f :
		rl_a110_t4_t1 = RG_quantized_block_rl_51 ;
	default :
		rl_a110_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a110_t4_t1 or rl_a110_t5 or FF_i )
	begin
	rl_a110_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a110_t4 = ( ( { 9{ FF_i } } & rl_a110_t5 )
		| ( { 9{ rl_a110_t4_c1 } } & rl_a110_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_52 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h01 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h02 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h03 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h04 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h05 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h06 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h07 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h08 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h09 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h0a :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h0b :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h0c :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h0d :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h0e :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h0f :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h10 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h11 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h12 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h13 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h14 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h15 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h16 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h17 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h18 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h19 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h1a :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h1b :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h1c :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h1d :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h1e :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h1f :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h20 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h21 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h22 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h23 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h24 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h25 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h26 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h27 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h28 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h29 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h2a :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h2b :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h2c :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h2d :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h2e :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h2f :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h30 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h31 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h32 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h33 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h34 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h35 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h36 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h37 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h38 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h39 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h3a :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h3b :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h3c :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h3d :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h3e :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h3f :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h40 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h41 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h42 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h43 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h44 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h45 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h46 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h47 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h48 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h49 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h4a :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h4b :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h4c :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h4d :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h4e :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h4f :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h50 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h51 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h52 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h53 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h54 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h55 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h56 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h57 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h58 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h59 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h5a :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h5b :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h5c :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h5d :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h5e :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h5f :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h60 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h61 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h62 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h63 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h64 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h65 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h66 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h67 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h68 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h69 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h6a :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h6b :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h6c :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h6d :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h6e :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h6f :
		rl_a111_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h70 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h71 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h72 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h73 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h74 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h75 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h76 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h77 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h78 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h79 :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h7a :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h7b :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h7c :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h7d :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h7e :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	7'h7f :
		rl_a111_t4_t1 = RG_quantized_block_rl_52 ;
	default :
		rl_a111_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a111_t4_t1 or rl_a111_t5 or FF_i )
	begin
	rl_a111_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a111_t4 = ( ( { 9{ FF_i } } & rl_a111_t5 )
		| ( { 9{ rl_a111_t4_c1 } } & rl_a111_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_53 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h01 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h02 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h03 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h04 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h05 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h06 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h07 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h08 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h09 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h0a :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h0b :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h0c :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h0d :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h0e :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h0f :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h10 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h11 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h12 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h13 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h14 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h15 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h16 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h17 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h18 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h19 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h1a :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h1b :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h1c :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h1d :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h1e :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h1f :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h20 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h21 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h22 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h23 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h24 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h25 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h26 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h27 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h28 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h29 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h2a :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h2b :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h2c :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h2d :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h2e :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h2f :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h30 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h31 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h32 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h33 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h34 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h35 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h36 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h37 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h38 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h39 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h3a :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h3b :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h3c :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h3d :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h3e :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h3f :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h40 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h41 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h42 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h43 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h44 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h45 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h46 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h47 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h48 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h49 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h4a :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h4b :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h4c :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h4d :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h4e :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h4f :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h50 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h51 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h52 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h53 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h54 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h55 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h56 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h57 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h58 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h59 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h5a :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h5b :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h5c :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h5d :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h5e :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h5f :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h60 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h61 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h62 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h63 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h64 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h65 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h66 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h67 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h68 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h69 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h6a :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h6b :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h6c :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h6d :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h6e :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h6f :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h70 :
		rl_a112_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h71 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h72 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h73 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h74 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h75 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h76 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h77 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h78 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h79 :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h7a :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h7b :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h7c :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h7d :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h7e :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	7'h7f :
		rl_a112_t4_t1 = RG_quantized_block_rl_53 ;
	default :
		rl_a112_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a112_t4_t1 or rl_a112_t5 or FF_i )
	begin
	rl_a112_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a112_t4 = ( ( { 9{ FF_i } } & rl_a112_t5 )
		| ( { 9{ rl_a112_t4_c1 } } & rl_a112_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_54 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h01 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h02 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h03 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h04 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h05 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h06 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h07 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h08 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h09 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h0a :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h0b :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h0c :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h0d :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h0e :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h0f :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h10 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h11 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h12 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h13 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h14 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h15 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h16 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h17 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h18 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h19 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h1a :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h1b :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h1c :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h1d :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h1e :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h1f :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h20 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h21 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h22 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h23 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h24 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h25 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h26 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h27 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h28 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h29 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h2a :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h2b :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h2c :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h2d :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h2e :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h2f :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h30 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h31 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h32 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h33 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h34 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h35 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h36 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h37 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h38 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h39 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h3a :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h3b :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h3c :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h3d :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h3e :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h3f :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h40 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h41 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h42 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h43 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h44 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h45 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h46 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h47 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h48 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h49 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h4a :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h4b :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h4c :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h4d :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h4e :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h4f :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h50 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h51 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h52 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h53 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h54 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h55 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h56 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h57 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h58 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h59 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h5a :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h5b :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h5c :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h5d :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h5e :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h5f :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h60 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h61 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h62 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h63 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h64 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h65 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h66 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h67 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h68 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h69 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h6a :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h6b :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h6c :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h6d :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h6e :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h6f :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h70 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h71 :
		rl_a113_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h72 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h73 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h74 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h75 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h76 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h77 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h78 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h79 :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h7a :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h7b :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h7c :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h7d :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h7e :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	7'h7f :
		rl_a113_t4_t1 = RG_quantized_block_rl_54 ;
	default :
		rl_a113_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a113_t4_t1 or rl_a113_t5 or FF_i )
	begin
	rl_a113_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a113_t4 = ( ( { 9{ FF_i } } & rl_a113_t5 )
		| ( { 9{ rl_a113_t4_c1 } } & rl_a113_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_55 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h01 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h02 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h03 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h04 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h05 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h06 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h07 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h08 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h09 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h0a :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h0b :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h0c :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h0d :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h0e :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h0f :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h10 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h11 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h12 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h13 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h14 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h15 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h16 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h17 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h18 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h19 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h1a :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h1b :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h1c :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h1d :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h1e :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h1f :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h20 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h21 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h22 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h23 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h24 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h25 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h26 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h27 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h28 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h29 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h2a :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h2b :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h2c :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h2d :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h2e :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h2f :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h30 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h31 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h32 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h33 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h34 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h35 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h36 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h37 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h38 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h39 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h3a :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h3b :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h3c :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h3d :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h3e :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h3f :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h40 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h41 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h42 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h43 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h44 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h45 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h46 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h47 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h48 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h49 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h4a :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h4b :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h4c :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h4d :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h4e :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h4f :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h50 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h51 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h52 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h53 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h54 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h55 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h56 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h57 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h58 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h59 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h5a :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h5b :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h5c :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h5d :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h5e :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h5f :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h60 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h61 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h62 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h63 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h64 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h65 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h66 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h67 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h68 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h69 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h6a :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h6b :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h6c :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h6d :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h6e :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h6f :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h70 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h71 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h72 :
		rl_a114_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h73 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h74 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h75 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h76 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h77 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h78 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h79 :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h7a :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h7b :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h7c :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h7d :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h7e :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	7'h7f :
		rl_a114_t4_t1 = RG_quantized_block_rl_55 ;
	default :
		rl_a114_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a114_t4_t1 or rl_a114_t5 or FF_i )
	begin
	rl_a114_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a114_t4 = ( ( { 9{ FF_i } } & rl_a114_t5 )
		| ( { 9{ rl_a114_t4_c1 } } & rl_a114_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_56 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h01 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h02 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h03 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h04 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h05 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h06 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h07 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h08 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h09 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h0a :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h0b :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h0c :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h0d :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h0e :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h0f :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h10 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h11 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h12 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h13 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h14 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h15 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h16 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h17 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h18 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h19 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h1a :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h1b :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h1c :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h1d :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h1e :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h1f :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h20 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h21 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h22 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h23 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h24 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h25 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h26 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h27 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h28 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h29 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h2a :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h2b :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h2c :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h2d :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h2e :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h2f :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h30 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h31 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h32 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h33 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h34 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h35 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h36 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h37 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h38 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h39 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h3a :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h3b :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h3c :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h3d :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h3e :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h3f :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h40 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h41 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h42 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h43 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h44 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h45 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h46 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h47 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h48 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h49 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h4a :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h4b :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h4c :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h4d :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h4e :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h4f :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h50 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h51 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h52 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h53 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h54 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h55 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h56 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h57 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h58 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h59 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h5a :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h5b :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h5c :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h5d :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h5e :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h5f :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h60 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h61 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h62 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h63 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h64 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h65 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h66 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h67 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h68 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h69 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h6a :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h6b :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h6c :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h6d :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h6e :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h6f :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h70 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h71 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h72 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h73 :
		rl_a115_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h74 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h75 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h76 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h77 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h78 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h79 :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h7a :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h7b :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h7c :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h7d :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h7e :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	7'h7f :
		rl_a115_t4_t1 = RG_quantized_block_rl_56 ;
	default :
		rl_a115_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a115_t4_t1 or rl_a115_t5 or FF_i )
	begin
	rl_a115_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a115_t4 = ( ( { 9{ FF_i } } & rl_a115_t5 )
		| ( { 9{ rl_a115_t4_c1 } } & rl_a115_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_242 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h01 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h02 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h03 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h04 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h05 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h06 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h07 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h08 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h09 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h0a :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h0b :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h0c :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h0d :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h0e :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h0f :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h10 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h11 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h12 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h13 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h14 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h15 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h16 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h17 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h18 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h19 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h1a :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h1b :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h1c :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h1d :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h1e :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h1f :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h20 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h21 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h22 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h23 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h24 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h25 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h26 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h27 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h28 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h29 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h2a :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h2b :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h2c :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h2d :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h2e :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h2f :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h30 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h31 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h32 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h33 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h34 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h35 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h36 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h37 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h38 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h39 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h3a :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h3b :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h3c :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h3d :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h3e :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h3f :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h40 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h41 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h42 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h43 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h44 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h45 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h46 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h47 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h48 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h49 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h4a :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h4b :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h4c :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h4d :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h4e :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h4f :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h50 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h51 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h52 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h53 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h54 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h55 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h56 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h57 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h58 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h59 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h5a :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h5b :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h5c :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h5d :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h5e :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h5f :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h60 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h61 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h62 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h63 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h64 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h65 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h66 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h67 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h68 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h69 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h6a :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h6b :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h6c :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h6d :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h6e :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h6f :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h70 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h71 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h72 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h73 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h74 :
		rl_a116_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h75 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h76 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h77 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h78 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h79 :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h7a :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h7b :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h7c :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h7d :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h7e :
		rl_a116_t4_t1 = RG_rl_242 ;
	7'h7f :
		rl_a116_t4_t1 = RG_rl_242 ;
	default :
		rl_a116_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a116_t4_t1 or rl_a116_t5 or FF_i )
	begin
	rl_a116_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a116_t4 = ( ( { 9{ FF_i } } & rl_a116_t5 )
		| ( { 9{ rl_a116_t4_c1 } } & rl_a116_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_57 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h01 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h02 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h03 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h04 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h05 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h06 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h07 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h08 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h09 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h0a :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h0b :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h0c :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h0d :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h0e :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h0f :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h10 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h11 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h12 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h13 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h14 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h15 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h16 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h17 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h18 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h19 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h1a :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h1b :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h1c :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h1d :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h1e :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h1f :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h20 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h21 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h22 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h23 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h24 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h25 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h26 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h27 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h28 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h29 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h2a :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h2b :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h2c :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h2d :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h2e :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h2f :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h30 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h31 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h32 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h33 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h34 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h35 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h36 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h37 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h38 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h39 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h3a :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h3b :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h3c :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h3d :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h3e :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h3f :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h40 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h41 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h42 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h43 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h44 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h45 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h46 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h47 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h48 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h49 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h4a :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h4b :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h4c :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h4d :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h4e :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h4f :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h50 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h51 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h52 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h53 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h54 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h55 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h56 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h57 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h58 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h59 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h5a :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h5b :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h5c :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h5d :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h5e :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h5f :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h60 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h61 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h62 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h63 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h64 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h65 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h66 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h67 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h68 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h69 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h6a :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h6b :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h6c :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h6d :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h6e :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h6f :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h70 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h71 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h72 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h73 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h74 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h75 :
		rl_a117_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h76 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h77 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h78 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h79 :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h7a :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h7b :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h7c :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h7d :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h7e :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	7'h7f :
		rl_a117_t4_t1 = RG_quantized_block_rl_57 ;
	default :
		rl_a117_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a117_t4_t1 or rl_a117_t5 or FF_i )
	begin
	rl_a117_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a117_t4 = ( ( { 9{ FF_i } } & rl_a117_t5 )
		| ( { 9{ rl_a117_t4_c1 } } & rl_a117_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_243 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h01 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h02 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h03 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h04 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h05 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h06 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h07 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h08 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h09 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h0a :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h0b :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h0c :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h0d :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h0e :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h0f :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h10 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h11 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h12 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h13 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h14 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h15 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h16 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h17 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h18 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h19 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h1a :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h1b :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h1c :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h1d :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h1e :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h1f :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h20 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h21 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h22 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h23 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h24 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h25 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h26 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h27 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h28 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h29 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h2a :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h2b :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h2c :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h2d :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h2e :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h2f :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h30 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h31 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h32 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h33 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h34 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h35 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h36 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h37 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h38 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h39 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h3a :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h3b :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h3c :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h3d :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h3e :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h3f :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h40 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h41 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h42 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h43 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h44 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h45 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h46 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h47 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h48 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h49 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h4a :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h4b :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h4c :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h4d :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h4e :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h4f :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h50 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h51 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h52 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h53 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h54 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h55 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h56 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h57 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h58 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h59 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h5a :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h5b :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h5c :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h5d :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h5e :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h5f :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h60 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h61 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h62 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h63 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h64 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h65 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h66 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h67 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h68 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h69 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h6a :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h6b :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h6c :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h6d :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h6e :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h6f :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h70 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h71 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h72 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h73 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h74 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h75 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h76 :
		rl_a118_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h77 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h78 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h79 :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h7a :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h7b :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h7c :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h7d :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h7e :
		rl_a118_t4_t1 = RG_rl_243 ;
	7'h7f :
		rl_a118_t4_t1 = RG_rl_243 ;
	default :
		rl_a118_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a118_t4_t1 or rl_a118_t5 or FF_i )
	begin
	rl_a118_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a118_t4 = ( ( { 9{ FF_i } } & rl_a118_t5 )
		| ( { 9{ rl_a118_t4_c1 } } & rl_a118_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_58 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h01 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h02 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h03 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h04 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h05 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h06 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h07 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h08 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h09 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h0a :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h0b :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h0c :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h0d :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h0e :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h0f :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h10 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h11 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h12 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h13 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h14 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h15 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h16 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h17 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h18 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h19 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h1a :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h1b :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h1c :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h1d :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h1e :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h1f :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h20 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h21 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h22 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h23 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h24 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h25 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h26 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h27 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h28 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h29 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h2a :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h2b :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h2c :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h2d :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h2e :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h2f :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h30 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h31 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h32 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h33 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h34 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h35 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h36 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h37 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h38 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h39 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h3a :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h3b :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h3c :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h3d :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h3e :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h3f :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h40 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h41 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h42 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h43 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h44 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h45 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h46 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h47 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h48 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h49 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h4a :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h4b :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h4c :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h4d :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h4e :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h4f :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h50 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h51 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h52 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h53 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h54 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h55 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h56 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h57 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h58 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h59 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h5a :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h5b :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h5c :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h5d :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h5e :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h5f :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h60 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h61 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h62 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h63 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h64 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h65 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h66 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h67 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h68 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h69 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h6a :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h6b :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h6c :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h6d :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h6e :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h6f :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h70 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h71 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h72 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h73 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h74 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h75 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h76 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h77 :
		rl_a119_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h78 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h79 :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h7a :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h7b :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h7c :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h7d :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h7e :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	7'h7f :
		rl_a119_t4_t1 = RG_quantized_block_rl_58 ;
	default :
		rl_a119_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a119_t4_t1 or rl_a119_t5 or FF_i )
	begin
	rl_a119_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a119_t4 = ( ( { 9{ FF_i } } & rl_a119_t5 )
		| ( { 9{ rl_a119_t4_c1 } } & rl_a119_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_244 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h01 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h02 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h03 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h04 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h05 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h06 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h07 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h08 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h09 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h0a :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h0b :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h0c :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h0d :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h0e :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h0f :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h10 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h11 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h12 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h13 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h14 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h15 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h16 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h17 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h18 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h19 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h1a :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h1b :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h1c :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h1d :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h1e :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h1f :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h20 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h21 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h22 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h23 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h24 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h25 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h26 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h27 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h28 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h29 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h2a :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h2b :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h2c :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h2d :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h2e :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h2f :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h30 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h31 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h32 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h33 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h34 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h35 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h36 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h37 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h38 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h39 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h3a :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h3b :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h3c :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h3d :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h3e :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h3f :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h40 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h41 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h42 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h43 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h44 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h45 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h46 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h47 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h48 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h49 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h4a :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h4b :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h4c :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h4d :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h4e :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h4f :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h50 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h51 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h52 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h53 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h54 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h55 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h56 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h57 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h58 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h59 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h5a :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h5b :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h5c :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h5d :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h5e :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h5f :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h60 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h61 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h62 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h63 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h64 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h65 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h66 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h67 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h68 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h69 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h6a :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h6b :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h6c :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h6d :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h6e :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h6f :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h70 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h71 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h72 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h73 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h74 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h75 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h76 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h77 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h78 :
		rl_a120_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h79 :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h7a :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h7b :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h7c :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h7d :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h7e :
		rl_a120_t4_t1 = RG_rl_244 ;
	7'h7f :
		rl_a120_t4_t1 = RG_rl_244 ;
	default :
		rl_a120_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a120_t4_t1 or rl_a120_t5 or FF_i )
	begin
	rl_a120_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a120_t4 = ( ( { 9{ FF_i } } & rl_a120_t5 )
		| ( { 9{ rl_a120_t4_c1 } } & rl_a120_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_59 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h01 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h02 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h03 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h04 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h05 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h06 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h07 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h08 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h09 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h0a :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h0b :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h0c :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h0d :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h0e :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h0f :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h10 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h11 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h12 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h13 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h14 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h15 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h16 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h17 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h18 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h19 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h1a :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h1b :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h1c :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h1d :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h1e :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h1f :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h20 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h21 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h22 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h23 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h24 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h25 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h26 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h27 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h28 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h29 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h2a :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h2b :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h2c :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h2d :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h2e :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h2f :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h30 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h31 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h32 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h33 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h34 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h35 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h36 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h37 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h38 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h39 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h3a :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h3b :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h3c :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h3d :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h3e :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h3f :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h40 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h41 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h42 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h43 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h44 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h45 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h46 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h47 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h48 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h49 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h4a :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h4b :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h4c :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h4d :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h4e :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h4f :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h50 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h51 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h52 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h53 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h54 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h55 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h56 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h57 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h58 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h59 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h5a :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h5b :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h5c :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h5d :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h5e :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h5f :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h60 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h61 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h62 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h63 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h64 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h65 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h66 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h67 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h68 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h69 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h6a :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h6b :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h6c :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h6d :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h6e :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h6f :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h70 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h71 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h72 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h73 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h74 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h75 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h76 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h77 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h78 :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h79 :
		rl_a121_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h7a :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h7b :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h7c :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h7d :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h7e :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	7'h7f :
		rl_a121_t4_t1 = RG_quantized_block_rl_59 ;
	default :
		rl_a121_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a121_t4_t1 or rl_a121_t5 or FF_i )
	begin
	rl_a121_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a121_t4 = ( ( { 9{ FF_i } } & rl_a121_t5 )
		| ( { 9{ rl_a121_t4_c1 } } & rl_a121_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_245 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h01 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h02 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h03 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h04 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h05 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h06 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h07 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h08 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h09 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h0a :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h0b :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h0c :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h0d :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h0e :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h0f :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h10 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h11 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h12 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h13 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h14 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h15 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h16 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h17 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h18 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h19 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h1a :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h1b :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h1c :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h1d :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h1e :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h1f :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h20 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h21 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h22 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h23 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h24 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h25 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h26 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h27 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h28 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h29 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h2a :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h2b :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h2c :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h2d :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h2e :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h2f :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h30 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h31 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h32 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h33 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h34 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h35 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h36 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h37 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h38 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h39 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h3a :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h3b :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h3c :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h3d :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h3e :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h3f :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h40 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h41 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h42 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h43 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h44 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h45 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h46 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h47 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h48 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h49 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h4a :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h4b :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h4c :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h4d :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h4e :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h4f :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h50 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h51 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h52 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h53 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h54 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h55 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h56 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h57 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h58 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h59 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h5a :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h5b :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h5c :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h5d :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h5e :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h5f :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h60 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h61 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h62 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h63 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h64 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h65 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h66 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h67 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h68 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h69 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h6a :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h6b :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h6c :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h6d :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h6e :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h6f :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h70 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h71 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h72 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h73 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h74 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h75 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h76 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h77 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h78 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h79 :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h7a :
		rl_a122_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h7b :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h7c :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h7d :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h7e :
		rl_a122_t4_t1 = RG_rl_245 ;
	7'h7f :
		rl_a122_t4_t1 = RG_rl_245 ;
	default :
		rl_a122_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a122_t4_t1 or rl_a122_t5 or FF_i )
	begin
	rl_a122_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a122_t4 = ( ( { 9{ FF_i } } & rl_a122_t5 )
		| ( { 9{ rl_a122_t4_c1 } } & rl_a122_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_60 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h01 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h02 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h03 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h04 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h05 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h06 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h07 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h08 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h09 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h0a :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h0b :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h0c :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h0d :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h0e :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h0f :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h10 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h11 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h12 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h13 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h14 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h15 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h16 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h17 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h18 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h19 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h1a :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h1b :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h1c :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h1d :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h1e :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h1f :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h20 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h21 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h22 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h23 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h24 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h25 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h26 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h27 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h28 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h29 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h2a :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h2b :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h2c :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h2d :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h2e :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h2f :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h30 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h31 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h32 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h33 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h34 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h35 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h36 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h37 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h38 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h39 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h3a :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h3b :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h3c :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h3d :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h3e :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h3f :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h40 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h41 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h42 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h43 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h44 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h45 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h46 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h47 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h48 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h49 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h4a :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h4b :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h4c :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h4d :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h4e :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h4f :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h50 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h51 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h52 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h53 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h54 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h55 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h56 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h57 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h58 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h59 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h5a :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h5b :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h5c :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h5d :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h5e :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h5f :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h60 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h61 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h62 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h63 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h64 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h65 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h66 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h67 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h68 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h69 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h6a :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h6b :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h6c :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h6d :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h6e :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h6f :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h70 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h71 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h72 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h73 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h74 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h75 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h76 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h77 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h78 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h79 :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h7a :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h7b :
		rl_a123_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h7c :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h7d :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h7e :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	7'h7f :
		rl_a123_t4_t1 = RG_quantized_block_rl_60 ;
	default :
		rl_a123_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a123_t4_t1 or rl_a123_t5 or FF_i )
	begin
	rl_a123_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a123_t4 = ( ( { 9{ FF_i } } & rl_a123_t5 )
		| ( { 9{ rl_a123_t4_c1 } } & rl_a123_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_rl_246 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h01 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h02 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h03 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h04 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h05 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h06 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h07 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h08 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h09 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h0a :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h0b :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h0c :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h0d :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h0e :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h0f :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h10 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h11 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h12 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h13 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h14 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h15 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h16 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h17 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h18 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h19 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h1a :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h1b :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h1c :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h1d :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h1e :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h1f :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h20 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h21 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h22 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h23 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h24 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h25 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h26 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h27 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h28 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h29 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h2a :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h2b :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h2c :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h2d :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h2e :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h2f :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h30 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h31 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h32 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h33 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h34 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h35 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h36 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h37 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h38 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h39 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h3a :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h3b :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h3c :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h3d :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h3e :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h3f :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h40 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h41 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h42 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h43 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h44 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h45 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h46 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h47 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h48 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h49 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h4a :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h4b :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h4c :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h4d :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h4e :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h4f :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h50 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h51 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h52 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h53 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h54 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h55 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h56 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h57 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h58 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h59 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h5a :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h5b :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h5c :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h5d :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h5e :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h5f :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h60 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h61 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h62 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h63 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h64 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h65 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h66 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h67 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h68 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h69 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h6a :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h6b :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h6c :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h6d :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h6e :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h6f :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h70 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h71 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h72 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h73 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h74 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h75 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h76 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h77 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h78 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h79 :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h7a :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h7b :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h7c :
		rl_a124_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h7d :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h7e :
		rl_a124_t4_t1 = RG_rl_246 ;
	7'h7f :
		rl_a124_t4_t1 = RG_rl_246 ;
	default :
		rl_a124_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a124_t4_t1 or rl_a124_t5 or FF_i )
	begin
	rl_a124_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a124_t4 = ( ( { 9{ FF_i } } & rl_a124_t5 )
		| ( { 9{ rl_a124_t4_c1 } } & rl_a124_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_61 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h01 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h02 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h03 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h04 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h05 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h06 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h07 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h08 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h09 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h0a :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h0b :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h0c :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h0d :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h0e :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h0f :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h10 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h11 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h12 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h13 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h14 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h15 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h16 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h17 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h18 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h19 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h1a :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h1b :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h1c :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h1d :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h1e :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h1f :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h20 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h21 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h22 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h23 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h24 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h25 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h26 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h27 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h28 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h29 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h2a :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h2b :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h2c :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h2d :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h2e :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h2f :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h30 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h31 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h32 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h33 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h34 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h35 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h36 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h37 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h38 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h39 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h3a :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h3b :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h3c :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h3d :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h3e :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h3f :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h40 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h41 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h42 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h43 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h44 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h45 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h46 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h47 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h48 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h49 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h4a :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h4b :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h4c :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h4d :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h4e :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h4f :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h50 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h51 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h52 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h53 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h54 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h55 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h56 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h57 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h58 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h59 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h5a :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h5b :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h5c :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h5d :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h5e :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h5f :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h60 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h61 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h62 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h63 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h64 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h65 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h66 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h67 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h68 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h69 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h6a :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h6b :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h6c :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h6d :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h6e :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h6f :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h70 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h71 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h72 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h73 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h74 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h75 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h76 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h77 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h78 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h79 :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h7a :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h7b :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h7c :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h7d :
		rl_a125_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h7e :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	7'h7f :
		rl_a125_t4_t1 = RG_quantized_block_rl_61 ;
	default :
		rl_a125_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a125_t4_t1 or rl_a125_t5 or FF_i )
	begin
	rl_a125_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a125_t4 = ( ( { 9{ FF_i } } & rl_a125_t5 )
		| ( { 9{ rl_a125_t4_c1 } } & rl_a125_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_previous_dc_rl_1 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h01 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h02 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h03 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h04 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h05 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h06 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h07 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h08 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h09 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h0a :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h0b :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h0c :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h0d :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h0e :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h0f :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h10 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h11 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h12 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h13 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h14 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h15 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h16 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h17 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h18 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h19 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h1a :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h1b :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h1c :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h1d :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h1e :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h1f :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h20 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h21 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h22 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h23 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h24 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h25 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h26 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h27 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h28 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h29 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h2a :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h2b :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h2c :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h2d :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h2e :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h2f :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h30 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h31 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h32 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h33 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h34 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h35 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h36 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h37 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h38 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h39 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h3a :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h3b :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h3c :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h3d :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h3e :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h3f :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h40 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h41 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h42 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h43 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h44 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h45 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h46 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h47 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h48 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h49 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h4a :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h4b :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h4c :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h4d :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h4e :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h4f :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h50 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h51 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h52 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h53 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h54 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h55 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h56 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h57 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h58 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h59 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h5a :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h5b :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h5c :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h5d :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h5e :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h5f :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h60 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h61 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h62 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h63 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h64 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h65 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h66 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h67 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h68 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h69 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h6a :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h6b :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h6c :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h6d :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h6e :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h6f :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h70 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h71 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h72 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h73 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h74 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h75 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h76 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h77 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h78 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h79 :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h7a :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h7b :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h7c :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h7d :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	7'h7e :
		rl_a126_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	7'h7f :
		rl_a126_t4_t1 = RG_previous_dc_rl_1 ;
	default :
		rl_a126_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a126_t4_t1 or rl_a126_t5 or FF_i )
	begin
	rl_a126_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a126_t4 = ( ( { 9{ FF_i } } & rl_a126_t5 )
		| ( { 9{ rl_a126_t4_c1 } } & rl_a126_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( zz_RD1 or RG_quantized_block_rl_62 or RG_k_01 )	// line#=../rle.cpp:74
	case ( RG_k_01 )
	7'h00 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h01 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h02 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h03 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h04 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h05 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h06 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h07 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h08 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h09 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h0a :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h0b :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h0c :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h0d :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h0e :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h0f :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h10 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h11 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h12 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h13 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h14 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h15 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h16 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h17 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h18 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h19 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h1a :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h1b :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h1c :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h1d :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h1e :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h1f :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h20 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h21 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h22 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h23 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h24 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h25 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h26 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h27 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h28 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h29 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h2a :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h2b :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h2c :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h2d :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h2e :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h2f :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h30 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h31 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h32 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h33 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h34 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h35 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h36 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h37 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h38 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h39 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h3a :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h3b :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h3c :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h3d :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h3e :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h3f :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h40 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h41 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h42 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h43 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h44 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h45 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h46 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h47 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h48 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h49 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h4a :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h4b :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h4c :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h4d :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h4e :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h4f :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h50 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h51 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h52 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h53 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h54 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h55 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h56 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h57 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h58 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h59 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h5a :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h5b :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h5c :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h5d :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h5e :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h5f :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h60 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h61 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h62 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h63 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h64 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h65 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h66 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h67 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h68 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h69 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h6a :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h6b :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h6c :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h6d :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h6e :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h6f :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h70 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h71 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h72 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h73 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h74 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h75 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h76 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h77 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h78 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h79 :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h7a :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h7b :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h7c :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h7d :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h7e :
		rl_a127_t4_t1 = RG_quantized_block_rl_62 ;
	7'h7f :
		rl_a127_t4_t1 = zz_RD1 ;	// line#=../rle.cpp:74
	default :
		rl_a127_t4_t1 = 9'hx ;
	endcase
always @ ( rl_a127_t4_t1 or rl_a127_t5 or FF_i )
	begin
	rl_a127_t4_c1 = ~FF_i ;	// line#=../rle.cpp:74
	rl_a127_t4 = ( ( { 9{ FF_i } } & rl_a127_t5 )
		| ( { 9{ rl_a127_t4_c1 } } & rl_a127_t4_t1 )	// line#=../rle.cpp:74
		) ;
	end
always @ ( FF_i or FF_len or RG_451 or RG_450 or RG_449 or RG_448 or RG_447 or RG_446 or 
	RG_445 or RG_444 or RG_443 or RG_442 or RG_441 or RG_440 or RG_439 or RG_438 or 
	RG_437 or RG_436 or RG_435 or RG_434 or RG_433 or RG_432 or RG_431 or RG_430 or 
	RG_429 or RG_428 or RG_427 or RG_426 or RG_425 or RG_424 or RG_423 or RG_422 or 
	RG_421 or RG_420 or RG_419 or RG_418 or RG_417 or RG_416 or RG_415 or RG_414 or 
	RG_413 or RG_412 or RG_411 or RG_410 or RG_409 or RG_408 or RG_407 or RG_406 or 
	RG_405 or RG_404 or RG_403 or RG_402 or RG_401 or RG_400 or RG_399 or RG_398 or 
	RG_397 or RG_396 or RG_395 or RG_394 or RG_393 or RG_392 or RG_391 or RG_390 or 
	RG_389 or RG_388 or RG_387 or RG_385 or RG_384 or RG_383 or RG_382 or RG_381 or 
	RG_380 or RG_379 or RG_378 or RG_377 or RG_376 or RG_375 or RG_374 or RG_373 or 
	RG_372 or RG_371 or RG_370 or RG_369 or RG_368 or RG_367 or RG_366 or RG_365 or 
	RG_364 or RG_363 or RG_362 or RG_361 or RG_360 or RG_359 or RG_358 or RG_357 or 
	RG_356 or RG_355 or RG_354 or RG_353 or RG_352 or RG_351 or RG_350 or RG_349 or 
	RG_348 or RG_347 or RG_346 or RG_345 or RG_344 or RG_343 or RG_342 or RG_341 or 
	RG_340 or RG_339 or RG_338 or RG_337 or RG_336 or RG_335 or RG_334 or RG_333 or 
	RG_332 or RG_331 or RG_330 or RG_329 or RG_328 or RG_327 or RG_326 or RG_325 or 
	RG_k_01 )	// line#=../rle.cpp:77,78
	case ( RG_k_01 )
	7'h00 :
		M_02_t_t1 = RG_325 ;	// line#=../rle.cpp:77,78
	7'h01 :
		M_02_t_t1 = RG_326 ;	// line#=../rle.cpp:77,78
	7'h02 :
		M_02_t_t1 = RG_327 ;	// line#=../rle.cpp:77,78
	7'h03 :
		M_02_t_t1 = RG_328 ;	// line#=../rle.cpp:77,78
	7'h04 :
		M_02_t_t1 = RG_329 ;	// line#=../rle.cpp:77,78
	7'h05 :
		M_02_t_t1 = RG_330 ;	// line#=../rle.cpp:77,78
	7'h06 :
		M_02_t_t1 = RG_331 ;	// line#=../rle.cpp:77,78
	7'h07 :
		M_02_t_t1 = RG_332 ;	// line#=../rle.cpp:77,78
	7'h08 :
		M_02_t_t1 = RG_333 ;	// line#=../rle.cpp:77,78
	7'h09 :
		M_02_t_t1 = RG_334 ;	// line#=../rle.cpp:77,78
	7'h0a :
		M_02_t_t1 = RG_335 ;	// line#=../rle.cpp:77,78
	7'h0b :
		M_02_t_t1 = RG_336 ;	// line#=../rle.cpp:77,78
	7'h0c :
		M_02_t_t1 = RG_337 ;	// line#=../rle.cpp:77,78
	7'h0d :
		M_02_t_t1 = RG_338 ;	// line#=../rle.cpp:77,78
	7'h0e :
		M_02_t_t1 = RG_339 ;	// line#=../rle.cpp:77,78
	7'h0f :
		M_02_t_t1 = RG_340 ;	// line#=../rle.cpp:77,78
	7'h10 :
		M_02_t_t1 = RG_341 ;	// line#=../rle.cpp:77,78
	7'h11 :
		M_02_t_t1 = RG_342 ;	// line#=../rle.cpp:77,78
	7'h12 :
		M_02_t_t1 = RG_343 ;	// line#=../rle.cpp:77,78
	7'h13 :
		M_02_t_t1 = RG_344 ;	// line#=../rle.cpp:77,78
	7'h14 :
		M_02_t_t1 = RG_345 ;	// line#=../rle.cpp:77,78
	7'h15 :
		M_02_t_t1 = RG_346 ;	// line#=../rle.cpp:77,78
	7'h16 :
		M_02_t_t1 = RG_347 ;	// line#=../rle.cpp:77,78
	7'h17 :
		M_02_t_t1 = RG_348 ;	// line#=../rle.cpp:77,78
	7'h18 :
		M_02_t_t1 = RG_349 ;	// line#=../rle.cpp:77,78
	7'h19 :
		M_02_t_t1 = RG_350 ;	// line#=../rle.cpp:77,78
	7'h1a :
		M_02_t_t1 = RG_351 ;	// line#=../rle.cpp:77,78
	7'h1b :
		M_02_t_t1 = RG_352 ;	// line#=../rle.cpp:77,78
	7'h1c :
		M_02_t_t1 = RG_353 ;	// line#=../rle.cpp:77,78
	7'h1d :
		M_02_t_t1 = RG_354 ;	// line#=../rle.cpp:77,78
	7'h1e :
		M_02_t_t1 = RG_355 ;	// line#=../rle.cpp:77,78
	7'h1f :
		M_02_t_t1 = RG_356 ;	// line#=../rle.cpp:77,78
	7'h20 :
		M_02_t_t1 = RG_357 ;	// line#=../rle.cpp:77,78
	7'h21 :
		M_02_t_t1 = RG_358 ;	// line#=../rle.cpp:77,78
	7'h22 :
		M_02_t_t1 = RG_359 ;	// line#=../rle.cpp:77,78
	7'h23 :
		M_02_t_t1 = RG_360 ;	// line#=../rle.cpp:77,78
	7'h24 :
		M_02_t_t1 = RG_361 ;	// line#=../rle.cpp:77,78
	7'h25 :
		M_02_t_t1 = RG_362 ;	// line#=../rle.cpp:77,78
	7'h26 :
		M_02_t_t1 = RG_363 ;	// line#=../rle.cpp:77,78
	7'h27 :
		M_02_t_t1 = RG_364 ;	// line#=../rle.cpp:77,78
	7'h28 :
		M_02_t_t1 = RG_365 ;	// line#=../rle.cpp:77,78
	7'h29 :
		M_02_t_t1 = RG_366 ;	// line#=../rle.cpp:77,78
	7'h2a :
		M_02_t_t1 = RG_367 ;	// line#=../rle.cpp:77,78
	7'h2b :
		M_02_t_t1 = RG_368 ;	// line#=../rle.cpp:77,78
	7'h2c :
		M_02_t_t1 = RG_369 ;	// line#=../rle.cpp:77,78
	7'h2d :
		M_02_t_t1 = RG_370 ;	// line#=../rle.cpp:77,78
	7'h2e :
		M_02_t_t1 = RG_371 ;	// line#=../rle.cpp:77,78
	7'h2f :
		M_02_t_t1 = RG_372 ;	// line#=../rle.cpp:77,78
	7'h30 :
		M_02_t_t1 = RG_373 ;	// line#=../rle.cpp:77,78
	7'h31 :
		M_02_t_t1 = RG_374 ;	// line#=../rle.cpp:77,78
	7'h32 :
		M_02_t_t1 = RG_375 ;	// line#=../rle.cpp:77,78
	7'h33 :
		M_02_t_t1 = RG_376 ;	// line#=../rle.cpp:77,78
	7'h34 :
		M_02_t_t1 = RG_377 ;	// line#=../rle.cpp:77,78
	7'h35 :
		M_02_t_t1 = RG_378 ;	// line#=../rle.cpp:77,78
	7'h36 :
		M_02_t_t1 = RG_379 ;	// line#=../rle.cpp:77,78
	7'h37 :
		M_02_t_t1 = RG_380 ;	// line#=../rle.cpp:77,78
	7'h38 :
		M_02_t_t1 = RG_381 ;	// line#=../rle.cpp:77,78
	7'h39 :
		M_02_t_t1 = RG_382 ;	// line#=../rle.cpp:77,78
	7'h3a :
		M_02_t_t1 = RG_383 ;	// line#=../rle.cpp:77,78
	7'h3b :
		M_02_t_t1 = RG_384 ;	// line#=../rle.cpp:77,78
	7'h3c :
		M_02_t_t1 = RG_385 ;	// line#=../rle.cpp:77,78
	7'h3d :
		M_02_t_t1 = RG_387 ;	// line#=../rle.cpp:77,78
	7'h3e :
		M_02_t_t1 = RG_388 ;	// line#=../rle.cpp:77,78
	7'h3f :
		M_02_t_t1 = RG_389 ;	// line#=../rle.cpp:77,78
	7'h40 :
		M_02_t_t1 = RG_390 ;	// line#=../rle.cpp:77,78
	7'h41 :
		M_02_t_t1 = RG_391 ;	// line#=../rle.cpp:77,78
	7'h42 :
		M_02_t_t1 = RG_392 ;	// line#=../rle.cpp:77,78
	7'h43 :
		M_02_t_t1 = RG_393 ;	// line#=../rle.cpp:77,78
	7'h44 :
		M_02_t_t1 = RG_394 ;	// line#=../rle.cpp:77,78
	7'h45 :
		M_02_t_t1 = RG_395 ;	// line#=../rle.cpp:77,78
	7'h46 :
		M_02_t_t1 = RG_396 ;	// line#=../rle.cpp:77,78
	7'h47 :
		M_02_t_t1 = RG_397 ;	// line#=../rle.cpp:77,78
	7'h48 :
		M_02_t_t1 = RG_398 ;	// line#=../rle.cpp:77,78
	7'h49 :
		M_02_t_t1 = RG_399 ;	// line#=../rle.cpp:77,78
	7'h4a :
		M_02_t_t1 = RG_400 ;	// line#=../rle.cpp:77,78
	7'h4b :
		M_02_t_t1 = RG_401 ;	// line#=../rle.cpp:77,78
	7'h4c :
		M_02_t_t1 = RG_402 ;	// line#=../rle.cpp:77,78
	7'h4d :
		M_02_t_t1 = RG_403 ;	// line#=../rle.cpp:77,78
	7'h4e :
		M_02_t_t1 = RG_404 ;	// line#=../rle.cpp:77,78
	7'h4f :
		M_02_t_t1 = RG_405 ;	// line#=../rle.cpp:77,78
	7'h50 :
		M_02_t_t1 = RG_406 ;	// line#=../rle.cpp:77,78
	7'h51 :
		M_02_t_t1 = RG_407 ;	// line#=../rle.cpp:77,78
	7'h52 :
		M_02_t_t1 = RG_408 ;	// line#=../rle.cpp:77,78
	7'h53 :
		M_02_t_t1 = RG_409 ;	// line#=../rle.cpp:77,78
	7'h54 :
		M_02_t_t1 = RG_410 ;	// line#=../rle.cpp:77,78
	7'h55 :
		M_02_t_t1 = RG_411 ;	// line#=../rle.cpp:77,78
	7'h56 :
		M_02_t_t1 = RG_412 ;	// line#=../rle.cpp:77,78
	7'h57 :
		M_02_t_t1 = RG_413 ;	// line#=../rle.cpp:77,78
	7'h58 :
		M_02_t_t1 = RG_414 ;	// line#=../rle.cpp:77,78
	7'h59 :
		M_02_t_t1 = RG_415 ;	// line#=../rle.cpp:77,78
	7'h5a :
		M_02_t_t1 = RG_416 ;	// line#=../rle.cpp:77,78
	7'h5b :
		M_02_t_t1 = RG_417 ;	// line#=../rle.cpp:77,78
	7'h5c :
		M_02_t_t1 = RG_418 ;	// line#=../rle.cpp:77,78
	7'h5d :
		M_02_t_t1 = RG_419 ;	// line#=../rle.cpp:77,78
	7'h5e :
		M_02_t_t1 = RG_420 ;	// line#=../rle.cpp:77,78
	7'h5f :
		M_02_t_t1 = RG_421 ;	// line#=../rle.cpp:77,78
	7'h60 :
		M_02_t_t1 = RG_422 ;	// line#=../rle.cpp:77,78
	7'h61 :
		M_02_t_t1 = RG_423 ;	// line#=../rle.cpp:77,78
	7'h62 :
		M_02_t_t1 = RG_424 ;	// line#=../rle.cpp:77,78
	7'h63 :
		M_02_t_t1 = RG_425 ;	// line#=../rle.cpp:77,78
	7'h64 :
		M_02_t_t1 = RG_426 ;	// line#=../rle.cpp:77,78
	7'h65 :
		M_02_t_t1 = RG_427 ;	// line#=../rle.cpp:77,78
	7'h66 :
		M_02_t_t1 = RG_428 ;	// line#=../rle.cpp:77,78
	7'h67 :
		M_02_t_t1 = RG_429 ;	// line#=../rle.cpp:77,78
	7'h68 :
		M_02_t_t1 = RG_430 ;	// line#=../rle.cpp:77,78
	7'h69 :
		M_02_t_t1 = RG_431 ;	// line#=../rle.cpp:77,78
	7'h6a :
		M_02_t_t1 = RG_432 ;	// line#=../rle.cpp:77,78
	7'h6b :
		M_02_t_t1 = RG_433 ;	// line#=../rle.cpp:77,78
	7'h6c :
		M_02_t_t1 = RG_434 ;	// line#=../rle.cpp:77,78
	7'h6d :
		M_02_t_t1 = RG_435 ;	// line#=../rle.cpp:77,78
	7'h6e :
		M_02_t_t1 = RG_436 ;	// line#=../rle.cpp:77,78
	7'h6f :
		M_02_t_t1 = RG_437 ;	// line#=../rle.cpp:77,78
	7'h70 :
		M_02_t_t1 = RG_438 ;	// line#=../rle.cpp:77,78
	7'h71 :
		M_02_t_t1 = RG_439 ;	// line#=../rle.cpp:77,78
	7'h72 :
		M_02_t_t1 = RG_440 ;	// line#=../rle.cpp:77,78
	7'h73 :
		M_02_t_t1 = RG_441 ;	// line#=../rle.cpp:77,78
	7'h74 :
		M_02_t_t1 = RG_442 ;	// line#=../rle.cpp:77,78
	7'h75 :
		M_02_t_t1 = RG_443 ;	// line#=../rle.cpp:77,78
	7'h76 :
		M_02_t_t1 = RG_444 ;	// line#=../rle.cpp:77,78
	7'h77 :
		M_02_t_t1 = RG_445 ;	// line#=../rle.cpp:77,78
	7'h78 :
		M_02_t_t1 = RG_446 ;	// line#=../rle.cpp:77,78
	7'h79 :
		M_02_t_t1 = RG_447 ;	// line#=../rle.cpp:77,78
	7'h7a :
		M_02_t_t1 = RG_448 ;	// line#=../rle.cpp:77,78
	7'h7b :
		M_02_t_t1 = RG_449 ;	// line#=../rle.cpp:77,78
	7'h7c :
		M_02_t_t1 = RG_450 ;	// line#=../rle.cpp:77,78
	7'h7d :
		M_02_t_t1 = RG_451 ;	// line#=../rle.cpp:77,78
	7'h7e :
		M_02_t_t1 = FF_len ;	// line#=../rle.cpp:77,78
	7'h7f :
		M_02_t_t1 = FF_i ;	// line#=../rle.cpp:77,78
	default :
		M_02_t_t1 = 1'hx ;
	endcase
always @ ( M_02_t_t1 or RG_324 or M_14_t128 )	// line#=../rle.cpp:77,78
	begin
	M_02_t_c1 = ~M_14_t128 ;	// line#=../rle.cpp:77,78
	M_02_t = ( ( { 1{ M_02_t_c1 } } & RG_324 )	// line#=../rle.cpp:77,78
		| ( { 1{ M_14_t128 } } & M_02_t_t1 )	// line#=../rle.cpp:77,78
		) ;
	end
always @ ( RG_rl_127 or RG_rl_126 or RG_rl_125 or RG_rl_124 or RG_rl_123 or RG_rl_122 or 
	RG_rl_121 or RG_rl_120 or RG_rl_119 or RG_rl_118 or RG_rl_117 or RG_rl_116 or 
	RG_rl_115 or RG_rl_114 or RG_rl_113 or RG_rl_112 or RG_rl_111 or RG_rl_110 or 
	RG_rl_109 or RG_rl_108 or RG_rl_107 or RG_rl_106 or RG_rl_105 or RG_rl_104 or 
	RG_rl_103 or RG_rl_102 or RG_rl_101 or RG_rl_100 or RG_rl_99 or RG_rl_98 or 
	RG_rl_97 or RG_rl_96 or RG_rl_95 or RG_rl_94 or RG_rl_93 or RG_rl_92 or 
	RG_rl_91 or RG_rl_90 or RG_rl_89 or RG_rl_88 or RG_rl_87 or RG_rl_86 or 
	RG_rl_85 or RG_rl_84 or RG_rl_83 or RG_rl_82 or RG_rl_81 or RG_rl_80 or 
	RG_rl_79 or RG_rl_78 or RG_rl_77 or RG_rl_76 or RG_rl_75 or RG_rl_74 or 
	RG_rl_73 or RG_rl_72 or RG_rl_71 or RG_rl_70 or RG_rl_69 or RG_rl_68 or 
	RG_rl_67 or RG_rl_66 or RG_rl_65 or RG_rl_64 or RG_rl_63 or RG_rl_62 or 
	RG_rl_61 or RG_rl_60 or RG_rl_59 or RG_rl_58 or RG_rl_57 or RG_rl_56 or 
	RG_rl_55 or RG_rl_54 or RG_rl_53 or RG_rl_52 or RG_rl_51 or RG_rl_50 or 
	RG_rl_49 or RG_rl_48 or RG_rl_47 or RG_rl_46 or RG_rl_45 or RG_rl_44 or 
	RG_rl_43 or RG_rl_42 or RG_rl_41 or RG_rl_40 or RG_rl_39 or RG_rl_38 or 
	RG_rl_37 or RG_rl_36 or RG_rl_35 or RG_rl_34 or RG_rl_33 or RG_rl_32 or 
	RG_rl_31 or RG_rl_30 or RG_rl_29 or RG_rl_28 or RG_rl_27 or RG_rl_26 or 
	RG_rl_25 or RG_rl_24 or RG_rl_23 or RG_rl_22 or RG_rl_21 or RG_rl_20 or 
	RG_rl_19 or RG_rl_18 or RG_rl_17 or RG_rl_16 or RG_rl_15 or RG_rl_14 or 
	RG_rl_13 or RG_rl_12 or RG_rl_11 or RG_rl_10 or RG_rl_9 or RG_rl_8 or RG_rl_7 or 
	RG_rl_6 or RG_rl_5 or RG_rl_4 or RG_rl_3 or RG_rl_2 or RG_rl_1 or RG_rl or 
	sub8u_7_11ot )	// line#=../rle.cpp:83,84
	case ( sub8u_7_11ot )
	7'h00 :
		M_03_t128_t1 = ~|RG_rl ;	// line#=../rle.cpp:83,84
	7'h01 :
		M_03_t128_t1 = ~|RG_rl_1 ;	// line#=../rle.cpp:83,84
	7'h02 :
		M_03_t128_t1 = ~|RG_rl_2 ;	// line#=../rle.cpp:83,84
	7'h03 :
		M_03_t128_t1 = ~|RG_rl_3 ;	// line#=../rle.cpp:83,84
	7'h04 :
		M_03_t128_t1 = ~|RG_rl_4 ;	// line#=../rle.cpp:83,84
	7'h05 :
		M_03_t128_t1 = ~|RG_rl_5 ;	// line#=../rle.cpp:83,84
	7'h06 :
		M_03_t128_t1 = ~|RG_rl_6 ;	// line#=../rle.cpp:83,84
	7'h07 :
		M_03_t128_t1 = ~|RG_rl_7 ;	// line#=../rle.cpp:83,84
	7'h08 :
		M_03_t128_t1 = ~|RG_rl_8 ;	// line#=../rle.cpp:83,84
	7'h09 :
		M_03_t128_t1 = ~|RG_rl_9 ;	// line#=../rle.cpp:83,84
	7'h0a :
		M_03_t128_t1 = ~|RG_rl_10 ;	// line#=../rle.cpp:83,84
	7'h0b :
		M_03_t128_t1 = ~|RG_rl_11 ;	// line#=../rle.cpp:83,84
	7'h0c :
		M_03_t128_t1 = ~|RG_rl_12 ;	// line#=../rle.cpp:83,84
	7'h0d :
		M_03_t128_t1 = ~|RG_rl_13 ;	// line#=../rle.cpp:83,84
	7'h0e :
		M_03_t128_t1 = ~|RG_rl_14 ;	// line#=../rle.cpp:83,84
	7'h0f :
		M_03_t128_t1 = ~|RG_rl_15 ;	// line#=../rle.cpp:83,84
	7'h10 :
		M_03_t128_t1 = ~|RG_rl_16 ;	// line#=../rle.cpp:83,84
	7'h11 :
		M_03_t128_t1 = ~|RG_rl_17 ;	// line#=../rle.cpp:83,84
	7'h12 :
		M_03_t128_t1 = ~|RG_rl_18 ;	// line#=../rle.cpp:83,84
	7'h13 :
		M_03_t128_t1 = ~|RG_rl_19 ;	// line#=../rle.cpp:83,84
	7'h14 :
		M_03_t128_t1 = ~|RG_rl_20 ;	// line#=../rle.cpp:83,84
	7'h15 :
		M_03_t128_t1 = ~|RG_rl_21 ;	// line#=../rle.cpp:83,84
	7'h16 :
		M_03_t128_t1 = ~|RG_rl_22 ;	// line#=../rle.cpp:83,84
	7'h17 :
		M_03_t128_t1 = ~|RG_rl_23 ;	// line#=../rle.cpp:83,84
	7'h18 :
		M_03_t128_t1 = ~|RG_rl_24 ;	// line#=../rle.cpp:83,84
	7'h19 :
		M_03_t128_t1 = ~|RG_rl_25 ;	// line#=../rle.cpp:83,84
	7'h1a :
		M_03_t128_t1 = ~|RG_rl_26 ;	// line#=../rle.cpp:83,84
	7'h1b :
		M_03_t128_t1 = ~|RG_rl_27 ;	// line#=../rle.cpp:83,84
	7'h1c :
		M_03_t128_t1 = ~|RG_rl_28 ;	// line#=../rle.cpp:83,84
	7'h1d :
		M_03_t128_t1 = ~|RG_rl_29 ;	// line#=../rle.cpp:83,84
	7'h1e :
		M_03_t128_t1 = ~|RG_rl_30 ;	// line#=../rle.cpp:83,84
	7'h1f :
		M_03_t128_t1 = ~|RG_rl_31 ;	// line#=../rle.cpp:83,84
	7'h20 :
		M_03_t128_t1 = ~|RG_rl_32 ;	// line#=../rle.cpp:83,84
	7'h21 :
		M_03_t128_t1 = ~|RG_rl_33 ;	// line#=../rle.cpp:83,84
	7'h22 :
		M_03_t128_t1 = ~|RG_rl_34 ;	// line#=../rle.cpp:83,84
	7'h23 :
		M_03_t128_t1 = ~|RG_rl_35 ;	// line#=../rle.cpp:83,84
	7'h24 :
		M_03_t128_t1 = ~|RG_rl_36 ;	// line#=../rle.cpp:83,84
	7'h25 :
		M_03_t128_t1 = ~|RG_rl_37 ;	// line#=../rle.cpp:83,84
	7'h26 :
		M_03_t128_t1 = ~|RG_rl_38 ;	// line#=../rle.cpp:83,84
	7'h27 :
		M_03_t128_t1 = ~|RG_rl_39 ;	// line#=../rle.cpp:83,84
	7'h28 :
		M_03_t128_t1 = ~|RG_rl_40 ;	// line#=../rle.cpp:83,84
	7'h29 :
		M_03_t128_t1 = ~|RG_rl_41 ;	// line#=../rle.cpp:83,84
	7'h2a :
		M_03_t128_t1 = ~|RG_rl_42 ;	// line#=../rle.cpp:83,84
	7'h2b :
		M_03_t128_t1 = ~|RG_rl_43 ;	// line#=../rle.cpp:83,84
	7'h2c :
		M_03_t128_t1 = ~|RG_rl_44 ;	// line#=../rle.cpp:83,84
	7'h2d :
		M_03_t128_t1 = ~|RG_rl_45 ;	// line#=../rle.cpp:83,84
	7'h2e :
		M_03_t128_t1 = ~|RG_rl_46 ;	// line#=../rle.cpp:83,84
	7'h2f :
		M_03_t128_t1 = ~|RG_rl_47 ;	// line#=../rle.cpp:83,84
	7'h30 :
		M_03_t128_t1 = ~|RG_rl_48 ;	// line#=../rle.cpp:83,84
	7'h31 :
		M_03_t128_t1 = ~|RG_rl_49 ;	// line#=../rle.cpp:83,84
	7'h32 :
		M_03_t128_t1 = ~|RG_rl_50 ;	// line#=../rle.cpp:83,84
	7'h33 :
		M_03_t128_t1 = ~|RG_rl_51 ;	// line#=../rle.cpp:83,84
	7'h34 :
		M_03_t128_t1 = ~|RG_rl_52 ;	// line#=../rle.cpp:83,84
	7'h35 :
		M_03_t128_t1 = ~|RG_rl_53 ;	// line#=../rle.cpp:83,84
	7'h36 :
		M_03_t128_t1 = ~|RG_rl_54 ;	// line#=../rle.cpp:83,84
	7'h37 :
		M_03_t128_t1 = ~|RG_rl_55 ;	// line#=../rle.cpp:83,84
	7'h38 :
		M_03_t128_t1 = ~|RG_rl_56 ;	// line#=../rle.cpp:83,84
	7'h39 :
		M_03_t128_t1 = ~|RG_rl_57 ;	// line#=../rle.cpp:83,84
	7'h3a :
		M_03_t128_t1 = ~|RG_rl_58 ;	// line#=../rle.cpp:83,84
	7'h3b :
		M_03_t128_t1 = ~|RG_rl_59 ;	// line#=../rle.cpp:83,84
	7'h3c :
		M_03_t128_t1 = ~|RG_rl_60 ;	// line#=../rle.cpp:83,84
	7'h3d :
		M_03_t128_t1 = ~|RG_rl_61 ;	// line#=../rle.cpp:83,84
	7'h3e :
		M_03_t128_t1 = ~|RG_rl_62 ;	// line#=../rle.cpp:83,84
	7'h3f :
		M_03_t128_t1 = ~|RG_rl_63 ;	// line#=../rle.cpp:83,84
	7'h40 :
		M_03_t128_t1 = ~|RG_rl_64 ;	// line#=../rle.cpp:83,84
	7'h41 :
		M_03_t128_t1 = ~|RG_rl_65 ;	// line#=../rle.cpp:83,84
	7'h42 :
		M_03_t128_t1 = ~|RG_rl_66 ;	// line#=../rle.cpp:83,84
	7'h43 :
		M_03_t128_t1 = ~|RG_rl_67 ;	// line#=../rle.cpp:83,84
	7'h44 :
		M_03_t128_t1 = ~|RG_rl_68 ;	// line#=../rle.cpp:83,84
	7'h45 :
		M_03_t128_t1 = ~|RG_rl_69 ;	// line#=../rle.cpp:83,84
	7'h46 :
		M_03_t128_t1 = ~|RG_rl_70 ;	// line#=../rle.cpp:83,84
	7'h47 :
		M_03_t128_t1 = ~|RG_rl_71 ;	// line#=../rle.cpp:83,84
	7'h48 :
		M_03_t128_t1 = ~|RG_rl_72 ;	// line#=../rle.cpp:83,84
	7'h49 :
		M_03_t128_t1 = ~|RG_rl_73 ;	// line#=../rle.cpp:83,84
	7'h4a :
		M_03_t128_t1 = ~|RG_rl_74 ;	// line#=../rle.cpp:83,84
	7'h4b :
		M_03_t128_t1 = ~|RG_rl_75 ;	// line#=../rle.cpp:83,84
	7'h4c :
		M_03_t128_t1 = ~|RG_rl_76 ;	// line#=../rle.cpp:83,84
	7'h4d :
		M_03_t128_t1 = ~|RG_rl_77 ;	// line#=../rle.cpp:83,84
	7'h4e :
		M_03_t128_t1 = ~|RG_rl_78 ;	// line#=../rle.cpp:83,84
	7'h4f :
		M_03_t128_t1 = ~|RG_rl_79 ;	// line#=../rle.cpp:83,84
	7'h50 :
		M_03_t128_t1 = ~|RG_rl_80 ;	// line#=../rle.cpp:83,84
	7'h51 :
		M_03_t128_t1 = ~|RG_rl_81 ;	// line#=../rle.cpp:83,84
	7'h52 :
		M_03_t128_t1 = ~|RG_rl_82 ;	// line#=../rle.cpp:83,84
	7'h53 :
		M_03_t128_t1 = ~|RG_rl_83 ;	// line#=../rle.cpp:83,84
	7'h54 :
		M_03_t128_t1 = ~|RG_rl_84 ;	// line#=../rle.cpp:83,84
	7'h55 :
		M_03_t128_t1 = ~|RG_rl_85 ;	// line#=../rle.cpp:83,84
	7'h56 :
		M_03_t128_t1 = ~|RG_rl_86 ;	// line#=../rle.cpp:83,84
	7'h57 :
		M_03_t128_t1 = ~|RG_rl_87 ;	// line#=../rle.cpp:83,84
	7'h58 :
		M_03_t128_t1 = ~|RG_rl_88 ;	// line#=../rle.cpp:83,84
	7'h59 :
		M_03_t128_t1 = ~|RG_rl_89 ;	// line#=../rle.cpp:83,84
	7'h5a :
		M_03_t128_t1 = ~|RG_rl_90 ;	// line#=../rle.cpp:83,84
	7'h5b :
		M_03_t128_t1 = ~|RG_rl_91 ;	// line#=../rle.cpp:83,84
	7'h5c :
		M_03_t128_t1 = ~|RG_rl_92 ;	// line#=../rle.cpp:83,84
	7'h5d :
		M_03_t128_t1 = ~|RG_rl_93 ;	// line#=../rle.cpp:83,84
	7'h5e :
		M_03_t128_t1 = ~|RG_rl_94 ;	// line#=../rle.cpp:83,84
	7'h5f :
		M_03_t128_t1 = ~|RG_rl_95 ;	// line#=../rle.cpp:83,84
	7'h60 :
		M_03_t128_t1 = ~|RG_rl_96 ;	// line#=../rle.cpp:83,84
	7'h61 :
		M_03_t128_t1 = ~|RG_rl_97 ;	// line#=../rle.cpp:83,84
	7'h62 :
		M_03_t128_t1 = ~|RG_rl_98 ;	// line#=../rle.cpp:83,84
	7'h63 :
		M_03_t128_t1 = ~|RG_rl_99 ;	// line#=../rle.cpp:83,84
	7'h64 :
		M_03_t128_t1 = ~|RG_rl_100 ;	// line#=../rle.cpp:83,84
	7'h65 :
		M_03_t128_t1 = ~|RG_rl_101 ;	// line#=../rle.cpp:83,84
	7'h66 :
		M_03_t128_t1 = ~|RG_rl_102 ;	// line#=../rle.cpp:83,84
	7'h67 :
		M_03_t128_t1 = ~|RG_rl_103 ;	// line#=../rle.cpp:83,84
	7'h68 :
		M_03_t128_t1 = ~|RG_rl_104 ;	// line#=../rle.cpp:83,84
	7'h69 :
		M_03_t128_t1 = ~|RG_rl_105 ;	// line#=../rle.cpp:83,84
	7'h6a :
		M_03_t128_t1 = ~|RG_rl_106 ;	// line#=../rle.cpp:83,84
	7'h6b :
		M_03_t128_t1 = ~|RG_rl_107 ;	// line#=../rle.cpp:83,84
	7'h6c :
		M_03_t128_t1 = ~|RG_rl_108 ;	// line#=../rle.cpp:83,84
	7'h6d :
		M_03_t128_t1 = ~|RG_rl_109 ;	// line#=../rle.cpp:83,84
	7'h6e :
		M_03_t128_t1 = ~|RG_rl_110 ;	// line#=../rle.cpp:83,84
	7'h6f :
		M_03_t128_t1 = ~|RG_rl_111 ;	// line#=../rle.cpp:83,84
	7'h70 :
		M_03_t128_t1 = ~|RG_rl_112 ;	// line#=../rle.cpp:83,84
	7'h71 :
		M_03_t128_t1 = ~|RG_rl_113 ;	// line#=../rle.cpp:83,84
	7'h72 :
		M_03_t128_t1 = ~|RG_rl_114 ;	// line#=../rle.cpp:83,84
	7'h73 :
		M_03_t128_t1 = ~|RG_rl_115 ;	// line#=../rle.cpp:83,84
	7'h74 :
		M_03_t128_t1 = ~|RG_rl_116 ;	// line#=../rle.cpp:83,84
	7'h75 :
		M_03_t128_t1 = ~|RG_rl_117 ;	// line#=../rle.cpp:83,84
	7'h76 :
		M_03_t128_t1 = ~|RG_rl_118 ;	// line#=../rle.cpp:83,84
	7'h77 :
		M_03_t128_t1 = ~|RG_rl_119 ;	// line#=../rle.cpp:83,84
	7'h78 :
		M_03_t128_t1 = ~|RG_rl_120 ;	// line#=../rle.cpp:83,84
	7'h79 :
		M_03_t128_t1 = ~|RG_rl_121 ;	// line#=../rle.cpp:83,84
	7'h7a :
		M_03_t128_t1 = ~|RG_rl_122 ;	// line#=../rle.cpp:83,84
	7'h7b :
		M_03_t128_t1 = ~|RG_rl_123 ;	// line#=../rle.cpp:83,84
	7'h7c :
		M_03_t128_t1 = ~|RG_rl_124 ;	// line#=../rle.cpp:83,84
	7'h7d :
		M_03_t128_t1 = ~|RG_rl_125 ;	// line#=../rle.cpp:83,84
	7'h7e :
		M_03_t128_t1 = ~|RG_rl_126 ;	// line#=../rle.cpp:83,84
	7'h7f :
		M_03_t128_t1 = ~|RG_rl_127 ;	// line#=../rle.cpp:83,84
	default :
		M_03_t128_t1 = 1'hx ;
	endcase
always @ ( M_03_t128_t1 or M_15_t128 )	// line#=../rle.cpp:83,84
	M_03_t128 = ( { 1{ M_15_t128 } } & M_03_t128_t1 )	// line#=../rle.cpp:83,84
		 ;	// line#=../rle.cpp:83,84
assign	JF_06 = ~M_03_t128 ;
assign	jpeg_out_a00_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a00_r_en )
		jpeg_out_a00_r <= RG_rl ;
assign	jpeg_out_a01_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a01_r_en )
		jpeg_out_a01_r <= RG_rl_1 ;
assign	jpeg_out_a02_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a02_r_en )
		jpeg_out_a02_r <= RG_rl_2 ;
assign	jpeg_out_a03_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a03_r_en )
		jpeg_out_a03_r <= RG_rl_3 ;
assign	jpeg_out_a04_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a04_r_en )
		jpeg_out_a04_r <= RG_rl_4 ;
assign	jpeg_out_a05_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a05_r_en )
		jpeg_out_a05_r <= RG_rl_5 ;
assign	jpeg_out_a06_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a06_r_en )
		jpeg_out_a06_r <= RG_rl_6 ;
assign	jpeg_out_a07_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a07_r_en )
		jpeg_out_a07_r <= RG_rl_7 ;
assign	jpeg_out_a08_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a08_r_en )
		jpeg_out_a08_r <= RG_rl_8 ;
assign	jpeg_out_a09_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a09_r_en )
		jpeg_out_a09_r <= RG_rl_9 ;
assign	jpeg_out_a10_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a10_r_en )
		jpeg_out_a10_r <= RG_rl_10 ;
assign	jpeg_out_a11_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a11_r_en )
		jpeg_out_a11_r <= RG_rl_11 ;
assign	jpeg_out_a12_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a12_r_en )
		jpeg_out_a12_r <= RG_rl_12 ;
assign	jpeg_out_a13_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a13_r_en )
		jpeg_out_a13_r <= RG_rl_13 ;
assign	jpeg_out_a14_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a14_r_en )
		jpeg_out_a14_r <= RG_rl_14 ;
assign	jpeg_out_a15_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a15_r_en )
		jpeg_out_a15_r <= RG_rl_15 ;
assign	jpeg_out_a16_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a16_r_en )
		jpeg_out_a16_r <= RG_rl_16 ;
assign	jpeg_out_a17_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a17_r_en )
		jpeg_out_a17_r <= RG_rl_17 ;
assign	jpeg_out_a18_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a18_r_en )
		jpeg_out_a18_r <= RG_rl_18 ;
assign	jpeg_out_a19_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a19_r_en )
		jpeg_out_a19_r <= RG_rl_19 ;
assign	jpeg_out_a20_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a20_r_en )
		jpeg_out_a20_r <= RG_rl_20 ;
assign	jpeg_out_a21_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a21_r_en )
		jpeg_out_a21_r <= RG_rl_21 ;
assign	jpeg_out_a22_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a22_r_en )
		jpeg_out_a22_r <= RG_rl_22 ;
assign	jpeg_out_a23_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a23_r_en )
		jpeg_out_a23_r <= RG_rl_23 ;
assign	jpeg_out_a24_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a24_r_en )
		jpeg_out_a24_r <= RG_rl_24 ;
assign	jpeg_out_a25_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a25_r_en )
		jpeg_out_a25_r <= RG_rl_25 ;
assign	jpeg_out_a26_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a26_r_en )
		jpeg_out_a26_r <= RG_rl_26 ;
assign	jpeg_out_a27_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a27_r_en )
		jpeg_out_a27_r <= RG_rl_27 ;
assign	jpeg_out_a28_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a28_r_en )
		jpeg_out_a28_r <= RG_rl_28 ;
assign	jpeg_out_a29_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a29_r_en )
		jpeg_out_a29_r <= RG_rl_29 ;
assign	jpeg_out_a30_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a30_r_en )
		jpeg_out_a30_r <= RG_rl_30 ;
assign	jpeg_out_a31_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a31_r_en )
		jpeg_out_a31_r <= RG_rl_31 ;
assign	jpeg_out_a32_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a32_r_en )
		jpeg_out_a32_r <= RG_rl_32 ;
assign	jpeg_out_a33_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a33_r_en )
		jpeg_out_a33_r <= RG_rl_33 ;
assign	jpeg_out_a34_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a34_r_en )
		jpeg_out_a34_r <= RG_rl_34 ;
assign	jpeg_out_a35_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a35_r_en )
		jpeg_out_a35_r <= RG_rl_35 ;
assign	jpeg_out_a36_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a36_r_en )
		jpeg_out_a36_r <= RG_rl_36 ;
assign	jpeg_out_a37_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a37_r_en )
		jpeg_out_a37_r <= RG_rl_37 ;
assign	jpeg_out_a38_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a38_r_en )
		jpeg_out_a38_r <= RG_rl_38 ;
assign	jpeg_out_a39_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a39_r_en )
		jpeg_out_a39_r <= RG_rl_39 ;
assign	jpeg_out_a40_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a40_r_en )
		jpeg_out_a40_r <= RG_rl_40 ;
assign	jpeg_out_a41_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a41_r_en )
		jpeg_out_a41_r <= RG_rl_41 ;
assign	jpeg_out_a42_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a42_r_en )
		jpeg_out_a42_r <= RG_rl_42 ;
assign	jpeg_out_a43_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a43_r_en )
		jpeg_out_a43_r <= RG_rl_43 ;
assign	jpeg_out_a44_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a44_r_en )
		jpeg_out_a44_r <= RG_rl_44 ;
assign	jpeg_out_a45_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a45_r_en )
		jpeg_out_a45_r <= RG_rl_45 ;
assign	jpeg_out_a46_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a46_r_en )
		jpeg_out_a46_r <= RG_rl_46 ;
assign	jpeg_out_a47_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a47_r_en )
		jpeg_out_a47_r <= RG_rl_47 ;
assign	jpeg_out_a48_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a48_r_en )
		jpeg_out_a48_r <= RG_rl_48 ;
assign	jpeg_out_a49_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a49_r_en )
		jpeg_out_a49_r <= RG_rl_49 ;
assign	jpeg_out_a50_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a50_r_en )
		jpeg_out_a50_r <= RG_rl_50 ;
assign	jpeg_out_a51_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a51_r_en )
		jpeg_out_a51_r <= RG_rl_51 ;
assign	jpeg_out_a52_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a52_r_en )
		jpeg_out_a52_r <= RG_rl_52 ;
assign	jpeg_out_a53_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a53_r_en )
		jpeg_out_a53_r <= RG_rl_53 ;
assign	jpeg_out_a54_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a54_r_en )
		jpeg_out_a54_r <= RG_rl_54 ;
assign	jpeg_out_a55_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a55_r_en )
		jpeg_out_a55_r <= RG_rl_55 ;
assign	jpeg_out_a56_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a56_r_en )
		jpeg_out_a56_r <= RG_rl_56 ;
assign	jpeg_out_a57_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a57_r_en )
		jpeg_out_a57_r <= RG_rl_57 ;
assign	jpeg_out_a58_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a58_r_en )
		jpeg_out_a58_r <= RG_rl_58 ;
assign	jpeg_out_a59_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a59_r_en )
		jpeg_out_a59_r <= RG_rl_59 ;
assign	jpeg_out_a60_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a60_r_en )
		jpeg_out_a60_r <= RG_rl_60 ;
assign	jpeg_out_a61_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a61_r_en )
		jpeg_out_a61_r <= RG_rl_61 ;
assign	jpeg_out_a62_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a62_r_en )
		jpeg_out_a62_r <= RG_rl_62 ;
assign	jpeg_out_a63_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a63_r_en )
		jpeg_out_a63_r <= RG_rl_63 ;
assign	jpeg_out_a64_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a64_r_en )
		jpeg_out_a64_r <= RG_rl_64 ;
assign	jpeg_out_a65_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a65_r_en )
		jpeg_out_a65_r <= RG_rl_65 ;
assign	jpeg_out_a66_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a66_r_en )
		jpeg_out_a66_r <= RG_rl_66 ;
assign	jpeg_out_a67_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a67_r_en )
		jpeg_out_a67_r <= RG_rl_67 ;
assign	jpeg_out_a68_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a68_r_en )
		jpeg_out_a68_r <= RG_rl_68 ;
assign	jpeg_out_a69_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a69_r_en )
		jpeg_out_a69_r <= RG_rl_69 ;
assign	jpeg_out_a70_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a70_r_en )
		jpeg_out_a70_r <= RG_rl_70 ;
assign	jpeg_out_a71_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a71_r_en )
		jpeg_out_a71_r <= RG_rl_71 ;
assign	jpeg_out_a72_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a72_r_en )
		jpeg_out_a72_r <= RG_rl_72 ;
assign	jpeg_out_a73_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a73_r_en )
		jpeg_out_a73_r <= RG_rl_73 ;
assign	jpeg_out_a74_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a74_r_en )
		jpeg_out_a74_r <= RG_rl_74 ;
assign	jpeg_out_a75_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a75_r_en )
		jpeg_out_a75_r <= RG_rl_75 ;
assign	jpeg_out_a76_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a76_r_en )
		jpeg_out_a76_r <= RG_rl_76 ;
assign	jpeg_out_a77_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a77_r_en )
		jpeg_out_a77_r <= RG_rl_77 ;
assign	jpeg_out_a78_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a78_r_en )
		jpeg_out_a78_r <= RG_rl_78 ;
assign	jpeg_out_a79_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a79_r_en )
		jpeg_out_a79_r <= RG_rl_79 ;
assign	jpeg_out_a80_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a80_r_en )
		jpeg_out_a80_r <= RG_rl_80 ;
assign	jpeg_out_a81_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a81_r_en )
		jpeg_out_a81_r <= RG_rl_81 ;
assign	jpeg_out_a82_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a82_r_en )
		jpeg_out_a82_r <= RG_rl_82 ;
assign	jpeg_out_a83_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a83_r_en )
		jpeg_out_a83_r <= RG_rl_83 ;
assign	jpeg_out_a84_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a84_r_en )
		jpeg_out_a84_r <= RG_rl_84 ;
assign	jpeg_out_a85_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a85_r_en )
		jpeg_out_a85_r <= RG_rl_85 ;
assign	jpeg_out_a86_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a86_r_en )
		jpeg_out_a86_r <= RG_rl_86 ;
assign	jpeg_out_a87_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a87_r_en )
		jpeg_out_a87_r <= RG_rl_87 ;
assign	jpeg_out_a88_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a88_r_en )
		jpeg_out_a88_r <= RG_rl_88 ;
assign	jpeg_out_a89_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a89_r_en )
		jpeg_out_a89_r <= RG_rl_89 ;
assign	jpeg_out_a90_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a90_r_en )
		jpeg_out_a90_r <= RG_rl_90 ;
assign	jpeg_out_a91_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a91_r_en )
		jpeg_out_a91_r <= RG_rl_91 ;
assign	jpeg_out_a92_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a92_r_en )
		jpeg_out_a92_r <= RG_rl_92 ;
assign	jpeg_out_a93_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a93_r_en )
		jpeg_out_a93_r <= RG_rl_93 ;
assign	jpeg_out_a94_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a94_r_en )
		jpeg_out_a94_r <= RG_rl_94 ;
assign	jpeg_out_a95_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a95_r_en )
		jpeg_out_a95_r <= RG_rl_95 ;
assign	jpeg_out_a96_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a96_r_en )
		jpeg_out_a96_r <= RG_rl_96 ;
assign	jpeg_out_a97_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a97_r_en )
		jpeg_out_a97_r <= RG_rl_97 ;
assign	jpeg_out_a98_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a98_r_en )
		jpeg_out_a98_r <= RG_rl_98 ;
assign	jpeg_out_a99_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a99_r_en )
		jpeg_out_a99_r <= RG_rl_99 ;
assign	jpeg_out_a100_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a100_r_en )
		jpeg_out_a100_r <= RG_rl_100 ;
assign	jpeg_out_a101_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a101_r_en )
		jpeg_out_a101_r <= RG_rl_101 ;
assign	jpeg_out_a102_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a102_r_en )
		jpeg_out_a102_r <= RG_rl_102 ;
assign	jpeg_out_a103_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a103_r_en )
		jpeg_out_a103_r <= RG_rl_103 ;
assign	jpeg_out_a104_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a104_r_en )
		jpeg_out_a104_r <= RG_rl_104 ;
assign	jpeg_out_a105_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a105_r_en )
		jpeg_out_a105_r <= RG_rl_105 ;
assign	jpeg_out_a106_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a106_r_en )
		jpeg_out_a106_r <= RG_rl_106 ;
assign	jpeg_out_a107_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a107_r_en )
		jpeg_out_a107_r <= RG_rl_107 ;
assign	jpeg_out_a108_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a108_r_en )
		jpeg_out_a108_r <= RG_rl_108 ;
assign	jpeg_out_a109_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a109_r_en )
		jpeg_out_a109_r <= RG_rl_109 ;
assign	jpeg_out_a110_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a110_r_en )
		jpeg_out_a110_r <= RG_rl_110 ;
assign	jpeg_out_a111_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a111_r_en )
		jpeg_out_a111_r <= RG_rl_111 ;
assign	jpeg_out_a112_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a112_r_en )
		jpeg_out_a112_r <= RG_rl_112 ;
assign	jpeg_out_a113_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a113_r_en )
		jpeg_out_a113_r <= RG_rl_113 ;
assign	jpeg_out_a114_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a114_r_en )
		jpeg_out_a114_r <= RG_rl_114 ;
assign	jpeg_out_a115_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a115_r_en )
		jpeg_out_a115_r <= RG_rl_115 ;
assign	jpeg_out_a116_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a116_r_en )
		jpeg_out_a116_r <= RG_rl_116 ;
assign	jpeg_out_a117_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a117_r_en )
		jpeg_out_a117_r <= RG_rl_117 ;
assign	jpeg_out_a118_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a118_r_en )
		jpeg_out_a118_r <= RG_rl_118 ;
assign	jpeg_out_a119_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a119_r_en )
		jpeg_out_a119_r <= RG_rl_119 ;
assign	jpeg_out_a120_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a120_r_en )
		jpeg_out_a120_r <= RG_rl_120 ;
assign	jpeg_out_a121_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a121_r_en )
		jpeg_out_a121_r <= RG_rl_121 ;
assign	jpeg_out_a122_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a122_r_en )
		jpeg_out_a122_r <= RG_rl_122 ;
assign	jpeg_out_a123_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a123_r_en )
		jpeg_out_a123_r <= RG_rl_123 ;
assign	jpeg_out_a124_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a124_r_en )
		jpeg_out_a124_r <= RG_rl_124 ;
assign	jpeg_out_a125_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a125_r_en )
		jpeg_out_a125_r <= RG_rl_125 ;
assign	jpeg_out_a126_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a126_r_en )
		jpeg_out_a126_r <= RG_rl_126 ;
assign	jpeg_out_a127_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:91
	if ( jpeg_out_a127_r_en )
		jpeg_out_a127_r <= RG_rl_127 ;
assign	jpeg_len_out_r_en = U_572 ;
always @ ( posedge clk )	// line#=../rle.cpp:93
	if ( jpeg_len_out_r_en )
		jpeg_len_out_r <= { 4'h0 , RG_len } ;
always @ ( U_572 )
	valid_r_t = ( { 1{ U_572 } } & 1'h1 )	// line#=../rle.cpp:95
		 ;	// line#=../rle.cpp:30
assign	valid_r_en = ( ST1_01d | U_572 ) ;
always @ ( posedge clk )
	if ( valid_r_en )
		valid_r <= valid_r_t ;	// line#=../rle.cpp:30,95
always @ ( RG_len or U_571 or len1_t3 or RG_315 or ST1_09d )	// line#=../rle.cpp:57,58
	begin
	sub8u1i1_c1 = ( ST1_09d & ( ~RG_315 ) ) ;	// line#=../rle.cpp:77,78
	sub8u1i1 = ( ( { 8{ sub8u1i1_c1 } } & { 1'h0 , len1_t3 [6:0] } )	// line#=../rle.cpp:77,78
		| ( { 8{ U_571 } } & RG_len )					// line#=../rle.cpp:86
		) ;
	end
assign	sub8u1i2 = 2'h2 ;	// line#=../rle.cpp:77,78,86
assign	incr8u1i1 = RG_len ;	// line#=../rle.cpp:68,73,79
always @ ( RG_len or FF_i or ST1_09d or RG_k_01 or U_87 or U_05 )	// line#=../rle.cpp:66,67
	begin
	incr8u3i1_c1 = ( U_05 | U_87 ) ;	// line#=../rle.cpp:111,140,141,142
	incr8u3i1_c2 = ( ST1_09d & ( ~FF_i ) ) ;	// line#=../rle.cpp:74
	incr8u3i1 = ( ( { 8{ incr8u3i1_c1 } } & { 2'h0 , RG_k_01 [5:0] } )	// line#=../rle.cpp:111,140,141,142
		| ( { 8{ incr8u3i1_c2 } } & RG_len )				// line#=../rle.cpp:74
		) ;
	end
assign	incr32s1i1 = RG_i_k_01 ;	// line#=../rle.cpp:64,119,129,140,141
					// ,150,160
assign	incr32s2i1 = RG_i_j_01 ;	// line#=../rle.cpp:63,114,125,140,141
					// ,145,156
assign	decr32s1i1 = RG_i_k_01 ;	// line#=../rle.cpp:124,140,141,155
assign	decr32s2i1 = RG_i_j_01 ;	// line#=../rle.cpp:130,140,141,161
always @ ( RG_i_j_01 or U_174 or CT_28 or ST1_07d )	// line#=../rle.cpp:61,62
	begin
	zz_RA1_c1 = ( ( ST1_07d & CT_28 ) | U_174 ) ;	// line#=../rle.cpp:61,62,74
	zz_RA1 = ( { 6{ zz_RA1_c1 } } & RG_i_j_01 [5:0] )	// line#=../rle.cpp:61,62,74
		 ;	// line#=../rle.cpp:52,53
	end
always @ ( RG_quantized_block_rl_7 or RG_quantized_block_rl_6 or RG_quantized_block_rl_5 or 
	RG_quantized_block_rl_4 or RG_quantized_block_rl_3 or RG_quantized_block_rl_2 or 
	RG_quantized_block_rl_1 or RG_quantized_block_rl or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_03 = RG_quantized_block_rl ;	// line#=../rle.cpp:111
	3'h1 :
		TR_03 = RG_quantized_block_rl_1 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_03 = RG_quantized_block_rl_2 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_03 = RG_quantized_block_rl_3 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_03 = RG_quantized_block_rl_4 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_03 = RG_quantized_block_rl_5 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_03 = RG_quantized_block_rl_6 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_03 = RG_quantized_block_rl_7 ;	// line#=../rle.cpp:111
	default :
		TR_03 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_15 or RG_quantized_block_rl_14 or RG_quantized_block_rl_13 or 
	RG_quantized_block_rl_12 or RG_quantized_block_rl_11 or RG_quantized_block_rl_10 or 
	RG_quantized_block_rl_9 or RG_quantized_block_rl_8 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_04 = RG_quantized_block_rl_8 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_04 = RG_quantized_block_rl_9 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_04 = RG_quantized_block_rl_10 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_04 = RG_quantized_block_rl_11 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_04 = RG_quantized_block_rl_12 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_04 = RG_quantized_block_rl_13 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_04 = RG_quantized_block_rl_14 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_04 = RG_quantized_block_rl_15 ;	// line#=../rle.cpp:111
	default :
		TR_04 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_23 or RG_quantized_block_rl_22 or RG_quantized_block_rl_21 or 
	RG_quantized_block_rl_20 or RG_quantized_block_rl_19 or RG_quantized_block_rl_18 or 
	RG_quantized_block_rl_17 or RG_quantized_block_rl_16 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_05 = RG_quantized_block_rl_16 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_05 = RG_quantized_block_rl_17 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_05 = RG_quantized_block_rl_18 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_05 = RG_quantized_block_rl_19 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_05 = RG_quantized_block_rl_20 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_05 = RG_quantized_block_rl_21 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_05 = RG_quantized_block_rl_22 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_05 = RG_quantized_block_rl_23 ;	// line#=../rle.cpp:111
	default :
		TR_05 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_31 or RG_quantized_block_rl_30 or RG_quantized_block_rl_29 or 
	RG_quantized_block_rl_28 or RG_quantized_block_rl_27 or RG_quantized_block_rl_26 or 
	RG_quantized_block_rl_25 or RG_quantized_block_rl_24 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_06 = RG_quantized_block_rl_24 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_06 = RG_quantized_block_rl_25 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_06 = RG_quantized_block_rl_26 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_06 = RG_quantized_block_rl_27 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_06 = RG_quantized_block_rl_28 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_06 = RG_quantized_block_rl_29 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_06 = RG_quantized_block_rl_30 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_06 = RG_quantized_block_rl_31 ;	// line#=../rle.cpp:111
	default :
		TR_06 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_39 or RG_quantized_block_rl_38 or RG_quantized_block_rl_37 or 
	RG_quantized_block_rl_36 or RG_quantized_block_rl_35 or RG_quantized_block_rl_34 or 
	RG_quantized_block_rl_33 or RG_quantized_block_rl_32 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_07 = RG_quantized_block_rl_32 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_07 = RG_quantized_block_rl_33 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_07 = RG_quantized_block_rl_34 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_07 = RG_quantized_block_rl_35 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_07 = RG_quantized_block_rl_36 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_07 = RG_quantized_block_rl_37 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_07 = RG_quantized_block_rl_38 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_07 = RG_quantized_block_rl_39 ;	// line#=../rle.cpp:111
	default :
		TR_07 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_47 or RG_quantized_block_rl_46 or RG_quantized_block_rl_45 or 
	RG_quantized_block_rl_44 or RG_quantized_block_rl_43 or RG_quantized_block_rl_42 or 
	RG_quantized_block_rl_41 or RG_quantized_block_rl_40 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_08 = RG_quantized_block_rl_40 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_08 = RG_quantized_block_rl_41 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_08 = RG_quantized_block_rl_42 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_08 = RG_quantized_block_rl_43 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_08 = RG_quantized_block_rl_44 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_08 = RG_quantized_block_rl_45 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_08 = RG_quantized_block_rl_46 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_08 = RG_quantized_block_rl_47 ;	// line#=../rle.cpp:111
	default :
		TR_08 = 9'hx ;
	endcase
always @ ( RG_quantized_block_rl_55 or RG_quantized_block_rl_54 or RG_quantized_block_rl_53 or 
	RG_quantized_block_rl_52 or RG_quantized_block_rl_51 or RG_quantized_block_rl_50 or 
	RG_quantized_block_rl_49 or RG_quantized_block_rl_48 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_09 = RG_quantized_block_rl_48 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_09 = RG_quantized_block_rl_49 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_09 = RG_quantized_block_rl_50 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_09 = RG_quantized_block_rl_51 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_09 = RG_quantized_block_rl_52 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_09 = RG_quantized_block_rl_53 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_09 = RG_quantized_block_rl_54 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_09 = RG_quantized_block_rl_55 ;	// line#=../rle.cpp:111
	default :
		TR_09 = 9'hx ;
	endcase
always @ ( RL_previous_dc_quantized_block or RG_quantized_block_rl_62 or RG_quantized_block_rl_61 or 
	RG_quantized_block_rl_60 or RG_quantized_block_rl_59 or RG_quantized_block_rl_58 or 
	RG_quantized_block_rl_57 or RG_quantized_block_rl_56 or RG_i_j_01 )	// line#=../rle.cpp:111
	case ( RG_i_j_01 [2:0] )
	3'h0 :
		TR_10 = RG_quantized_block_rl_56 ;	// line#=../rle.cpp:111
	3'h1 :
		TR_10 = RG_quantized_block_rl_57 ;	// line#=../rle.cpp:111
	3'h2 :
		TR_10 = RG_quantized_block_rl_58 ;	// line#=../rle.cpp:111
	3'h3 :
		TR_10 = RG_quantized_block_rl_59 ;	// line#=../rle.cpp:111
	3'h4 :
		TR_10 = RG_quantized_block_rl_60 ;	// line#=../rle.cpp:111
	3'h5 :
		TR_10 = RG_quantized_block_rl_61 ;	// line#=../rle.cpp:111
	3'h6 :
		TR_10 = RG_quantized_block_rl_62 ;	// line#=../rle.cpp:111
	3'h7 :
		TR_10 = RL_previous_dc_quantized_block ;	// line#=../rle.cpp:111
	default :
		TR_10 = 9'hx ;
	endcase
always @ ( U_96 or U_95 or U_94 or U_93 or U_92 or U_91 or U_90 or U_89 or TR_10 or 
	U_14 or TR_09 or U_13 or TR_08 or U_12 or TR_07 or U_11 or TR_06 or U_10 or 
	TR_05 or U_09 or TR_04 or U_08 or TR_03 or U_07 )
	zz_WD2 = ( ( { 9{ U_07 } } & TR_03 )	// line#=../rle.cpp:111
		| ( { 9{ U_08 } } & TR_04 )	// line#=../rle.cpp:111
		| ( { 9{ U_09 } } & TR_05 )	// line#=../rle.cpp:111
		| ( { 9{ U_10 } } & TR_06 )	// line#=../rle.cpp:111
		| ( { 9{ U_11 } } & TR_07 )	// line#=../rle.cpp:111
		| ( { 9{ U_12 } } & TR_08 )	// line#=../rle.cpp:111
		| ( { 9{ U_13 } } & TR_09 )	// line#=../rle.cpp:111
		| ( { 9{ U_14 } } & TR_10 )	// line#=../rle.cpp:111
		| ( { 9{ U_89 } } & TR_03 )	// line#=../rle.cpp:140,141,142
		| ( { 9{ U_90 } } & TR_04 )	// line#=../rle.cpp:140,141,142
		| ( { 9{ U_91 } } & TR_05 )	// line#=../rle.cpp:140,141,142
		| ( { 9{ U_92 } } & TR_06 )	// line#=../rle.cpp:140,141,142
		| ( { 9{ U_93 } } & TR_07 )	// line#=../rle.cpp:140,141,142
		| ( { 9{ U_94 } } & TR_08 )	// line#=../rle.cpp:140,141,142
		| ( { 9{ U_95 } } & TR_09 )	// line#=../rle.cpp:140,141,142
		| ( { 9{ U_96 } } & TR_10 )	// line#=../rle.cpp:140,141,142
		) ;
assign	M_174 = ~|( RG_i_j_01 [2:0] ^ 3'h1 ) ;	// line#=../rle.cpp:111,140,141,142
assign	M_176 = ~|RG_i_j_01 [2:0] ;	// line#=../rle.cpp:111,140,141,142
assign	M_178 = ~|( RG_i_j_01 [2:0] ^ 3'h2 ) ;	// line#=../rle.cpp:111,140,141,142
assign	M_180 = ~|( RG_i_j_01 [2:0] ^ 3'h7 ) ;	// line#=../rle.cpp:111,140,141,142
assign	M_182 = ~|( RG_i_j_01 [2:0] ^ 3'h4 ) ;	// line#=../rle.cpp:111,140,141,142
assign	M_184 = ~|( RG_i_j_01 [2:0] ^ 3'h3 ) ;	// line#=../rle.cpp:111,140,141,142
assign	M_186 = ~|( RG_i_j_01 [2:0] ^ 3'h5 ) ;	// line#=../rle.cpp:111,140,141,142
assign	M_188 = ~|( RG_i_j_01 [2:0] ^ 3'h6 ) ;	// line#=../rle.cpp:111,140,141,142
assign	zz_WE2 = ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( 
	( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( ( U_14 & M_180 ) | ( U_14 & M_188 ) ) | 
	( U_14 & M_186 ) ) | ( U_14 & M_182 ) ) | ( U_14 & M_184 ) ) | ( U_14 & M_178 ) ) | 
	( U_14 & M_174 ) ) | ( U_14 & M_176 ) ) | ( U_13 & M_180 ) ) | ( U_13 & M_188 ) ) | 
	( U_13 & M_186 ) ) | ( U_13 & M_182 ) ) | ( U_13 & M_184 ) ) | ( U_13 & M_178 ) ) | 
	( U_13 & M_174 ) ) | ( U_13 & M_176 ) ) | ( U_12 & M_180 ) ) | ( U_12 & M_188 ) ) | 
	( U_12 & M_186 ) ) | ( U_12 & M_182 ) ) | ( U_12 & M_184 ) ) | ( U_12 & M_178 ) ) | 
	( U_12 & M_174 ) ) | ( U_12 & M_176 ) ) | ( U_11 & M_180 ) ) | ( U_11 & M_188 ) ) | 
	( U_11 & M_186 ) ) | ( U_11 & M_182 ) ) | ( U_11 & M_184 ) ) | ( U_11 & M_178 ) ) | 
	( U_11 & M_174 ) ) | ( U_11 & M_176 ) ) | ( U_10 & M_180 ) ) | ( U_10 & M_188 ) ) | 
	( U_10 & M_186 ) ) | ( U_10 & M_182 ) ) | ( U_10 & M_184 ) ) | ( U_10 & M_178 ) ) | 
	( U_10 & M_174 ) ) | ( U_10 & M_176 ) ) | ( U_09 & M_180 ) ) | ( U_09 & M_188 ) ) | 
	( U_09 & M_186 ) ) | ( U_09 & M_182 ) ) | ( U_09 & M_184 ) ) | ( U_09 & M_178 ) ) | 
	( U_09 & M_174 ) ) | ( U_09 & M_176 ) ) | ( U_08 & M_180 ) ) | ( U_08 & M_188 ) ) | 
	( U_08 & M_186 ) ) | ( U_08 & M_182 ) ) | ( U_08 & M_184 ) ) | ( U_08 & M_178 ) ) | 
	( U_08 & M_174 ) ) | ( U_08 & M_176 ) ) | ( U_07 & M_180 ) ) | ( U_07 & M_188 ) ) | 
	( U_07 & M_186 ) ) | ( U_07 & M_182 ) ) | ( U_07 & M_184 ) ) | ( U_07 & M_178 ) ) | 
	( U_07 & M_174 ) ) | ( U_07 & M_176 ) ) | ( U_89 & M_176 ) ) | ( U_89 & M_174 ) ) | 
	( U_89 & M_178 ) ) | ( U_89 & M_184 ) ) | ( U_89 & M_182 ) ) | ( U_89 & M_186 ) ) | 
	( U_89 & M_188 ) ) | ( U_89 & M_180 ) ) | ( U_90 & M_176 ) ) | ( U_90 & M_174 ) ) | 
	( U_90 & M_178 ) ) | ( U_90 & M_184 ) ) | ( U_90 & M_182 ) ) | ( U_90 & M_186 ) ) | 
	( U_90 & M_188 ) ) | ( U_90 & M_180 ) ) | ( U_91 & M_176 ) ) | ( U_91 & M_174 ) ) | 
	( U_91 & M_178 ) ) | ( U_91 & M_184 ) ) | ( U_91 & M_182 ) ) | ( U_91 & M_186 ) ) | 
	( U_91 & M_188 ) ) | ( U_91 & M_180 ) ) | ( U_92 & M_176 ) ) | ( U_92 & M_174 ) ) | 
	( U_92 & M_178 ) ) | ( U_92 & M_184 ) ) | ( U_92 & M_182 ) ) | ( U_92 & M_186 ) ) | 
	( U_92 & M_188 ) ) | ( U_92 & M_180 ) ) | ( U_93 & M_176 ) ) | ( U_93 & M_174 ) ) | 
	( U_93 & M_178 ) ) | ( U_93 & M_184 ) ) | ( U_93 & M_182 ) ) | ( U_93 & M_186 ) ) | 
	( U_93 & M_188 ) ) | ( U_93 & M_180 ) ) | ( U_94 & M_176 ) ) | ( U_94 & M_174 ) ) | 
	( U_94 & M_178 ) ) | ( U_94 & M_184 ) ) | ( U_94 & M_182 ) ) | ( U_94 & M_186 ) ) | 
	( U_94 & M_188 ) ) | ( U_94 & M_180 ) ) | ( U_95 & M_176 ) ) | ( U_95 & M_174 ) ) | 
	( U_95 & M_178 ) ) | ( U_95 & M_184 ) ) | ( U_95 & M_182 ) ) | ( U_95 & M_186 ) ) | 
	( U_95 & M_188 ) ) | ( U_95 & M_180 ) ) | ( U_96 & M_176 ) ) | ( U_96 & M_174 ) ) | 
	( U_96 & M_178 ) ) | ( U_96 & M_184 ) ) | ( U_96 & M_182 ) ) | ( U_96 & M_186 ) ) | 
	( U_96 & M_188 ) ) | ( U_96 & M_180 ) ) ;

endmodule

module jpeg_sub8u_7_1 ( i1 ,i2 ,o1 );
input	[6:0]	i1 ;
input	[1:0]	i2 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - { 5'h00 , i2 } ) ;

endmodule

module jpeg_sub8u_7 ( i1 ,i2 ,o1 );
input	[6:0]	i1 ;
input	[2:0]	i2 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - { 4'h0 , i2 } ) ;

endmodule

module jpeg_decr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_decr8u_7 ( i1 ,o1 );
input	[6:0]	i1 ;
output	[6:0]	o1 ;

assign	o1 = ( i1 - 1'h1 ) ;

endmodule

module jpeg_incr32s ( i1 ,o1 );
input	[31:0]	i1 ;
output	[31:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr8u ( i1 ,o1 );
input	[7:0]	i1 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_incr4s ( i1 ,o1 );
input	[3:0]	i1 ;
output	[3:0]	o1 ;

assign	o1 = ( i1 + 1'h1 ) ;

endmodule

module jpeg_lop8u_1 ( i1 ,i2 ,o1 );
input	[5:0]	i1 ;
input	[5:0]	i2 ;
output		o1 ;
wire		M_01 ;

assign	M_01 = ( i1 < i2 ) ;
assign	o1 = M_01 ;

endmodule

module jpeg_sub12s_9 ( i1 ,i2 ,o1 );
input	[8:0]	i1 ;
input	[8:0]	i2 ;
output	[8:0]	o1 ;

assign	o1 = ( i1 - i2 ) ;

endmodule

module jpeg_sub8u ( i1 ,i2 ,o1 );
input	[7:0]	i1 ;
input	[1:0]	i2 ;
output	[7:0]	o1 ;

assign	o1 = ( i1 - { 6'h00 , i2 } ) ;

endmodule

module jpeg_MEMB9W64 ( RA1 ,RD1 ,RCLK1 ,WA2 ,WD2 ,WE2 ,WCLK2 );
input	[5:0]	RA1 ;
output	[8:0]	RD1 ;
input		RCLK1 ;
input	[5:0]	WA2 ;
input	[8:0]	WD2 ;
input		WE2 ;
input		WCLK2 ;

jpeg_MEMB9W64_sub INST_MEMB9W64_sub_1 ( .RD1(RD1) ,.WE2(WE2) ,.WD2(WD2) ,.RA1(RA1) ,
	.WA2(WA2) ,.RCLK1(RCLK1) ,.WCLK2(WCLK2) );

endmodule

(* ram_extract = "yes" *)
module jpeg_MEMB9W64_sub ( RD1 ,WE2 ,WD2 ,RA1 ,WA2 ,RCLK1 ,WCLK2 );
output	[8:0]	RD1 ;
input		WE2 ;
input	[8:0]	WD2 ;
input	[5:0]	RA1 ;
input	[5:0]	WA2 ;
input		RCLK1 ;
input		WCLK2 ;
wire		Wen1_wire ;
reg	[8:0]	Rd1_sr	[0:0] ;
(* ram_style = "block" *)reg	[8:0]	MEMB9W64_r	[0:63] ;

assign	RD1 = Rd1_sr[0] ;
assign	Wen1_wire = WE2 ;

always @ ( posedge RCLK1 )
	begin
	Rd1_sr [0] <= MEMB9W64_r[RA1] ;
	end

always @ ( posedge WCLK2 )
	begin
	if ( Wen1_wire )
		begin
		MEMB9W64_r [WA2] <= WD2 ;
		end
	end

endmodule
